-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jan 27 2023 14:59:52

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "zim" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of zim
entity zim is
port (
    VAC_DRDY : in std_logic;
    IAC_FLT1 : out std_logic;
    DDS_SCK : out std_logic;
    ICE_IOR_166 : in std_logic;
    ICE_IOR_119 : in std_logic;
    DDS_MOSI : out std_logic;
    VAC_MISO : in std_logic;
    DDS_MOSI1 : out std_logic;
    ICE_IOR_146 : in std_logic;
    VDC_CLK : out std_logic;
    ICE_IOT_222 : in std_logic;
    IAC_CS : out std_logic;
    ICE_IOL_18B : in std_logic;
    ICE_IOL_13A : in std_logic;
    ICE_IOB_81 : in std_logic;
    VAC_OSR1 : out std_logic;
    IAC_MOSI : out std_logic;
    DDS_CS1 : out std_logic;
    ICE_IOL_4B : in std_logic;
    ICE_IOB_94 : in std_logic;
    VAC_CS : out std_logic;
    VAC_CLK : out std_logic;
    ICE_SPI_CE0 : in std_logic;
    ICE_IOR_167 : in std_logic;
    ICE_IOR_118 : in std_logic;
    RTD_SDO : in std_logic;
    IAC_OSR0 : out std_logic;
    VDC_SCLK : out std_logic;
    VAC_FLT1 : out std_logic;
    ICE_SPI_MOSI : in std_logic;
    ICE_IOR_165 : in std_logic;
    ICE_IOR_147 : in std_logic;
    ICE_IOL_14A : in std_logic;
    ICE_IOL_13B : in std_logic;
    ICE_IOB_91 : in std_logic;
    ICE_GPMO_0 : in std_logic;
    DDS_RNG_0 : out std_logic;
    VDC_RNG0 : out std_logic;
    ICE_SPI_SCLK : in std_logic;
    ICE_IOR_152 : in std_logic;
    ICE_IOL_12A : in std_logic;
    RTD_DRDY : in std_logic;
    ICE_SPI_MISO : out std_logic;
    ICE_IOT_177 : in std_logic;
    ICE_IOR_141 : in std_logic;
    ICE_IOB_80 : in std_logic;
    ICE_IOB_102 : in std_logic;
    ICE_GPMO_2 : in std_logic;
    ICE_GPMI_0 : out std_logic;
    IAC_MISO : in std_logic;
    VAC_OSR0 : out std_logic;
    VAC_MOSI : out std_logic;
    TEST_LED : out std_logic;
    ICE_IOR_148 : in std_logic;
    STAT_COMM : out std_logic;
    ICE_SYSCLK : in std_logic;
    ICE_IOR_161 : in std_logic;
    ICE_IOB_95 : in std_logic;
    ICE_IOB_82 : in std_logic;
    ICE_IOB_104 : in std_logic;
    IAC_CLK : out std_logic;
    DDS_CS : out std_logic;
    SELIRNG0 : out std_logic;
    RTD_SDI : out std_logic;
    ICE_IOT_221 : in std_logic;
    ICE_IOT_197 : in std_logic;
    DDS_MCLK : out std_logic;
    RTD_SCLK : out std_logic;
    RTD_CS : out std_logic;
    ICE_IOR_137 : in std_logic;
    IAC_OSR1 : out std_logic;
    VAC_FLT0 : out std_logic;
    ICE_IOR_144 : in std_logic;
    ICE_IOR_128 : in std_logic;
    ICE_GPMO_1 : in std_logic;
    IAC_SCLK : out std_logic;
    EIS_SYNCCLK : in std_logic;
    ICE_IOR_139 : in std_logic;
    ICE_IOL_4A : in std_logic;
    VAC_SCLK : out std_logic;
    THERMOSTAT : in std_logic;
    ICE_IOR_164 : in std_logic;
    ICE_IOB_103 : in std_logic;
    AMPV_POW : out std_logic;
    VDC_SDO : in std_logic;
    ICE_IOT_174 : in std_logic;
    ICE_IOR_140 : in std_logic;
    ICE_IOB_96 : in std_logic;
    CONT_SD : out std_logic;
    AC_ADC_SYNC : out std_logic;
    SELIRNG1 : out std_logic;
    ICE_IOL_12B : in std_logic;
    ICE_IOR_160 : in std_logic;
    ICE_IOR_136 : in std_logic;
    DDS_MCLK1 : out std_logic;
    ICE_IOT_198 : in std_logic;
    ICE_IOT_173 : in std_logic;
    IAC_DRDY : in std_logic;
    ICE_IOT_178 : in std_logic;
    ICE_IOR_138 : in std_logic;
    ICE_IOR_120 : in std_logic;
    IAC_FLT0 : out std_logic;
    DDS_SCK1 : out std_logic);
end zim;

-- Architecture of zim
-- View name is \INTERFACE\
architecture \INTERFACE\ of zim is

signal \N__58652\ : std_logic;
signal \N__58651\ : std_logic;
signal \N__58650\ : std_logic;
signal \N__58643\ : std_logic;
signal \N__58642\ : std_logic;
signal \N__58641\ : std_logic;
signal \N__58634\ : std_logic;
signal \N__58633\ : std_logic;
signal \N__58632\ : std_logic;
signal \N__58625\ : std_logic;
signal \N__58624\ : std_logic;
signal \N__58623\ : std_logic;
signal \N__58616\ : std_logic;
signal \N__58615\ : std_logic;
signal \N__58614\ : std_logic;
signal \N__58607\ : std_logic;
signal \N__58606\ : std_logic;
signal \N__58605\ : std_logic;
signal \N__58598\ : std_logic;
signal \N__58597\ : std_logic;
signal \N__58596\ : std_logic;
signal \N__58589\ : std_logic;
signal \N__58588\ : std_logic;
signal \N__58587\ : std_logic;
signal \N__58580\ : std_logic;
signal \N__58579\ : std_logic;
signal \N__58578\ : std_logic;
signal \N__58571\ : std_logic;
signal \N__58570\ : std_logic;
signal \N__58569\ : std_logic;
signal \N__58562\ : std_logic;
signal \N__58561\ : std_logic;
signal \N__58560\ : std_logic;
signal \N__58553\ : std_logic;
signal \N__58552\ : std_logic;
signal \N__58551\ : std_logic;
signal \N__58544\ : std_logic;
signal \N__58543\ : std_logic;
signal \N__58542\ : std_logic;
signal \N__58535\ : std_logic;
signal \N__58534\ : std_logic;
signal \N__58533\ : std_logic;
signal \N__58526\ : std_logic;
signal \N__58525\ : std_logic;
signal \N__58524\ : std_logic;
signal \N__58517\ : std_logic;
signal \N__58516\ : std_logic;
signal \N__58515\ : std_logic;
signal \N__58508\ : std_logic;
signal \N__58507\ : std_logic;
signal \N__58506\ : std_logic;
signal \N__58499\ : std_logic;
signal \N__58498\ : std_logic;
signal \N__58497\ : std_logic;
signal \N__58490\ : std_logic;
signal \N__58489\ : std_logic;
signal \N__58488\ : std_logic;
signal \N__58481\ : std_logic;
signal \N__58480\ : std_logic;
signal \N__58479\ : std_logic;
signal \N__58472\ : std_logic;
signal \N__58471\ : std_logic;
signal \N__58470\ : std_logic;
signal \N__58463\ : std_logic;
signal \N__58462\ : std_logic;
signal \N__58461\ : std_logic;
signal \N__58454\ : std_logic;
signal \N__58453\ : std_logic;
signal \N__58452\ : std_logic;
signal \N__58445\ : std_logic;
signal \N__58444\ : std_logic;
signal \N__58443\ : std_logic;
signal \N__58436\ : std_logic;
signal \N__58435\ : std_logic;
signal \N__58434\ : std_logic;
signal \N__58427\ : std_logic;
signal \N__58426\ : std_logic;
signal \N__58425\ : std_logic;
signal \N__58418\ : std_logic;
signal \N__58417\ : std_logic;
signal \N__58416\ : std_logic;
signal \N__58409\ : std_logic;
signal \N__58408\ : std_logic;
signal \N__58407\ : std_logic;
signal \N__58400\ : std_logic;
signal \N__58399\ : std_logic;
signal \N__58398\ : std_logic;
signal \N__58391\ : std_logic;
signal \N__58390\ : std_logic;
signal \N__58389\ : std_logic;
signal \N__58382\ : std_logic;
signal \N__58381\ : std_logic;
signal \N__58380\ : std_logic;
signal \N__58373\ : std_logic;
signal \N__58372\ : std_logic;
signal \N__58371\ : std_logic;
signal \N__58364\ : std_logic;
signal \N__58363\ : std_logic;
signal \N__58362\ : std_logic;
signal \N__58355\ : std_logic;
signal \N__58354\ : std_logic;
signal \N__58353\ : std_logic;
signal \N__58346\ : std_logic;
signal \N__58345\ : std_logic;
signal \N__58344\ : std_logic;
signal \N__58337\ : std_logic;
signal \N__58336\ : std_logic;
signal \N__58335\ : std_logic;
signal \N__58328\ : std_logic;
signal \N__58327\ : std_logic;
signal \N__58326\ : std_logic;
signal \N__58319\ : std_logic;
signal \N__58318\ : std_logic;
signal \N__58317\ : std_logic;
signal \N__58310\ : std_logic;
signal \N__58309\ : std_logic;
signal \N__58308\ : std_logic;
signal \N__58301\ : std_logic;
signal \N__58300\ : std_logic;
signal \N__58299\ : std_logic;
signal \N__58292\ : std_logic;
signal \N__58291\ : std_logic;
signal \N__58290\ : std_logic;
signal \N__58283\ : std_logic;
signal \N__58282\ : std_logic;
signal \N__58281\ : std_logic;
signal \N__58274\ : std_logic;
signal \N__58273\ : std_logic;
signal \N__58272\ : std_logic;
signal \N__58265\ : std_logic;
signal \N__58264\ : std_logic;
signal \N__58263\ : std_logic;
signal \N__58256\ : std_logic;
signal \N__58255\ : std_logic;
signal \N__58254\ : std_logic;
signal \N__58247\ : std_logic;
signal \N__58246\ : std_logic;
signal \N__58245\ : std_logic;
signal \N__58238\ : std_logic;
signal \N__58237\ : std_logic;
signal \N__58236\ : std_logic;
signal \N__58229\ : std_logic;
signal \N__58228\ : std_logic;
signal \N__58227\ : std_logic;
signal \N__58220\ : std_logic;
signal \N__58219\ : std_logic;
signal \N__58218\ : std_logic;
signal \N__58211\ : std_logic;
signal \N__58210\ : std_logic;
signal \N__58209\ : std_logic;
signal \N__58202\ : std_logic;
signal \N__58201\ : std_logic;
signal \N__58200\ : std_logic;
signal \N__58193\ : std_logic;
signal \N__58192\ : std_logic;
signal \N__58191\ : std_logic;
signal \N__58184\ : std_logic;
signal \N__58183\ : std_logic;
signal \N__58182\ : std_logic;
signal \N__58175\ : std_logic;
signal \N__58174\ : std_logic;
signal \N__58173\ : std_logic;
signal \N__58166\ : std_logic;
signal \N__58165\ : std_logic;
signal \N__58164\ : std_logic;
signal \N__58157\ : std_logic;
signal \N__58156\ : std_logic;
signal \N__58155\ : std_logic;
signal \N__58148\ : std_logic;
signal \N__58147\ : std_logic;
signal \N__58146\ : std_logic;
signal \N__58139\ : std_logic;
signal \N__58138\ : std_logic;
signal \N__58137\ : std_logic;
signal \N__58130\ : std_logic;
signal \N__58129\ : std_logic;
signal \N__58128\ : std_logic;
signal \N__58121\ : std_logic;
signal \N__58120\ : std_logic;
signal \N__58119\ : std_logic;
signal \N__58112\ : std_logic;
signal \N__58111\ : std_logic;
signal \N__58110\ : std_logic;
signal \N__58103\ : std_logic;
signal \N__58102\ : std_logic;
signal \N__58101\ : std_logic;
signal \N__58094\ : std_logic;
signal \N__58093\ : std_logic;
signal \N__58092\ : std_logic;
signal \N__58085\ : std_logic;
signal \N__58084\ : std_logic;
signal \N__58083\ : std_logic;
signal \N__58076\ : std_logic;
signal \N__58075\ : std_logic;
signal \N__58074\ : std_logic;
signal \N__58067\ : std_logic;
signal \N__58066\ : std_logic;
signal \N__58065\ : std_logic;
signal \N__58058\ : std_logic;
signal \N__58057\ : std_logic;
signal \N__58056\ : std_logic;
signal \N__58049\ : std_logic;
signal \N__58048\ : std_logic;
signal \N__58047\ : std_logic;
signal \N__58040\ : std_logic;
signal \N__58039\ : std_logic;
signal \N__58038\ : std_logic;
signal \N__58031\ : std_logic;
signal \N__58030\ : std_logic;
signal \N__58029\ : std_logic;
signal \N__58022\ : std_logic;
signal \N__58021\ : std_logic;
signal \N__58020\ : std_logic;
signal \N__58013\ : std_logic;
signal \N__58012\ : std_logic;
signal \N__58011\ : std_logic;
signal \N__58004\ : std_logic;
signal \N__58003\ : std_logic;
signal \N__58002\ : std_logic;
signal \N__57995\ : std_logic;
signal \N__57994\ : std_logic;
signal \N__57993\ : std_logic;
signal \N__57986\ : std_logic;
signal \N__57985\ : std_logic;
signal \N__57984\ : std_logic;
signal \N__57977\ : std_logic;
signal \N__57976\ : std_logic;
signal \N__57975\ : std_logic;
signal \N__57968\ : std_logic;
signal \N__57967\ : std_logic;
signal \N__57966\ : std_logic;
signal \N__57959\ : std_logic;
signal \N__57958\ : std_logic;
signal \N__57957\ : std_logic;
signal \N__57950\ : std_logic;
signal \N__57949\ : std_logic;
signal \N__57948\ : std_logic;
signal \N__57941\ : std_logic;
signal \N__57940\ : std_logic;
signal \N__57939\ : std_logic;
signal \N__57932\ : std_logic;
signal \N__57931\ : std_logic;
signal \N__57930\ : std_logic;
signal \N__57923\ : std_logic;
signal \N__57922\ : std_logic;
signal \N__57921\ : std_logic;
signal \N__57914\ : std_logic;
signal \N__57913\ : std_logic;
signal \N__57912\ : std_logic;
signal \N__57905\ : std_logic;
signal \N__57904\ : std_logic;
signal \N__57903\ : std_logic;
signal \N__57896\ : std_logic;
signal \N__57895\ : std_logic;
signal \N__57894\ : std_logic;
signal \N__57887\ : std_logic;
signal \N__57886\ : std_logic;
signal \N__57885\ : std_logic;
signal \N__57878\ : std_logic;
signal \N__57877\ : std_logic;
signal \N__57876\ : std_logic;
signal \N__57869\ : std_logic;
signal \N__57868\ : std_logic;
signal \N__57867\ : std_logic;
signal \N__57860\ : std_logic;
signal \N__57859\ : std_logic;
signal \N__57858\ : std_logic;
signal \N__57851\ : std_logic;
signal \N__57850\ : std_logic;
signal \N__57849\ : std_logic;
signal \N__57842\ : std_logic;
signal \N__57841\ : std_logic;
signal \N__57840\ : std_logic;
signal \N__57833\ : std_logic;
signal \N__57832\ : std_logic;
signal \N__57831\ : std_logic;
signal \N__57824\ : std_logic;
signal \N__57823\ : std_logic;
signal \N__57822\ : std_logic;
signal \N__57815\ : std_logic;
signal \N__57814\ : std_logic;
signal \N__57813\ : std_logic;
signal \N__57806\ : std_logic;
signal \N__57805\ : std_logic;
signal \N__57804\ : std_logic;
signal \N__57797\ : std_logic;
signal \N__57796\ : std_logic;
signal \N__57795\ : std_logic;
signal \N__57788\ : std_logic;
signal \N__57787\ : std_logic;
signal \N__57786\ : std_logic;
signal \N__57779\ : std_logic;
signal \N__57778\ : std_logic;
signal \N__57777\ : std_logic;
signal \N__57770\ : std_logic;
signal \N__57769\ : std_logic;
signal \N__57768\ : std_logic;
signal \N__57761\ : std_logic;
signal \N__57760\ : std_logic;
signal \N__57759\ : std_logic;
signal \N__57752\ : std_logic;
signal \N__57751\ : std_logic;
signal \N__57750\ : std_logic;
signal \N__57743\ : std_logic;
signal \N__57742\ : std_logic;
signal \N__57741\ : std_logic;
signal \N__57734\ : std_logic;
signal \N__57733\ : std_logic;
signal \N__57732\ : std_logic;
signal \N__57715\ : std_logic;
signal \N__57714\ : std_logic;
signal \N__57711\ : std_logic;
signal \N__57708\ : std_logic;
signal \N__57705\ : std_logic;
signal \N__57700\ : std_logic;
signal \N__57697\ : std_logic;
signal \N__57694\ : std_logic;
signal \N__57693\ : std_logic;
signal \N__57690\ : std_logic;
signal \N__57687\ : std_logic;
signal \N__57684\ : std_logic;
signal \N__57679\ : std_logic;
signal \N__57676\ : std_logic;
signal \N__57673\ : std_logic;
signal \N__57670\ : std_logic;
signal \N__57669\ : std_logic;
signal \N__57666\ : std_logic;
signal \N__57663\ : std_logic;
signal \N__57660\ : std_logic;
signal \N__57655\ : std_logic;
signal \N__57652\ : std_logic;
signal \N__57651\ : std_logic;
signal \N__57648\ : std_logic;
signal \N__57645\ : std_logic;
signal \N__57642\ : std_logic;
signal \N__57637\ : std_logic;
signal \N__57634\ : std_logic;
signal \N__57633\ : std_logic;
signal \N__57630\ : std_logic;
signal \N__57627\ : std_logic;
signal \N__57624\ : std_logic;
signal \N__57619\ : std_logic;
signal \N__57616\ : std_logic;
signal \N__57615\ : std_logic;
signal \N__57612\ : std_logic;
signal \N__57609\ : std_logic;
signal \N__57606\ : std_logic;
signal \N__57601\ : std_logic;
signal \N__57598\ : std_logic;
signal \N__57595\ : std_logic;
signal \N__57592\ : std_logic;
signal \N__57589\ : std_logic;
signal \N__57588\ : std_logic;
signal \N__57583\ : std_logic;
signal \N__57580\ : std_logic;
signal \N__57577\ : std_logic;
signal \N__57574\ : std_logic;
signal \N__57571\ : std_logic;
signal \N__57568\ : std_logic;
signal \N__57567\ : std_logic;
signal \N__57564\ : std_logic;
signal \N__57561\ : std_logic;
signal \N__57558\ : std_logic;
signal \N__57553\ : std_logic;
signal \N__57552\ : std_logic;
signal \N__57551\ : std_logic;
signal \N__57550\ : std_logic;
signal \N__57549\ : std_logic;
signal \N__57548\ : std_logic;
signal \N__57547\ : std_logic;
signal \N__57544\ : std_logic;
signal \N__57543\ : std_logic;
signal \N__57542\ : std_logic;
signal \N__57541\ : std_logic;
signal \N__57540\ : std_logic;
signal \N__57539\ : std_logic;
signal \N__57538\ : std_logic;
signal \N__57537\ : std_logic;
signal \N__57536\ : std_logic;
signal \N__57535\ : std_logic;
signal \N__57534\ : std_logic;
signal \N__57533\ : std_logic;
signal \N__57532\ : std_logic;
signal \N__57531\ : std_logic;
signal \N__57526\ : std_logic;
signal \N__57525\ : std_logic;
signal \N__57524\ : std_logic;
signal \N__57523\ : std_logic;
signal \N__57522\ : std_logic;
signal \N__57521\ : std_logic;
signal \N__57516\ : std_logic;
signal \N__57513\ : std_logic;
signal \N__57510\ : std_logic;
signal \N__57507\ : std_logic;
signal \N__57504\ : std_logic;
signal \N__57503\ : std_logic;
signal \N__57502\ : std_logic;
signal \N__57497\ : std_logic;
signal \N__57494\ : std_logic;
signal \N__57493\ : std_logic;
signal \N__57490\ : std_logic;
signal \N__57489\ : std_logic;
signal \N__57486\ : std_logic;
signal \N__57485\ : std_logic;
signal \N__57484\ : std_logic;
signal \N__57483\ : std_logic;
signal \N__57482\ : std_logic;
signal \N__57481\ : std_logic;
signal \N__57480\ : std_logic;
signal \N__57479\ : std_logic;
signal \N__57472\ : std_logic;
signal \N__57469\ : std_logic;
signal \N__57466\ : std_logic;
signal \N__57465\ : std_logic;
signal \N__57464\ : std_logic;
signal \N__57463\ : std_logic;
signal \N__57462\ : std_logic;
signal \N__57459\ : std_logic;
signal \N__57456\ : std_logic;
signal \N__57453\ : std_logic;
signal \N__57450\ : std_logic;
signal \N__57449\ : std_logic;
signal \N__57448\ : std_logic;
signal \N__57447\ : std_logic;
signal \N__57446\ : std_logic;
signal \N__57445\ : std_logic;
signal \N__57444\ : std_logic;
signal \N__57443\ : std_logic;
signal \N__57442\ : std_logic;
signal \N__57441\ : std_logic;
signal \N__57440\ : std_logic;
signal \N__57437\ : std_logic;
signal \N__57436\ : std_logic;
signal \N__57433\ : std_logic;
signal \N__57430\ : std_logic;
signal \N__57427\ : std_logic;
signal \N__57422\ : std_logic;
signal \N__57419\ : std_logic;
signal \N__57414\ : std_logic;
signal \N__57411\ : std_logic;
signal \N__57410\ : std_logic;
signal \N__57409\ : std_logic;
signal \N__57408\ : std_logic;
signal \N__57407\ : std_logic;
signal \N__57404\ : std_logic;
signal \N__57399\ : std_logic;
signal \N__57396\ : std_logic;
signal \N__57395\ : std_logic;
signal \N__57394\ : std_logic;
signal \N__57393\ : std_logic;
signal \N__57392\ : std_logic;
signal \N__57391\ : std_logic;
signal \N__57390\ : std_logic;
signal \N__57389\ : std_logic;
signal \N__57388\ : std_logic;
signal \N__57387\ : std_logic;
signal \N__57386\ : std_logic;
signal \N__57383\ : std_logic;
signal \N__57380\ : std_logic;
signal \N__57377\ : std_logic;
signal \N__57374\ : std_logic;
signal \N__57371\ : std_logic;
signal \N__57370\ : std_logic;
signal \N__57367\ : std_logic;
signal \N__57364\ : std_logic;
signal \N__57359\ : std_logic;
signal \N__57356\ : std_logic;
signal \N__57353\ : std_logic;
signal \N__57350\ : std_logic;
signal \N__57347\ : std_logic;
signal \N__57346\ : std_logic;
signal \N__57345\ : std_logic;
signal \N__57342\ : std_logic;
signal \N__57341\ : std_logic;
signal \N__57334\ : std_logic;
signal \N__57331\ : std_logic;
signal \N__57328\ : std_logic;
signal \N__57323\ : std_logic;
signal \N__57318\ : std_logic;
signal \N__57315\ : std_logic;
signal \N__57312\ : std_logic;
signal \N__57311\ : std_logic;
signal \N__57310\ : std_logic;
signal \N__57305\ : std_logic;
signal \N__57300\ : std_logic;
signal \N__57297\ : std_logic;
signal \N__57294\ : std_logic;
signal \N__57291\ : std_logic;
signal \N__57288\ : std_logic;
signal \N__57279\ : std_logic;
signal \N__57274\ : std_logic;
signal \N__57271\ : std_logic;
signal \N__57262\ : std_logic;
signal \N__57259\ : std_logic;
signal \N__57254\ : std_logic;
signal \N__57251\ : std_logic;
signal \N__57250\ : std_logic;
signal \N__57243\ : std_logic;
signal \N__57242\ : std_logic;
signal \N__57241\ : std_logic;
signal \N__57238\ : std_logic;
signal \N__57233\ : std_logic;
signal \N__57230\ : std_logic;
signal \N__57225\ : std_logic;
signal \N__57220\ : std_logic;
signal \N__57215\ : std_logic;
signal \N__57212\ : std_logic;
signal \N__57209\ : std_logic;
signal \N__57206\ : std_logic;
signal \N__57193\ : std_logic;
signal \N__57192\ : std_logic;
signal \N__57191\ : std_logic;
signal \N__57190\ : std_logic;
signal \N__57189\ : std_logic;
signal \N__57188\ : std_logic;
signal \N__57187\ : std_logic;
signal \N__57186\ : std_logic;
signal \N__57185\ : std_logic;
signal \N__57184\ : std_logic;
signal \N__57183\ : std_logic;
signal \N__57182\ : std_logic;
signal \N__57181\ : std_logic;
signal \N__57172\ : std_logic;
signal \N__57163\ : std_logic;
signal \N__57160\ : std_logic;
signal \N__57157\ : std_logic;
signal \N__57154\ : std_logic;
signal \N__57149\ : std_logic;
signal \N__57142\ : std_logic;
signal \N__57135\ : std_logic;
signal \N__57126\ : std_logic;
signal \N__57119\ : std_logic;
signal \N__57116\ : std_logic;
signal \N__57113\ : std_logic;
signal \N__57108\ : std_logic;
signal \N__57091\ : std_logic;
signal \N__57086\ : std_logic;
signal \N__57081\ : std_logic;
signal \N__57074\ : std_logic;
signal \N__57071\ : std_logic;
signal \N__57064\ : std_logic;
signal \N__57061\ : std_logic;
signal \N__57058\ : std_logic;
signal \N__57055\ : std_logic;
signal \N__57050\ : std_logic;
signal \N__57045\ : std_logic;
signal \N__57040\ : std_logic;
signal \N__57037\ : std_logic;
signal \N__57032\ : std_logic;
signal \N__57029\ : std_logic;
signal \N__57018\ : std_logic;
signal \N__56989\ : std_logic;
signal \N__56988\ : std_logic;
signal \N__56985\ : std_logic;
signal \N__56984\ : std_logic;
signal \N__56983\ : std_logic;
signal \N__56982\ : std_logic;
signal \N__56979\ : std_logic;
signal \N__56978\ : std_logic;
signal \N__56977\ : std_logic;
signal \N__56974\ : std_logic;
signal \N__56969\ : std_logic;
signal \N__56968\ : std_logic;
signal \N__56967\ : std_logic;
signal \N__56966\ : std_logic;
signal \N__56965\ : std_logic;
signal \N__56964\ : std_logic;
signal \N__56961\ : std_logic;
signal \N__56960\ : std_logic;
signal \N__56959\ : std_logic;
signal \N__56958\ : std_logic;
signal \N__56957\ : std_logic;
signal \N__56956\ : std_logic;
signal \N__56955\ : std_logic;
signal \N__56954\ : std_logic;
signal \N__56953\ : std_logic;
signal \N__56952\ : std_logic;
signal \N__56951\ : std_logic;
signal \N__56950\ : std_logic;
signal \N__56949\ : std_logic;
signal \N__56946\ : std_logic;
signal \N__56945\ : std_logic;
signal \N__56942\ : std_logic;
signal \N__56941\ : std_logic;
signal \N__56940\ : std_logic;
signal \N__56939\ : std_logic;
signal \N__56938\ : std_logic;
signal \N__56935\ : std_logic;
signal \N__56934\ : std_logic;
signal \N__56933\ : std_logic;
signal \N__56932\ : std_logic;
signal \N__56931\ : std_logic;
signal \N__56930\ : std_logic;
signal \N__56929\ : std_logic;
signal \N__56928\ : std_logic;
signal \N__56927\ : std_logic;
signal \N__56922\ : std_logic;
signal \N__56921\ : std_logic;
signal \N__56918\ : std_logic;
signal \N__56915\ : std_logic;
signal \N__56914\ : std_logic;
signal \N__56913\ : std_logic;
signal \N__56912\ : std_logic;
signal \N__56911\ : std_logic;
signal \N__56910\ : std_logic;
signal \N__56909\ : std_logic;
signal \N__56908\ : std_logic;
signal \N__56907\ : std_logic;
signal \N__56906\ : std_logic;
signal \N__56905\ : std_logic;
signal \N__56904\ : std_logic;
signal \N__56903\ : std_logic;
signal \N__56902\ : std_logic;
signal \N__56901\ : std_logic;
signal \N__56898\ : std_logic;
signal \N__56897\ : std_logic;
signal \N__56894\ : std_logic;
signal \N__56891\ : std_logic;
signal \N__56890\ : std_logic;
signal \N__56889\ : std_logic;
signal \N__56888\ : std_logic;
signal \N__56887\ : std_logic;
signal \N__56886\ : std_logic;
signal \N__56885\ : std_logic;
signal \N__56884\ : std_logic;
signal \N__56883\ : std_logic;
signal \N__56880\ : std_logic;
signal \N__56875\ : std_logic;
signal \N__56868\ : std_logic;
signal \N__56867\ : std_logic;
signal \N__56866\ : std_logic;
signal \N__56865\ : std_logic;
signal \N__56860\ : std_logic;
signal \N__56855\ : std_logic;
signal \N__56848\ : std_logic;
signal \N__56845\ : std_logic;
signal \N__56842\ : std_logic;
signal \N__56841\ : std_logic;
signal \N__56840\ : std_logic;
signal \N__56837\ : std_logic;
signal \N__56834\ : std_logic;
signal \N__56833\ : std_logic;
signal \N__56832\ : std_logic;
signal \N__56831\ : std_logic;
signal \N__56824\ : std_logic;
signal \N__56811\ : std_logic;
signal \N__56804\ : std_logic;
signal \N__56803\ : std_logic;
signal \N__56802\ : std_logic;
signal \N__56801\ : std_logic;
signal \N__56800\ : std_logic;
signal \N__56799\ : std_logic;
signal \N__56798\ : std_logic;
signal \N__56797\ : std_logic;
signal \N__56794\ : std_logic;
signal \N__56791\ : std_logic;
signal \N__56786\ : std_logic;
signal \N__56781\ : std_logic;
signal \N__56778\ : std_logic;
signal \N__56775\ : std_logic;
signal \N__56772\ : std_logic;
signal \N__56763\ : std_logic;
signal \N__56760\ : std_logic;
signal \N__56757\ : std_logic;
signal \N__56754\ : std_logic;
signal \N__56749\ : std_logic;
signal \N__56746\ : std_logic;
signal \N__56743\ : std_logic;
signal \N__56738\ : std_logic;
signal \N__56733\ : std_logic;
signal \N__56730\ : std_logic;
signal \N__56727\ : std_logic;
signal \N__56726\ : std_logic;
signal \N__56725\ : std_logic;
signal \N__56722\ : std_logic;
signal \N__56717\ : std_logic;
signal \N__56714\ : std_logic;
signal \N__56707\ : std_logic;
signal \N__56700\ : std_logic;
signal \N__56699\ : std_logic;
signal \N__56698\ : std_logic;
signal \N__56695\ : std_logic;
signal \N__56694\ : std_logic;
signal \N__56693\ : std_logic;
signal \N__56690\ : std_logic;
signal \N__56687\ : std_logic;
signal \N__56686\ : std_logic;
signal \N__56685\ : std_logic;
signal \N__56684\ : std_logic;
signal \N__56683\ : std_logic;
signal \N__56678\ : std_logic;
signal \N__56675\ : std_logic;
signal \N__56672\ : std_logic;
signal \N__56667\ : std_logic;
signal \N__56662\ : std_logic;
signal \N__56659\ : std_logic;
signal \N__56652\ : std_logic;
signal \N__56649\ : std_logic;
signal \N__56646\ : std_logic;
signal \N__56643\ : std_logic;
signal \N__56642\ : std_logic;
signal \N__56641\ : std_logic;
signal \N__56640\ : std_logic;
signal \N__56639\ : std_logic;
signal \N__56638\ : std_logic;
signal \N__56637\ : std_logic;
signal \N__56636\ : std_logic;
signal \N__56635\ : std_logic;
signal \N__56634\ : std_logic;
signal \N__56625\ : std_logic;
signal \N__56616\ : std_logic;
signal \N__56607\ : std_logic;
signal \N__56598\ : std_logic;
signal \N__56595\ : std_logic;
signal \N__56584\ : std_logic;
signal \N__56579\ : std_logic;
signal \N__56568\ : std_logic;
signal \N__56567\ : std_logic;
signal \N__56564\ : std_logic;
signal \N__56563\ : std_logic;
signal \N__56562\ : std_logic;
signal \N__56559\ : std_logic;
signal \N__56556\ : std_logic;
signal \N__56551\ : std_logic;
signal \N__56546\ : std_logic;
signal \N__56543\ : std_logic;
signal \N__56536\ : std_logic;
signal \N__56533\ : std_logic;
signal \N__56528\ : std_logic;
signal \N__56517\ : std_logic;
signal \N__56512\ : std_logic;
signal \N__56509\ : std_logic;
signal \N__56502\ : std_logic;
signal \N__56499\ : std_logic;
signal \N__56490\ : std_logic;
signal \N__56487\ : std_logic;
signal \N__56480\ : std_logic;
signal \N__56471\ : std_logic;
signal \N__56462\ : std_logic;
signal \N__56451\ : std_logic;
signal \N__56446\ : std_logic;
signal \N__56441\ : std_logic;
signal \N__56416\ : std_logic;
signal \N__56413\ : std_logic;
signal \N__56410\ : std_logic;
signal \N__56407\ : std_logic;
signal \N__56404\ : std_logic;
signal \N__56401\ : std_logic;
signal \N__56398\ : std_logic;
signal \N__56397\ : std_logic;
signal \N__56394\ : std_logic;
signal \N__56391\ : std_logic;
signal \N__56388\ : std_logic;
signal \N__56387\ : std_logic;
signal \N__56382\ : std_logic;
signal \N__56379\ : std_logic;
signal \N__56374\ : std_logic;
signal \N__56371\ : std_logic;
signal \N__56368\ : std_logic;
signal \N__56365\ : std_logic;
signal \N__56362\ : std_logic;
signal \N__56359\ : std_logic;
signal \N__56356\ : std_logic;
signal \N__56353\ : std_logic;
signal \N__56350\ : std_logic;
signal \N__56347\ : std_logic;
signal \N__56346\ : std_logic;
signal \N__56345\ : std_logic;
signal \N__56344\ : std_logic;
signal \N__56343\ : std_logic;
signal \N__56342\ : std_logic;
signal \N__56341\ : std_logic;
signal \N__56340\ : std_logic;
signal \N__56339\ : std_logic;
signal \N__56338\ : std_logic;
signal \N__56337\ : std_logic;
signal \N__56336\ : std_logic;
signal \N__56335\ : std_logic;
signal \N__56334\ : std_logic;
signal \N__56331\ : std_logic;
signal \N__56326\ : std_logic;
signal \N__56321\ : std_logic;
signal \N__56318\ : std_logic;
signal \N__56317\ : std_logic;
signal \N__56316\ : std_logic;
signal \N__56315\ : std_logic;
signal \N__56312\ : std_logic;
signal \N__56311\ : std_logic;
signal \N__56310\ : std_logic;
signal \N__56309\ : std_logic;
signal \N__56308\ : std_logic;
signal \N__56301\ : std_logic;
signal \N__56296\ : std_logic;
signal \N__56291\ : std_logic;
signal \N__56290\ : std_logic;
signal \N__56289\ : std_logic;
signal \N__56288\ : std_logic;
signal \N__56287\ : std_logic;
signal \N__56284\ : std_logic;
signal \N__56281\ : std_logic;
signal \N__56278\ : std_logic;
signal \N__56275\ : std_logic;
signal \N__56274\ : std_logic;
signal \N__56273\ : std_logic;
signal \N__56272\ : std_logic;
signal \N__56271\ : std_logic;
signal \N__56270\ : std_logic;
signal \N__56269\ : std_logic;
signal \N__56266\ : std_logic;
signal \N__56265\ : std_logic;
signal \N__56264\ : std_logic;
signal \N__56261\ : std_logic;
signal \N__56260\ : std_logic;
signal \N__56259\ : std_logic;
signal \N__56258\ : std_logic;
signal \N__56257\ : std_logic;
signal \N__56256\ : std_logic;
signal \N__56253\ : std_logic;
signal \N__56248\ : std_logic;
signal \N__56245\ : std_logic;
signal \N__56240\ : std_logic;
signal \N__56233\ : std_logic;
signal \N__56228\ : std_logic;
signal \N__56225\ : std_logic;
signal \N__56222\ : std_logic;
signal \N__56213\ : std_logic;
signal \N__56210\ : std_logic;
signal \N__56207\ : std_logic;
signal \N__56204\ : std_logic;
signal \N__56201\ : std_logic;
signal \N__56198\ : std_logic;
signal \N__56195\ : std_logic;
signal \N__56192\ : std_logic;
signal \N__56187\ : std_logic;
signal \N__56184\ : std_logic;
signal \N__56181\ : std_logic;
signal \N__56176\ : std_logic;
signal \N__56173\ : std_logic;
signal \N__56170\ : std_logic;
signal \N__56169\ : std_logic;
signal \N__56166\ : std_logic;
signal \N__56161\ : std_logic;
signal \N__56156\ : std_logic;
signal \N__56147\ : std_logic;
signal \N__56146\ : std_logic;
signal \N__56145\ : std_logic;
signal \N__56144\ : std_logic;
signal \N__56139\ : std_logic;
signal \N__56134\ : std_logic;
signal \N__56131\ : std_logic;
signal \N__56118\ : std_logic;
signal \N__56115\ : std_logic;
signal \N__56112\ : std_logic;
signal \N__56109\ : std_logic;
signal \N__56106\ : std_logic;
signal \N__56103\ : std_logic;
signal \N__56098\ : std_logic;
signal \N__56091\ : std_logic;
signal \N__56082\ : std_logic;
signal \N__56065\ : std_logic;
signal \N__56062\ : std_logic;
signal \N__56059\ : std_logic;
signal \N__56056\ : std_logic;
signal \N__56053\ : std_logic;
signal \N__56050\ : std_logic;
signal \N__56047\ : std_logic;
signal \N__56044\ : std_logic;
signal \N__56041\ : std_logic;
signal \N__56040\ : std_logic;
signal \N__56037\ : std_logic;
signal \N__56034\ : std_logic;
signal \N__56031\ : std_logic;
signal \N__56030\ : std_logic;
signal \N__56029\ : std_logic;
signal \N__56028\ : std_logic;
signal \N__56027\ : std_logic;
signal \N__56026\ : std_logic;
signal \N__56025\ : std_logic;
signal \N__56024\ : std_logic;
signal \N__56023\ : std_logic;
signal \N__56022\ : std_logic;
signal \N__56019\ : std_logic;
signal \N__56018\ : std_logic;
signal \N__56017\ : std_logic;
signal \N__56016\ : std_logic;
signal \N__56015\ : std_logic;
signal \N__55984\ : std_logic;
signal \N__55981\ : std_logic;
signal \N__55978\ : std_logic;
signal \N__55977\ : std_logic;
signal \N__55974\ : std_logic;
signal \N__55971\ : std_logic;
signal \N__55966\ : std_logic;
signal \N__55963\ : std_logic;
signal \N__55962\ : std_logic;
signal \N__55959\ : std_logic;
signal \N__55956\ : std_logic;
signal \N__55953\ : std_logic;
signal \N__55950\ : std_logic;
signal \N__55949\ : std_logic;
signal \N__55944\ : std_logic;
signal \N__55941\ : std_logic;
signal \N__55938\ : std_logic;
signal \N__55933\ : std_logic;
signal \N__55930\ : std_logic;
signal \N__55927\ : std_logic;
signal \N__55924\ : std_logic;
signal \N__55921\ : std_logic;
signal \N__55918\ : std_logic;
signal \N__55915\ : std_logic;
signal \N__55912\ : std_logic;
signal \N__55909\ : std_logic;
signal \N__55906\ : std_logic;
signal \N__55905\ : std_logic;
signal \N__55902\ : std_logic;
signal \N__55899\ : std_logic;
signal \N__55896\ : std_logic;
signal \N__55893\ : std_logic;
signal \N__55888\ : std_logic;
signal \N__55887\ : std_logic;
signal \N__55886\ : std_logic;
signal \N__55885\ : std_logic;
signal \N__55884\ : std_logic;
signal \N__55883\ : std_logic;
signal \N__55882\ : std_logic;
signal \N__55881\ : std_logic;
signal \N__55880\ : std_logic;
signal \N__55879\ : std_logic;
signal \N__55878\ : std_logic;
signal \N__55875\ : std_logic;
signal \N__55874\ : std_logic;
signal \N__55873\ : std_logic;
signal \N__55872\ : std_logic;
signal \N__55871\ : std_logic;
signal \N__55870\ : std_logic;
signal \N__55869\ : std_logic;
signal \N__55868\ : std_logic;
signal \N__55867\ : std_logic;
signal \N__55866\ : std_logic;
signal \N__55863\ : std_logic;
signal \N__55862\ : std_logic;
signal \N__55861\ : std_logic;
signal \N__55860\ : std_logic;
signal \N__55845\ : std_logic;
signal \N__55840\ : std_logic;
signal \N__55833\ : std_logic;
signal \N__55832\ : std_logic;
signal \N__55827\ : std_logic;
signal \N__55816\ : std_logic;
signal \N__55813\ : std_logic;
signal \N__55810\ : std_logic;
signal \N__55807\ : std_logic;
signal \N__55804\ : std_logic;
signal \N__55801\ : std_logic;
signal \N__55796\ : std_logic;
signal \N__55795\ : std_logic;
signal \N__55792\ : std_logic;
signal \N__55787\ : std_logic;
signal \N__55784\ : std_logic;
signal \N__55781\ : std_logic;
signal \N__55776\ : std_logic;
signal \N__55771\ : std_logic;
signal \N__55768\ : std_logic;
signal \N__55765\ : std_logic;
signal \N__55760\ : std_logic;
signal \N__55753\ : std_logic;
signal \N__55744\ : std_logic;
signal \N__55741\ : std_logic;
signal \N__55740\ : std_logic;
signal \N__55739\ : std_logic;
signal \N__55738\ : std_logic;
signal \N__55737\ : std_logic;
signal \N__55734\ : std_logic;
signal \N__55731\ : std_logic;
signal \N__55728\ : std_logic;
signal \N__55725\ : std_logic;
signal \N__55722\ : std_logic;
signal \N__55713\ : std_logic;
signal \N__55712\ : std_logic;
signal \N__55711\ : std_logic;
signal \N__55708\ : std_logic;
signal \N__55705\ : std_logic;
signal \N__55700\ : std_logic;
signal \N__55697\ : std_logic;
signal \N__55696\ : std_logic;
signal \N__55695\ : std_logic;
signal \N__55690\ : std_logic;
signal \N__55687\ : std_logic;
signal \N__55682\ : std_logic;
signal \N__55679\ : std_logic;
signal \N__55672\ : std_logic;
signal \N__55669\ : std_logic;
signal \N__55668\ : std_logic;
signal \N__55667\ : std_logic;
signal \N__55666\ : std_logic;
signal \N__55665\ : std_logic;
signal \N__55664\ : std_logic;
signal \N__55663\ : std_logic;
signal \N__55662\ : std_logic;
signal \N__55661\ : std_logic;
signal \N__55660\ : std_logic;
signal \N__55659\ : std_logic;
signal \N__55656\ : std_logic;
signal \N__55655\ : std_logic;
signal \N__55640\ : std_logic;
signal \N__55635\ : std_logic;
signal \N__55634\ : std_logic;
signal \N__55633\ : std_logic;
signal \N__55632\ : std_logic;
signal \N__55631\ : std_logic;
signal \N__55630\ : std_logic;
signal \N__55629\ : std_logic;
signal \N__55628\ : std_logic;
signal \N__55627\ : std_logic;
signal \N__55626\ : std_logic;
signal \N__55623\ : std_logic;
signal \N__55622\ : std_logic;
signal \N__55621\ : std_logic;
signal \N__55620\ : std_logic;
signal \N__55617\ : std_logic;
signal \N__55614\ : std_logic;
signal \N__55613\ : std_logic;
signal \N__55608\ : std_logic;
signal \N__55603\ : std_logic;
signal \N__55592\ : std_logic;
signal \N__55589\ : std_logic;
signal \N__55586\ : std_logic;
signal \N__55585\ : std_logic;
signal \N__55582\ : std_logic;
signal \N__55579\ : std_logic;
signal \N__55574\ : std_logic;
signal \N__55571\ : std_logic;
signal \N__55568\ : std_logic;
signal \N__55567\ : std_logic;
signal \N__55566\ : std_logic;
signal \N__55563\ : std_logic;
signal \N__55556\ : std_logic;
signal \N__55553\ : std_logic;
signal \N__55550\ : std_logic;
signal \N__55547\ : std_logic;
signal \N__55540\ : std_logic;
signal \N__55537\ : std_logic;
signal \N__55534\ : std_logic;
signal \N__55529\ : std_logic;
signal \N__55524\ : std_logic;
signal \N__55515\ : std_logic;
signal \N__55504\ : std_logic;
signal \N__55501\ : std_logic;
signal \N__55498\ : std_logic;
signal \N__55495\ : std_logic;
signal \N__55492\ : std_logic;
signal \N__55489\ : std_logic;
signal \N__55486\ : std_logic;
signal \N__55483\ : std_logic;
signal \N__55480\ : std_logic;
signal \N__55477\ : std_logic;
signal \N__55474\ : std_logic;
signal \N__55473\ : std_logic;
signal \N__55472\ : std_logic;
signal \N__55469\ : std_logic;
signal \N__55466\ : std_logic;
signal \N__55465\ : std_logic;
signal \N__55464\ : std_logic;
signal \N__55463\ : std_logic;
signal \N__55462\ : std_logic;
signal \N__55461\ : std_logic;
signal \N__55460\ : std_logic;
signal \N__55459\ : std_logic;
signal \N__55458\ : std_logic;
signal \N__55455\ : std_logic;
signal \N__55452\ : std_logic;
signal \N__55443\ : std_logic;
signal \N__55438\ : std_logic;
signal \N__55437\ : std_logic;
signal \N__55432\ : std_logic;
signal \N__55431\ : std_logic;
signal \N__55430\ : std_logic;
signal \N__55429\ : std_logic;
signal \N__55428\ : std_logic;
signal \N__55427\ : std_logic;
signal \N__55426\ : std_logic;
signal \N__55425\ : std_logic;
signal \N__55424\ : std_logic;
signal \N__55423\ : std_logic;
signal \N__55422\ : std_logic;
signal \N__55421\ : std_logic;
signal \N__55418\ : std_logic;
signal \N__55415\ : std_logic;
signal \N__55410\ : std_logic;
signal \N__55409\ : std_logic;
signal \N__55408\ : std_logic;
signal \N__55407\ : std_logic;
signal \N__55406\ : std_logic;
signal \N__55405\ : std_logic;
signal \N__55404\ : std_logic;
signal \N__55403\ : std_logic;
signal \N__55402\ : std_logic;
signal \N__55401\ : std_logic;
signal \N__55398\ : std_logic;
signal \N__55395\ : std_logic;
signal \N__55392\ : std_logic;
signal \N__55389\ : std_logic;
signal \N__55384\ : std_logic;
signal \N__55383\ : std_logic;
signal \N__55382\ : std_logic;
signal \N__55379\ : std_logic;
signal \N__55378\ : std_logic;
signal \N__55377\ : std_logic;
signal \N__55362\ : std_logic;
signal \N__55355\ : std_logic;
signal \N__55350\ : std_logic;
signal \N__55347\ : std_logic;
signal \N__55342\ : std_logic;
signal \N__55333\ : std_logic;
signal \N__55328\ : std_logic;
signal \N__55321\ : std_logic;
signal \N__55318\ : std_logic;
signal \N__55315\ : std_logic;
signal \N__55312\ : std_logic;
signal \N__55307\ : std_logic;
signal \N__55304\ : std_logic;
signal \N__55299\ : std_logic;
signal \N__55294\ : std_logic;
signal \N__55291\ : std_logic;
signal \N__55284\ : std_logic;
signal \N__55281\ : std_logic;
signal \N__55274\ : std_logic;
signal \N__55271\ : std_logic;
signal \N__55268\ : std_logic;
signal \N__55263\ : std_logic;
signal \N__55258\ : std_logic;
signal \N__55255\ : std_logic;
signal \N__55246\ : std_logic;
signal \N__55245\ : std_logic;
signal \N__55244\ : std_logic;
signal \N__55243\ : std_logic;
signal \N__55242\ : std_logic;
signal \N__55241\ : std_logic;
signal \N__55240\ : std_logic;
signal \N__55239\ : std_logic;
signal \N__55238\ : std_logic;
signal \N__55237\ : std_logic;
signal \N__55236\ : std_logic;
signal \N__55235\ : std_logic;
signal \N__55234\ : std_logic;
signal \N__55233\ : std_logic;
signal \N__55232\ : std_logic;
signal \N__55231\ : std_logic;
signal \N__55230\ : std_logic;
signal \N__55229\ : std_logic;
signal \N__55228\ : std_logic;
signal \N__55227\ : std_logic;
signal \N__55226\ : std_logic;
signal \N__55225\ : std_logic;
signal \N__55224\ : std_logic;
signal \N__55223\ : std_logic;
signal \N__55222\ : std_logic;
signal \N__55221\ : std_logic;
signal \N__55220\ : std_logic;
signal \N__55219\ : std_logic;
signal \N__55218\ : std_logic;
signal \N__55217\ : std_logic;
signal \N__55216\ : std_logic;
signal \N__55215\ : std_logic;
signal \N__55214\ : std_logic;
signal \N__55213\ : std_logic;
signal \N__55212\ : std_logic;
signal \N__55211\ : std_logic;
signal \N__55210\ : std_logic;
signal \N__55209\ : std_logic;
signal \N__55208\ : std_logic;
signal \N__55207\ : std_logic;
signal \N__55206\ : std_logic;
signal \N__55205\ : std_logic;
signal \N__55204\ : std_logic;
signal \N__55203\ : std_logic;
signal \N__55202\ : std_logic;
signal \N__55201\ : std_logic;
signal \N__55200\ : std_logic;
signal \N__55199\ : std_logic;
signal \N__55198\ : std_logic;
signal \N__55197\ : std_logic;
signal \N__55196\ : std_logic;
signal \N__55195\ : std_logic;
signal \N__55194\ : std_logic;
signal \N__55193\ : std_logic;
signal \N__55192\ : std_logic;
signal \N__55191\ : std_logic;
signal \N__55190\ : std_logic;
signal \N__55189\ : std_logic;
signal \N__55188\ : std_logic;
signal \N__55187\ : std_logic;
signal \N__55186\ : std_logic;
signal \N__55185\ : std_logic;
signal \N__55184\ : std_logic;
signal \N__55183\ : std_logic;
signal \N__55182\ : std_logic;
signal \N__55181\ : std_logic;
signal \N__55180\ : std_logic;
signal \N__55179\ : std_logic;
signal \N__55178\ : std_logic;
signal \N__55177\ : std_logic;
signal \N__55176\ : std_logic;
signal \N__55175\ : std_logic;
signal \N__55174\ : std_logic;
signal \N__55173\ : std_logic;
signal \N__55172\ : std_logic;
signal \N__55171\ : std_logic;
signal \N__55170\ : std_logic;
signal \N__55169\ : std_logic;
signal \N__55168\ : std_logic;
signal \N__55167\ : std_logic;
signal \N__55166\ : std_logic;
signal \N__55165\ : std_logic;
signal \N__55164\ : std_logic;
signal \N__55163\ : std_logic;
signal \N__55162\ : std_logic;
signal \N__55161\ : std_logic;
signal \N__55160\ : std_logic;
signal \N__55159\ : std_logic;
signal \N__55158\ : std_logic;
signal \N__55157\ : std_logic;
signal \N__55156\ : std_logic;
signal \N__55155\ : std_logic;
signal \N__55154\ : std_logic;
signal \N__55153\ : std_logic;
signal \N__55152\ : std_logic;
signal \N__55151\ : std_logic;
signal \N__55150\ : std_logic;
signal \N__55149\ : std_logic;
signal \N__55148\ : std_logic;
signal \N__55147\ : std_logic;
signal \N__55146\ : std_logic;
signal \N__55145\ : std_logic;
signal \N__55144\ : std_logic;
signal \N__55143\ : std_logic;
signal \N__55142\ : std_logic;
signal \N__55141\ : std_logic;
signal \N__55140\ : std_logic;
signal \N__55139\ : std_logic;
signal \N__55138\ : std_logic;
signal \N__55137\ : std_logic;
signal \N__55136\ : std_logic;
signal \N__55135\ : std_logic;
signal \N__55134\ : std_logic;
signal \N__55133\ : std_logic;
signal \N__55132\ : std_logic;
signal \N__55131\ : std_logic;
signal \N__55130\ : std_logic;
signal \N__55129\ : std_logic;
signal \N__55128\ : std_logic;
signal \N__55127\ : std_logic;
signal \N__55126\ : std_logic;
signal \N__55125\ : std_logic;
signal \N__55124\ : std_logic;
signal \N__55123\ : std_logic;
signal \N__55122\ : std_logic;
signal \N__55121\ : std_logic;
signal \N__55120\ : std_logic;
signal \N__55119\ : std_logic;
signal \N__55118\ : std_logic;
signal \N__55117\ : std_logic;
signal \N__55116\ : std_logic;
signal \N__55115\ : std_logic;
signal \N__55114\ : std_logic;
signal \N__55113\ : std_logic;
signal \N__55112\ : std_logic;
signal \N__55111\ : std_logic;
signal \N__55110\ : std_logic;
signal \N__55109\ : std_logic;
signal \N__55108\ : std_logic;
signal \N__55107\ : std_logic;
signal \N__55106\ : std_logic;
signal \N__55105\ : std_logic;
signal \N__55104\ : std_logic;
signal \N__55103\ : std_logic;
signal \N__55102\ : std_logic;
signal \N__55101\ : std_logic;
signal \N__55100\ : std_logic;
signal \N__55099\ : std_logic;
signal \N__55098\ : std_logic;
signal \N__55097\ : std_logic;
signal \N__55096\ : std_logic;
signal \N__55095\ : std_logic;
signal \N__55094\ : std_logic;
signal \N__55093\ : std_logic;
signal \N__55092\ : std_logic;
signal \N__55091\ : std_logic;
signal \N__55090\ : std_logic;
signal \N__55089\ : std_logic;
signal \N__55088\ : std_logic;
signal \N__55087\ : std_logic;
signal \N__55086\ : std_logic;
signal \N__55085\ : std_logic;
signal \N__55084\ : std_logic;
signal \N__55083\ : std_logic;
signal \N__55082\ : std_logic;
signal \N__55081\ : std_logic;
signal \N__55080\ : std_logic;
signal \N__55079\ : std_logic;
signal \N__55078\ : std_logic;
signal \N__55077\ : std_logic;
signal \N__55076\ : std_logic;
signal \N__55075\ : std_logic;
signal \N__55074\ : std_logic;
signal \N__54727\ : std_logic;
signal \N__54724\ : std_logic;
signal \N__54723\ : std_logic;
signal \N__54722\ : std_logic;
signal \N__54721\ : std_logic;
signal \N__54720\ : std_logic;
signal \N__54719\ : std_logic;
signal \N__54718\ : std_logic;
signal \N__54717\ : std_logic;
signal \N__54716\ : std_logic;
signal \N__54715\ : std_logic;
signal \N__54714\ : std_logic;
signal \N__54713\ : std_logic;
signal \N__54712\ : std_logic;
signal \N__54711\ : std_logic;
signal \N__54710\ : std_logic;
signal \N__54709\ : std_logic;
signal \N__54706\ : std_logic;
signal \N__54705\ : std_logic;
signal \N__54704\ : std_logic;
signal \N__54703\ : std_logic;
signal \N__54702\ : std_logic;
signal \N__54701\ : std_logic;
signal \N__54700\ : std_logic;
signal \N__54699\ : std_logic;
signal \N__54696\ : std_logic;
signal \N__54695\ : std_logic;
signal \N__54694\ : std_logic;
signal \N__54693\ : std_logic;
signal \N__54690\ : std_logic;
signal \N__54687\ : std_logic;
signal \N__54684\ : std_logic;
signal \N__54681\ : std_logic;
signal \N__54676\ : std_logic;
signal \N__54675\ : std_logic;
signal \N__54674\ : std_logic;
signal \N__54673\ : std_logic;
signal \N__54672\ : std_logic;
signal \N__54671\ : std_logic;
signal \N__54670\ : std_logic;
signal \N__54669\ : std_logic;
signal \N__54668\ : std_logic;
signal \N__54667\ : std_logic;
signal \N__54666\ : std_logic;
signal \N__54665\ : std_logic;
signal \N__54664\ : std_logic;
signal \N__54663\ : std_logic;
signal \N__54662\ : std_logic;
signal \N__54661\ : std_logic;
signal \N__54660\ : std_logic;
signal \N__54659\ : std_logic;
signal \N__54658\ : std_logic;
signal \N__54657\ : std_logic;
signal \N__54656\ : std_logic;
signal \N__54653\ : std_logic;
signal \N__54650\ : std_logic;
signal \N__54649\ : std_logic;
signal \N__54646\ : std_logic;
signal \N__54645\ : std_logic;
signal \N__54642\ : std_logic;
signal \N__54639\ : std_logic;
signal \N__54636\ : std_logic;
signal \N__54635\ : std_logic;
signal \N__54632\ : std_logic;
signal \N__54629\ : std_logic;
signal \N__54626\ : std_logic;
signal \N__54625\ : std_logic;
signal \N__54624\ : std_logic;
signal \N__54623\ : std_logic;
signal \N__54620\ : std_logic;
signal \N__54617\ : std_logic;
signal \N__54612\ : std_logic;
signal \N__54611\ : std_logic;
signal \N__54610\ : std_logic;
signal \N__54609\ : std_logic;
signal \N__54604\ : std_logic;
signal \N__54601\ : std_logic;
signal \N__54600\ : std_logic;
signal \N__54599\ : std_logic;
signal \N__54598\ : std_logic;
signal \N__54597\ : std_logic;
signal \N__54596\ : std_logic;
signal \N__54593\ : std_logic;
signal \N__54592\ : std_logic;
signal \N__54591\ : std_logic;
signal \N__54590\ : std_logic;
signal \N__54589\ : std_logic;
signal \N__54588\ : std_logic;
signal \N__54585\ : std_logic;
signal \N__54584\ : std_logic;
signal \N__54581\ : std_logic;
signal \N__54580\ : std_logic;
signal \N__54577\ : std_logic;
signal \N__54576\ : std_logic;
signal \N__54571\ : std_logic;
signal \N__54564\ : std_logic;
signal \N__54563\ : std_logic;
signal \N__54562\ : std_logic;
signal \N__54561\ : std_logic;
signal \N__54558\ : std_logic;
signal \N__54555\ : std_logic;
signal \N__54550\ : std_logic;
signal \N__54545\ : std_logic;
signal \N__54544\ : std_logic;
signal \N__54541\ : std_logic;
signal \N__54538\ : std_logic;
signal \N__54537\ : std_logic;
signal \N__54536\ : std_logic;
signal \N__54535\ : std_logic;
signal \N__54522\ : std_logic;
signal \N__54511\ : std_logic;
signal \N__54508\ : std_logic;
signal \N__54495\ : std_logic;
signal \N__54490\ : std_logic;
signal \N__54489\ : std_logic;
signal \N__54488\ : std_logic;
signal \N__54487\ : std_logic;
signal \N__54486\ : std_logic;
signal \N__54485\ : std_logic;
signal \N__54482\ : std_logic;
signal \N__54475\ : std_logic;
signal \N__54472\ : std_logic;
signal \N__54467\ : std_logic;
signal \N__54460\ : std_logic;
signal \N__54455\ : std_logic;
signal \N__54452\ : std_logic;
signal \N__54451\ : std_logic;
signal \N__54448\ : std_logic;
signal \N__54445\ : std_logic;
signal \N__54442\ : std_logic;
signal \N__54441\ : std_logic;
signal \N__54440\ : std_logic;
signal \N__54437\ : std_logic;
signal \N__54434\ : std_logic;
signal \N__54433\ : std_logic;
signal \N__54430\ : std_logic;
signal \N__54427\ : std_logic;
signal \N__54424\ : std_logic;
signal \N__54421\ : std_logic;
signal \N__54416\ : std_logic;
signal \N__54399\ : std_logic;
signal \N__54394\ : std_logic;
signal \N__54389\ : std_logic;
signal \N__54388\ : std_logic;
signal \N__54387\ : std_logic;
signal \N__54384\ : std_logic;
signal \N__54381\ : std_logic;
signal \N__54376\ : std_logic;
signal \N__54373\ : std_logic;
signal \N__54372\ : std_logic;
signal \N__54369\ : std_logic;
signal \N__54368\ : std_logic;
signal \N__54367\ : std_logic;
signal \N__54364\ : std_logic;
signal \N__54361\ : std_logic;
signal \N__54358\ : std_logic;
signal \N__54355\ : std_logic;
signal \N__54352\ : std_logic;
signal \N__54341\ : std_logic;
signal \N__54336\ : std_logic;
signal \N__54329\ : std_logic;
signal \N__54318\ : std_logic;
signal \N__54315\ : std_logic;
signal \N__54312\ : std_logic;
signal \N__54309\ : std_logic;
signal \N__54306\ : std_logic;
signal \N__54301\ : std_logic;
signal \N__54298\ : std_logic;
signal \N__54295\ : std_logic;
signal \N__54288\ : std_logic;
signal \N__54285\ : std_logic;
signal \N__54280\ : std_logic;
signal \N__54275\ : std_logic;
signal \N__54268\ : std_logic;
signal \N__54263\ : std_logic;
signal \N__54260\ : std_logic;
signal \N__54253\ : std_logic;
signal \N__54250\ : std_logic;
signal \N__54249\ : std_logic;
signal \N__54246\ : std_logic;
signal \N__54245\ : std_logic;
signal \N__54244\ : std_logic;
signal \N__54241\ : std_logic;
signal \N__54240\ : std_logic;
signal \N__54239\ : std_logic;
signal \N__54238\ : std_logic;
signal \N__54235\ : std_logic;
signal \N__54228\ : std_logic;
signal \N__54223\ : std_logic;
signal \N__54220\ : std_logic;
signal \N__54211\ : std_logic;
signal \N__54200\ : std_logic;
signal \N__54193\ : std_logic;
signal \N__54184\ : std_logic;
signal \N__54177\ : std_logic;
signal \N__54176\ : std_logic;
signal \N__54175\ : std_logic;
signal \N__54172\ : std_logic;
signal \N__54169\ : std_logic;
signal \N__54166\ : std_logic;
signal \N__54157\ : std_logic;
signal \N__54154\ : std_logic;
signal \N__54143\ : std_logic;
signal \N__54138\ : std_logic;
signal \N__54135\ : std_logic;
signal \N__54132\ : std_logic;
signal \N__54127\ : std_logic;
signal \N__54106\ : std_logic;
signal \N__54105\ : std_logic;
signal \N__54104\ : std_logic;
signal \N__54103\ : std_logic;
signal \N__54102\ : std_logic;
signal \N__54101\ : std_logic;
signal \N__54100\ : std_logic;
signal \N__54099\ : std_logic;
signal \N__54098\ : std_logic;
signal \N__54097\ : std_logic;
signal \N__54096\ : std_logic;
signal \N__54095\ : std_logic;
signal \N__54094\ : std_logic;
signal \N__54093\ : std_logic;
signal \N__54092\ : std_logic;
signal \N__54091\ : std_logic;
signal \N__54090\ : std_logic;
signal \N__54089\ : std_logic;
signal \N__54088\ : std_logic;
signal \N__54087\ : std_logic;
signal \N__54086\ : std_logic;
signal \N__54085\ : std_logic;
signal \N__54084\ : std_logic;
signal \N__54083\ : std_logic;
signal \N__54082\ : std_logic;
signal \N__54081\ : std_logic;
signal \N__54080\ : std_logic;
signal \N__54079\ : std_logic;
signal \N__54076\ : std_logic;
signal \N__54067\ : std_logic;
signal \N__54064\ : std_logic;
signal \N__54061\ : std_logic;
signal \N__54052\ : std_logic;
signal \N__54051\ : std_logic;
signal \N__54048\ : std_logic;
signal \N__54045\ : std_logic;
signal \N__54042\ : std_logic;
signal \N__54039\ : std_logic;
signal \N__54036\ : std_logic;
signal \N__54035\ : std_logic;
signal \N__54034\ : std_logic;
signal \N__54033\ : std_logic;
signal \N__54032\ : std_logic;
signal \N__54031\ : std_logic;
signal \N__54028\ : std_logic;
signal \N__54027\ : std_logic;
signal \N__54010\ : std_logic;
signal \N__54005\ : std_logic;
signal \N__54002\ : std_logic;
signal \N__54001\ : std_logic;
signal \N__54000\ : std_logic;
signal \N__53997\ : std_logic;
signal \N__53988\ : std_logic;
signal \N__53987\ : std_logic;
signal \N__53986\ : std_logic;
signal \N__53985\ : std_logic;
signal \N__53984\ : std_logic;
signal \N__53983\ : std_logic;
signal \N__53982\ : std_logic;
signal \N__53981\ : std_logic;
signal \N__53980\ : std_logic;
signal \N__53979\ : std_logic;
signal \N__53978\ : std_logic;
signal \N__53977\ : std_logic;
signal \N__53976\ : std_logic;
signal \N__53975\ : std_logic;
signal \N__53972\ : std_logic;
signal \N__53967\ : std_logic;
signal \N__53964\ : std_logic;
signal \N__53961\ : std_logic;
signal \N__53958\ : std_logic;
signal \N__53957\ : std_logic;
signal \N__53956\ : std_logic;
signal \N__53953\ : std_logic;
signal \N__53950\ : std_logic;
signal \N__53949\ : std_logic;
signal \N__53948\ : std_logic;
signal \N__53947\ : std_logic;
signal \N__53946\ : std_logic;
signal \N__53945\ : std_logic;
signal \N__53944\ : std_logic;
signal \N__53943\ : std_logic;
signal \N__53942\ : std_logic;
signal \N__53941\ : std_logic;
signal \N__53940\ : std_logic;
signal \N__53939\ : std_logic;
signal \N__53938\ : std_logic;
signal \N__53937\ : std_logic;
signal \N__53936\ : std_logic;
signal \N__53935\ : std_logic;
signal \N__53932\ : std_logic;
signal \N__53929\ : std_logic;
signal \N__53926\ : std_logic;
signal \N__53923\ : std_logic;
signal \N__53920\ : std_logic;
signal \N__53913\ : std_logic;
signal \N__53910\ : std_logic;
signal \N__53909\ : std_logic;
signal \N__53908\ : std_logic;
signal \N__53905\ : std_logic;
signal \N__53904\ : std_logic;
signal \N__53903\ : std_logic;
signal \N__53902\ : std_logic;
signal \N__53901\ : std_logic;
signal \N__53900\ : std_logic;
signal \N__53895\ : std_logic;
signal \N__53892\ : std_logic;
signal \N__53889\ : std_logic;
signal \N__53886\ : std_logic;
signal \N__53885\ : std_logic;
signal \N__53884\ : std_logic;
signal \N__53883\ : std_logic;
signal \N__53882\ : std_logic;
signal \N__53881\ : std_logic;
signal \N__53878\ : std_logic;
signal \N__53875\ : std_logic;
signal \N__53874\ : std_logic;
signal \N__53873\ : std_logic;
signal \N__53872\ : std_logic;
signal \N__53871\ : std_logic;
signal \N__53854\ : std_logic;
signal \N__53851\ : std_logic;
signal \N__53848\ : std_logic;
signal \N__53843\ : std_logic;
signal \N__53840\ : std_logic;
signal \N__53839\ : std_logic;
signal \N__53838\ : std_logic;
signal \N__53837\ : std_logic;
signal \N__53834\ : std_logic;
signal \N__53831\ : std_logic;
signal \N__53830\ : std_logic;
signal \N__53829\ : std_logic;
signal \N__53828\ : std_logic;
signal \N__53823\ : std_logic;
signal \N__53806\ : std_logic;
signal \N__53791\ : std_logic;
signal \N__53780\ : std_logic;
signal \N__53777\ : std_logic;
signal \N__53774\ : std_logic;
signal \N__53771\ : std_logic;
signal \N__53768\ : std_logic;
signal \N__53765\ : std_logic;
signal \N__53756\ : std_logic;
signal \N__53753\ : std_logic;
signal \N__53750\ : std_logic;
signal \N__53743\ : std_logic;
signal \N__53742\ : std_logic;
signal \N__53741\ : std_logic;
signal \N__53740\ : std_logic;
signal \N__53733\ : std_logic;
signal \N__53728\ : std_logic;
signal \N__53723\ : std_logic;
signal \N__53720\ : std_logic;
signal \N__53713\ : std_logic;
signal \N__53704\ : std_logic;
signal \N__53701\ : std_logic;
signal \N__53696\ : std_logic;
signal \N__53693\ : std_logic;
signal \N__53688\ : std_logic;
signal \N__53687\ : std_logic;
signal \N__53686\ : std_logic;
signal \N__53685\ : std_logic;
signal \N__53682\ : std_logic;
signal \N__53681\ : std_logic;
signal \N__53680\ : std_logic;
signal \N__53679\ : std_logic;
signal \N__53676\ : std_logic;
signal \N__53673\ : std_logic;
signal \N__53670\ : std_logic;
signal \N__53659\ : std_logic;
signal \N__53658\ : std_logic;
signal \N__53657\ : std_logic;
signal \N__53656\ : std_logic;
signal \N__53655\ : std_logic;
signal \N__53654\ : std_logic;
signal \N__53645\ : std_logic;
signal \N__53638\ : std_logic;
signal \N__53637\ : std_logic;
signal \N__53630\ : std_logic;
signal \N__53623\ : std_logic;
signal \N__53608\ : std_logic;
signal \N__53601\ : std_logic;
signal \N__53592\ : std_logic;
signal \N__53587\ : std_logic;
signal \N__53582\ : std_logic;
signal \N__53571\ : std_logic;
signal \N__53568\ : std_logic;
signal \N__53565\ : std_logic;
signal \N__53562\ : std_logic;
signal \N__53555\ : std_logic;
signal \N__53536\ : std_logic;
signal \N__53533\ : std_logic;
signal \N__53532\ : std_logic;
signal \N__53531\ : std_logic;
signal \N__53530\ : std_logic;
signal \N__53529\ : std_logic;
signal \N__53526\ : std_logic;
signal \N__53523\ : std_logic;
signal \N__53522\ : std_logic;
signal \N__53521\ : std_logic;
signal \N__53518\ : std_logic;
signal \N__53513\ : std_logic;
signal \N__53512\ : std_logic;
signal \N__53511\ : std_logic;
signal \N__53510\ : std_logic;
signal \N__53509\ : std_logic;
signal \N__53506\ : std_logic;
signal \N__53503\ : std_logic;
signal \N__53500\ : std_logic;
signal \N__53499\ : std_logic;
signal \N__53498\ : std_logic;
signal \N__53497\ : std_logic;
signal \N__53496\ : std_logic;
signal \N__53495\ : std_logic;
signal \N__53494\ : std_logic;
signal \N__53493\ : std_logic;
signal \N__53492\ : std_logic;
signal \N__53491\ : std_logic;
signal \N__53490\ : std_logic;
signal \N__53489\ : std_logic;
signal \N__53488\ : std_logic;
signal \N__53487\ : std_logic;
signal \N__53486\ : std_logic;
signal \N__53485\ : std_logic;
signal \N__53482\ : std_logic;
signal \N__53479\ : std_logic;
signal \N__53476\ : std_logic;
signal \N__53475\ : std_logic;
signal \N__53474\ : std_logic;
signal \N__53467\ : std_logic;
signal \N__53466\ : std_logic;
signal \N__53463\ : std_logic;
signal \N__53462\ : std_logic;
signal \N__53461\ : std_logic;
signal \N__53454\ : std_logic;
signal \N__53451\ : std_logic;
signal \N__53450\ : std_logic;
signal \N__53449\ : std_logic;
signal \N__53448\ : std_logic;
signal \N__53439\ : std_logic;
signal \N__53438\ : std_logic;
signal \N__53437\ : std_logic;
signal \N__53432\ : std_logic;
signal \N__53421\ : std_logic;
signal \N__53418\ : std_logic;
signal \N__53417\ : std_logic;
signal \N__53414\ : std_logic;
signal \N__53411\ : std_logic;
signal \N__53408\ : std_logic;
signal \N__53403\ : std_logic;
signal \N__53398\ : std_logic;
signal \N__53395\ : std_logic;
signal \N__53392\ : std_logic;
signal \N__53389\ : std_logic;
signal \N__53384\ : std_logic;
signal \N__53379\ : std_logic;
signal \N__53372\ : std_logic;
signal \N__53371\ : std_logic;
signal \N__53368\ : std_logic;
signal \N__53365\ : std_logic;
signal \N__53362\ : std_logic;
signal \N__53361\ : std_logic;
signal \N__53358\ : std_logic;
signal \N__53353\ : std_logic;
signal \N__53350\ : std_logic;
signal \N__53345\ : std_logic;
signal \N__53340\ : std_logic;
signal \N__53337\ : std_logic;
signal \N__53332\ : std_logic;
signal \N__53327\ : std_logic;
signal \N__53324\ : std_logic;
signal \N__53321\ : std_logic;
signal \N__53318\ : std_logic;
signal \N__53311\ : std_logic;
signal \N__53308\ : std_logic;
signal \N__53303\ : std_logic;
signal \N__53300\ : std_logic;
signal \N__53291\ : std_logic;
signal \N__53288\ : std_logic;
signal \N__53285\ : std_logic;
signal \N__53266\ : std_logic;
signal \N__53263\ : std_logic;
signal \N__53260\ : std_logic;
signal \N__53259\ : std_logic;
signal \N__53258\ : std_logic;
signal \N__53255\ : std_logic;
signal \N__53250\ : std_logic;
signal \N__53247\ : std_logic;
signal \N__53244\ : std_logic;
signal \N__53239\ : std_logic;
signal \N__53236\ : std_logic;
signal \N__53233\ : std_logic;
signal \N__53230\ : std_logic;
signal \N__53229\ : std_logic;
signal \N__53228\ : std_logic;
signal \N__53225\ : std_logic;
signal \N__53222\ : std_logic;
signal \N__53219\ : std_logic;
signal \N__53212\ : std_logic;
signal \N__53209\ : std_logic;
signal \N__53206\ : std_logic;
signal \N__53203\ : std_logic;
signal \N__53200\ : std_logic;
signal \N__53199\ : std_logic;
signal \N__53194\ : std_logic;
signal \N__53193\ : std_logic;
signal \N__53190\ : std_logic;
signal \N__53187\ : std_logic;
signal \N__53184\ : std_logic;
signal \N__53181\ : std_logic;
signal \N__53176\ : std_logic;
signal \N__53173\ : std_logic;
signal \N__53170\ : std_logic;
signal \N__53167\ : std_logic;
signal \N__53164\ : std_logic;
signal \N__53161\ : std_logic;
signal \N__53160\ : std_logic;
signal \N__53157\ : std_logic;
signal \N__53154\ : std_logic;
signal \N__53149\ : std_logic;
signal \N__53148\ : std_logic;
signal \N__53145\ : std_logic;
signal \N__53142\ : std_logic;
signal \N__53139\ : std_logic;
signal \N__53136\ : std_logic;
signal \N__53131\ : std_logic;
signal \N__53128\ : std_logic;
signal \N__53125\ : std_logic;
signal \N__53122\ : std_logic;
signal \N__53119\ : std_logic;
signal \N__53116\ : std_logic;
signal \N__53113\ : std_logic;
signal \N__53110\ : std_logic;
signal \N__53107\ : std_logic;
signal \N__53104\ : std_logic;
signal \N__53103\ : std_logic;
signal \N__53100\ : std_logic;
signal \N__53097\ : std_logic;
signal \N__53094\ : std_logic;
signal \N__53089\ : std_logic;
signal \N__53088\ : std_logic;
signal \N__53085\ : std_logic;
signal \N__53082\ : std_logic;
signal \N__53079\ : std_logic;
signal \N__53074\ : std_logic;
signal \N__53071\ : std_logic;
signal \N__53068\ : std_logic;
signal \N__53067\ : std_logic;
signal \N__53064\ : std_logic;
signal \N__53061\ : std_logic;
signal \N__53058\ : std_logic;
signal \N__53053\ : std_logic;
signal \N__53052\ : std_logic;
signal \N__53049\ : std_logic;
signal \N__53046\ : std_logic;
signal \N__53043\ : std_logic;
signal \N__53038\ : std_logic;
signal \N__53035\ : std_logic;
signal \N__53032\ : std_logic;
signal \N__53029\ : std_logic;
signal \N__53026\ : std_logic;
signal \N__53025\ : std_logic;
signal \N__53022\ : std_logic;
signal \N__53019\ : std_logic;
signal \N__53018\ : std_logic;
signal \N__53015\ : std_logic;
signal \N__53012\ : std_logic;
signal \N__53009\ : std_logic;
signal \N__53006\ : std_logic;
signal \N__53005\ : std_logic;
signal \N__53002\ : std_logic;
signal \N__52999\ : std_logic;
signal \N__52996\ : std_logic;
signal \N__52993\ : std_logic;
signal \N__52990\ : std_logic;
signal \N__52985\ : std_logic;
signal \N__52982\ : std_logic;
signal \N__52979\ : std_logic;
signal \N__52976\ : std_logic;
signal \N__52969\ : std_logic;
signal \N__52966\ : std_logic;
signal \N__52963\ : std_logic;
signal \N__52960\ : std_logic;
signal \N__52957\ : std_logic;
signal \N__52954\ : std_logic;
signal \N__52953\ : std_logic;
signal \N__52952\ : std_logic;
signal \N__52949\ : std_logic;
signal \N__52946\ : std_logic;
signal \N__52943\ : std_logic;
signal \N__52942\ : std_logic;
signal \N__52941\ : std_logic;
signal \N__52938\ : std_logic;
signal \N__52933\ : std_logic;
signal \N__52930\ : std_logic;
signal \N__52927\ : std_logic;
signal \N__52924\ : std_logic;
signal \N__52917\ : std_logic;
signal \N__52914\ : std_logic;
signal \N__52911\ : std_logic;
signal \N__52906\ : std_logic;
signal \N__52903\ : std_logic;
signal \N__52900\ : std_logic;
signal \N__52897\ : std_logic;
signal \N__52894\ : std_logic;
signal \N__52891\ : std_logic;
signal \N__52888\ : std_logic;
signal \N__52887\ : std_logic;
signal \N__52886\ : std_logic;
signal \N__52883\ : std_logic;
signal \N__52880\ : std_logic;
signal \N__52879\ : std_logic;
signal \N__52878\ : std_logic;
signal \N__52877\ : std_logic;
signal \N__52874\ : std_logic;
signal \N__52873\ : std_logic;
signal \N__52868\ : std_logic;
signal \N__52865\ : std_logic;
signal \N__52862\ : std_logic;
signal \N__52861\ : std_logic;
signal \N__52860\ : std_logic;
signal \N__52857\ : std_logic;
signal \N__52854\ : std_logic;
signal \N__52851\ : std_logic;
signal \N__52844\ : std_logic;
signal \N__52841\ : std_logic;
signal \N__52838\ : std_logic;
signal \N__52837\ : std_logic;
signal \N__52836\ : std_logic;
signal \N__52835\ : std_logic;
signal \N__52832\ : std_logic;
signal \N__52831\ : std_logic;
signal \N__52830\ : std_logic;
signal \N__52829\ : std_logic;
signal \N__52828\ : std_logic;
signal \N__52823\ : std_logic;
signal \N__52816\ : std_logic;
signal \N__52813\ : std_logic;
signal \N__52812\ : std_logic;
signal \N__52811\ : std_logic;
signal \N__52810\ : std_logic;
signal \N__52809\ : std_logic;
signal \N__52806\ : std_logic;
signal \N__52805\ : std_logic;
signal \N__52804\ : std_logic;
signal \N__52803\ : std_logic;
signal \N__52802\ : std_logic;
signal \N__52801\ : std_logic;
signal \N__52800\ : std_logic;
signal \N__52799\ : std_logic;
signal \N__52796\ : std_logic;
signal \N__52795\ : std_logic;
signal \N__52794\ : std_logic;
signal \N__52793\ : std_logic;
signal \N__52792\ : std_logic;
signal \N__52791\ : std_logic;
signal \N__52788\ : std_logic;
signal \N__52785\ : std_logic;
signal \N__52784\ : std_logic;
signal \N__52781\ : std_logic;
signal \N__52780\ : std_logic;
signal \N__52777\ : std_logic;
signal \N__52776\ : std_logic;
signal \N__52773\ : std_logic;
signal \N__52766\ : std_logic;
signal \N__52763\ : std_logic;
signal \N__52762\ : std_logic;
signal \N__52759\ : std_logic;
signal \N__52758\ : std_logic;
signal \N__52755\ : std_logic;
signal \N__52754\ : std_logic;
signal \N__52751\ : std_logic;
signal \N__52750\ : std_logic;
signal \N__52749\ : std_logic;
signal \N__52748\ : std_logic;
signal \N__52747\ : std_logic;
signal \N__52744\ : std_logic;
signal \N__52737\ : std_logic;
signal \N__52728\ : std_logic;
signal \N__52725\ : std_logic;
signal \N__52724\ : std_logic;
signal \N__52723\ : std_logic;
signal \N__52720\ : std_logic;
signal \N__52719\ : std_logic;
signal \N__52716\ : std_logic;
signal \N__52715\ : std_logic;
signal \N__52712\ : std_logic;
signal \N__52711\ : std_logic;
signal \N__52708\ : std_logic;
signal \N__52707\ : std_logic;
signal \N__52704\ : std_logic;
signal \N__52701\ : std_logic;
signal \N__52686\ : std_logic;
signal \N__52683\ : std_logic;
signal \N__52668\ : std_logic;
signal \N__52667\ : std_logic;
signal \N__52664\ : std_logic;
signal \N__52663\ : std_logic;
signal \N__52660\ : std_logic;
signal \N__52659\ : std_logic;
signal \N__52656\ : std_logic;
signal \N__52655\ : std_logic;
signal \N__52652\ : std_logic;
signal \N__52649\ : std_logic;
signal \N__52644\ : std_logic;
signal \N__52641\ : std_logic;
signal \N__52638\ : std_logic;
signal \N__52635\ : std_logic;
signal \N__52632\ : std_logic;
signal \N__52615\ : std_logic;
signal \N__52610\ : std_logic;
signal \N__52605\ : std_logic;
signal \N__52588\ : std_logic;
signal \N__52585\ : std_logic;
signal \N__52582\ : std_logic;
signal \N__52577\ : std_logic;
signal \N__52574\ : std_logic;
signal \N__52571\ : std_logic;
signal \N__52568\ : std_logic;
signal \N__52561\ : std_logic;
signal \N__52556\ : std_logic;
signal \N__52551\ : std_logic;
signal \N__52546\ : std_logic;
signal \N__52543\ : std_logic;
signal \N__52534\ : std_logic;
signal \N__52531\ : std_logic;
signal \N__52528\ : std_logic;
signal \N__52525\ : std_logic;
signal \N__52522\ : std_logic;
signal \N__52519\ : std_logic;
signal \N__52518\ : std_logic;
signal \N__52515\ : std_logic;
signal \N__52512\ : std_logic;
signal \N__52507\ : std_logic;
signal \N__52504\ : std_logic;
signal \N__52501\ : std_logic;
signal \N__52498\ : std_logic;
signal \N__52497\ : std_logic;
signal \N__52494\ : std_logic;
signal \N__52491\ : std_logic;
signal \N__52486\ : std_logic;
signal \N__52483\ : std_logic;
signal \N__52482\ : std_logic;
signal \N__52479\ : std_logic;
signal \N__52476\ : std_logic;
signal \N__52471\ : std_logic;
signal \N__52468\ : std_logic;
signal \N__52465\ : std_logic;
signal \N__52462\ : std_logic;
signal \N__52461\ : std_logic;
signal \N__52458\ : std_logic;
signal \N__52455\ : std_logic;
signal \N__52452\ : std_logic;
signal \N__52449\ : std_logic;
signal \N__52444\ : std_logic;
signal \N__52443\ : std_logic;
signal \N__52442\ : std_logic;
signal \N__52441\ : std_logic;
signal \N__52438\ : std_logic;
signal \N__52437\ : std_logic;
signal \N__52434\ : std_logic;
signal \N__52431\ : std_logic;
signal \N__52430\ : std_logic;
signal \N__52427\ : std_logic;
signal \N__52426\ : std_logic;
signal \N__52425\ : std_logic;
signal \N__52424\ : std_logic;
signal \N__52421\ : std_logic;
signal \N__52418\ : std_logic;
signal \N__52417\ : std_logic;
signal \N__52416\ : std_logic;
signal \N__52415\ : std_logic;
signal \N__52414\ : std_logic;
signal \N__52413\ : std_logic;
signal \N__52408\ : std_logic;
signal \N__52407\ : std_logic;
signal \N__52404\ : std_logic;
signal \N__52401\ : std_logic;
signal \N__52398\ : std_logic;
signal \N__52395\ : std_logic;
signal \N__52392\ : std_logic;
signal \N__52391\ : std_logic;
signal \N__52386\ : std_logic;
signal \N__52383\ : std_logic;
signal \N__52380\ : std_logic;
signal \N__52379\ : std_logic;
signal \N__52376\ : std_logic;
signal \N__52375\ : std_logic;
signal \N__52372\ : std_logic;
signal \N__52369\ : std_logic;
signal \N__52368\ : std_logic;
signal \N__52365\ : std_logic;
signal \N__52364\ : std_logic;
signal \N__52361\ : std_logic;
signal \N__52360\ : std_logic;
signal \N__52353\ : std_logic;
signal \N__52348\ : std_logic;
signal \N__52345\ : std_logic;
signal \N__52340\ : std_logic;
signal \N__52337\ : std_logic;
signal \N__52334\ : std_logic;
signal \N__52331\ : std_logic;
signal \N__52328\ : std_logic;
signal \N__52323\ : std_logic;
signal \N__52320\ : std_logic;
signal \N__52319\ : std_logic;
signal \N__52316\ : std_logic;
signal \N__52313\ : std_logic;
signal \N__52310\ : std_logic;
signal \N__52307\ : std_logic;
signal \N__52304\ : std_logic;
signal \N__52293\ : std_logic;
signal \N__52288\ : std_logic;
signal \N__52283\ : std_logic;
signal \N__52280\ : std_logic;
signal \N__52277\ : std_logic;
signal \N__52274\ : std_logic;
signal \N__52267\ : std_logic;
signal \N__52264\ : std_logic;
signal \N__52257\ : std_logic;
signal \N__52246\ : std_logic;
signal \N__52243\ : std_logic;
signal \N__52240\ : std_logic;
signal \N__52237\ : std_logic;
signal \N__52234\ : std_logic;
signal \N__52233\ : std_logic;
signal \N__52232\ : std_logic;
signal \N__52229\ : std_logic;
signal \N__52226\ : std_logic;
signal \N__52223\ : std_logic;
signal \N__52220\ : std_logic;
signal \N__52217\ : std_logic;
signal \N__52214\ : std_logic;
signal \N__52211\ : std_logic;
signal \N__52208\ : std_logic;
signal \N__52205\ : std_logic;
signal \N__52198\ : std_logic;
signal \N__52195\ : std_logic;
signal \N__52194\ : std_logic;
signal \N__52193\ : std_logic;
signal \N__52192\ : std_logic;
signal \N__52191\ : std_logic;
signal \N__52190\ : std_logic;
signal \N__52189\ : std_logic;
signal \N__52186\ : std_logic;
signal \N__52185\ : std_logic;
signal \N__52182\ : std_logic;
signal \N__52181\ : std_logic;
signal \N__52178\ : std_logic;
signal \N__52177\ : std_logic;
signal \N__52176\ : std_logic;
signal \N__52175\ : std_logic;
signal \N__52174\ : std_logic;
signal \N__52173\ : std_logic;
signal \N__52172\ : std_logic;
signal \N__52171\ : std_logic;
signal \N__52170\ : std_logic;
signal \N__52169\ : std_logic;
signal \N__52168\ : std_logic;
signal \N__52167\ : std_logic;
signal \N__52166\ : std_logic;
signal \N__52163\ : std_logic;
signal \N__52162\ : std_logic;
signal \N__52161\ : std_logic;
signal \N__52160\ : std_logic;
signal \N__52159\ : std_logic;
signal \N__52158\ : std_logic;
signal \N__52151\ : std_logic;
signal \N__52148\ : std_logic;
signal \N__52147\ : std_logic;
signal \N__52140\ : std_logic;
signal \N__52135\ : std_logic;
signal \N__52132\ : std_logic;
signal \N__52125\ : std_logic;
signal \N__52124\ : std_logic;
signal \N__52123\ : std_logic;
signal \N__52120\ : std_logic;
signal \N__52117\ : std_logic;
signal \N__52114\ : std_logic;
signal \N__52113\ : std_logic;
signal \N__52112\ : std_logic;
signal \N__52111\ : std_logic;
signal \N__52110\ : std_logic;
signal \N__52109\ : std_logic;
signal \N__52108\ : std_logic;
signal \N__52105\ : std_logic;
signal \N__52102\ : std_logic;
signal \N__52099\ : std_logic;
signal \N__52096\ : std_logic;
signal \N__52093\ : std_logic;
signal \N__52092\ : std_logic;
signal \N__52091\ : std_logic;
signal \N__52088\ : std_logic;
signal \N__52087\ : std_logic;
signal \N__52084\ : std_logic;
signal \N__52081\ : std_logic;
signal \N__52078\ : std_logic;
signal \N__52077\ : std_logic;
signal \N__52074\ : std_logic;
signal \N__52069\ : std_logic;
signal \N__52066\ : std_logic;
signal \N__52065\ : std_logic;
signal \N__52064\ : std_logic;
signal \N__52063\ : std_logic;
signal \N__52062\ : std_logic;
signal \N__52061\ : std_logic;
signal \N__52060\ : std_logic;
signal \N__52059\ : std_logic;
signal \N__52050\ : std_logic;
signal \N__52047\ : std_logic;
signal \N__52044\ : std_logic;
signal \N__52043\ : std_logic;
signal \N__52042\ : std_logic;
signal \N__52037\ : std_logic;
signal \N__52034\ : std_logic;
signal \N__52033\ : std_logic;
signal \N__52030\ : std_logic;
signal \N__52027\ : std_logic;
signal \N__52024\ : std_logic;
signal \N__52017\ : std_logic;
signal \N__52012\ : std_logic;
signal \N__52007\ : std_logic;
signal \N__52004\ : std_logic;
signal \N__52001\ : std_logic;
signal \N__51998\ : std_logic;
signal \N__51995\ : std_logic;
signal \N__51986\ : std_logic;
signal \N__51985\ : std_logic;
signal \N__51984\ : std_logic;
signal \N__51983\ : std_logic;
signal \N__51980\ : std_logic;
signal \N__51979\ : std_logic;
signal \N__51978\ : std_logic;
signal \N__51977\ : std_logic;
signal \N__51976\ : std_logic;
signal \N__51975\ : std_logic;
signal \N__51974\ : std_logic;
signal \N__51971\ : std_logic;
signal \N__51968\ : std_logic;
signal \N__51963\ : std_logic;
signal \N__51958\ : std_logic;
signal \N__51955\ : std_logic;
signal \N__51952\ : std_logic;
signal \N__51951\ : std_logic;
signal \N__51950\ : std_logic;
signal \N__51945\ : std_logic;
signal \N__51942\ : std_logic;
signal \N__51937\ : std_logic;
signal \N__51934\ : std_logic;
signal \N__51931\ : std_logic;
signal \N__51930\ : std_logic;
signal \N__51929\ : std_logic;
signal \N__51924\ : std_logic;
signal \N__51921\ : std_logic;
signal \N__51920\ : std_logic;
signal \N__51919\ : std_logic;
signal \N__51916\ : std_logic;
signal \N__51915\ : std_logic;
signal \N__51914\ : std_logic;
signal \N__51907\ : std_logic;
signal \N__51900\ : std_logic;
signal \N__51895\ : std_logic;
signal \N__51894\ : std_logic;
signal \N__51893\ : std_logic;
signal \N__51888\ : std_logic;
signal \N__51885\ : std_logic;
signal \N__51882\ : std_logic;
signal \N__51881\ : std_logic;
signal \N__51878\ : std_logic;
signal \N__51873\ : std_logic;
signal \N__51870\ : std_logic;
signal \N__51861\ : std_logic;
signal \N__51852\ : std_logic;
signal \N__51849\ : std_logic;
signal \N__51842\ : std_logic;
signal \N__51835\ : std_logic;
signal \N__51826\ : std_logic;
signal \N__51823\ : std_logic;
signal \N__51818\ : std_logic;
signal \N__51815\ : std_logic;
signal \N__51812\ : std_logic;
signal \N__51807\ : std_logic;
signal \N__51800\ : std_logic;
signal \N__51795\ : std_logic;
signal \N__51792\ : std_logic;
signal \N__51787\ : std_logic;
signal \N__51786\ : std_logic;
signal \N__51783\ : std_logic;
signal \N__51782\ : std_logic;
signal \N__51763\ : std_logic;
signal \N__51758\ : std_logic;
signal \N__51755\ : std_logic;
signal \N__51752\ : std_logic;
signal \N__51747\ : std_logic;
signal \N__51740\ : std_logic;
signal \N__51737\ : std_logic;
signal \N__51734\ : std_logic;
signal \N__51731\ : std_logic;
signal \N__51728\ : std_logic;
signal \N__51725\ : std_logic;
signal \N__51716\ : std_logic;
signal \N__51703\ : std_logic;
signal \N__51700\ : std_logic;
signal \N__51697\ : std_logic;
signal \N__51694\ : std_logic;
signal \N__51691\ : std_logic;
signal \N__51688\ : std_logic;
signal \N__51685\ : std_logic;
signal \N__51684\ : std_logic;
signal \N__51681\ : std_logic;
signal \N__51678\ : std_logic;
signal \N__51677\ : std_logic;
signal \N__51674\ : std_logic;
signal \N__51671\ : std_logic;
signal \N__51668\ : std_logic;
signal \N__51665\ : std_logic;
signal \N__51660\ : std_logic;
signal \N__51659\ : std_logic;
signal \N__51656\ : std_logic;
signal \N__51653\ : std_logic;
signal \N__51650\ : std_logic;
signal \N__51643\ : std_logic;
signal \N__51642\ : std_logic;
signal \N__51641\ : std_logic;
signal \N__51640\ : std_logic;
signal \N__51639\ : std_logic;
signal \N__51638\ : std_logic;
signal \N__51633\ : std_logic;
signal \N__51632\ : std_logic;
signal \N__51631\ : std_logic;
signal \N__51630\ : std_logic;
signal \N__51629\ : std_logic;
signal \N__51628\ : std_logic;
signal \N__51627\ : std_logic;
signal \N__51626\ : std_logic;
signal \N__51625\ : std_logic;
signal \N__51624\ : std_logic;
signal \N__51623\ : std_logic;
signal \N__51622\ : std_logic;
signal \N__51621\ : std_logic;
signal \N__51620\ : std_logic;
signal \N__51619\ : std_logic;
signal \N__51610\ : std_logic;
signal \N__51607\ : std_logic;
signal \N__51606\ : std_logic;
signal \N__51605\ : std_logic;
signal \N__51604\ : std_logic;
signal \N__51601\ : std_logic;
signal \N__51592\ : std_logic;
signal \N__51583\ : std_logic;
signal \N__51580\ : std_logic;
signal \N__51579\ : std_logic;
signal \N__51578\ : std_logic;
signal \N__51577\ : std_logic;
signal \N__51570\ : std_logic;
signal \N__51567\ : std_logic;
signal \N__51564\ : std_logic;
signal \N__51561\ : std_logic;
signal \N__51554\ : std_logic;
signal \N__51551\ : std_logic;
signal \N__51544\ : std_logic;
signal \N__51541\ : std_logic;
signal \N__51538\ : std_logic;
signal \N__51537\ : std_logic;
signal \N__51534\ : std_logic;
signal \N__51533\ : std_logic;
signal \N__51530\ : std_logic;
signal \N__51529\ : std_logic;
signal \N__51526\ : std_logic;
signal \N__51519\ : std_logic;
signal \N__51518\ : std_logic;
signal \N__51517\ : std_logic;
signal \N__51516\ : std_logic;
signal \N__51515\ : std_logic;
signal \N__51510\ : std_logic;
signal \N__51505\ : std_logic;
signal \N__51498\ : std_logic;
signal \N__51495\ : std_logic;
signal \N__51492\ : std_logic;
signal \N__51487\ : std_logic;
signal \N__51478\ : std_logic;
signal \N__51473\ : std_logic;
signal \N__51460\ : std_logic;
signal \N__51457\ : std_logic;
signal \N__51454\ : std_logic;
signal \N__51451\ : std_logic;
signal \N__51448\ : std_logic;
signal \N__51445\ : std_logic;
signal \N__51442\ : std_logic;
signal \N__51439\ : std_logic;
signal \N__51438\ : std_logic;
signal \N__51435\ : std_logic;
signal \N__51432\ : std_logic;
signal \N__51431\ : std_logic;
signal \N__51430\ : std_logic;
signal \N__51429\ : std_logic;
signal \N__51428\ : std_logic;
signal \N__51425\ : std_logic;
signal \N__51420\ : std_logic;
signal \N__51417\ : std_logic;
signal \N__51414\ : std_logic;
signal \N__51411\ : std_logic;
signal \N__51406\ : std_logic;
signal \N__51403\ : std_logic;
signal \N__51400\ : std_logic;
signal \N__51397\ : std_logic;
signal \N__51394\ : std_logic;
signal \N__51391\ : std_logic;
signal \N__51386\ : std_logic;
signal \N__51383\ : std_logic;
signal \N__51376\ : std_logic;
signal \N__51375\ : std_logic;
signal \N__51372\ : std_logic;
signal \N__51369\ : std_logic;
signal \N__51364\ : std_logic;
signal \N__51361\ : std_logic;
signal \N__51358\ : std_logic;
signal \N__51355\ : std_logic;
signal \N__51352\ : std_logic;
signal \N__51349\ : std_logic;
signal \N__51346\ : std_logic;
signal \N__51343\ : std_logic;
signal \N__51342\ : std_logic;
signal \N__51339\ : std_logic;
signal \N__51336\ : std_logic;
signal \N__51331\ : std_logic;
signal \N__51330\ : std_logic;
signal \N__51327\ : std_logic;
signal \N__51326\ : std_logic;
signal \N__51323\ : std_logic;
signal \N__51320\ : std_logic;
signal \N__51317\ : std_logic;
signal \N__51310\ : std_logic;
signal \N__51307\ : std_logic;
signal \N__51304\ : std_logic;
signal \N__51301\ : std_logic;
signal \N__51298\ : std_logic;
signal \N__51297\ : std_logic;
signal \N__51294\ : std_logic;
signal \N__51293\ : std_logic;
signal \N__51290\ : std_logic;
signal \N__51287\ : std_logic;
signal \N__51286\ : std_logic;
signal \N__51285\ : std_logic;
signal \N__51284\ : std_logic;
signal \N__51283\ : std_logic;
signal \N__51282\ : std_logic;
signal \N__51279\ : std_logic;
signal \N__51276\ : std_logic;
signal \N__51273\ : std_logic;
signal \N__51268\ : std_logic;
signal \N__51265\ : std_logic;
signal \N__51264\ : std_logic;
signal \N__51263\ : std_logic;
signal \N__51262\ : std_logic;
signal \N__51261\ : std_logic;
signal \N__51260\ : std_logic;
signal \N__51259\ : std_logic;
signal \N__51254\ : std_logic;
signal \N__51251\ : std_logic;
signal \N__51244\ : std_logic;
signal \N__51241\ : std_logic;
signal \N__51240\ : std_logic;
signal \N__51239\ : std_logic;
signal \N__51238\ : std_logic;
signal \N__51235\ : std_logic;
signal \N__51234\ : std_logic;
signal \N__51231\ : std_logic;
signal \N__51230\ : std_logic;
signal \N__51229\ : std_logic;
signal \N__51228\ : std_logic;
signal \N__51227\ : std_logic;
signal \N__51226\ : std_logic;
signal \N__51225\ : std_logic;
signal \N__51222\ : std_logic;
signal \N__51221\ : std_logic;
signal \N__51220\ : std_logic;
signal \N__51219\ : std_logic;
signal \N__51218\ : std_logic;
signal \N__51217\ : std_logic;
signal \N__51214\ : std_logic;
signal \N__51211\ : std_logic;
signal \N__51210\ : std_logic;
signal \N__51209\ : std_logic;
signal \N__51208\ : std_logic;
signal \N__51207\ : std_logic;
signal \N__51206\ : std_logic;
signal \N__51205\ : std_logic;
signal \N__51204\ : std_logic;
signal \N__51201\ : std_logic;
signal \N__51200\ : std_logic;
signal \N__51199\ : std_logic;
signal \N__51198\ : std_logic;
signal \N__51197\ : std_logic;
signal \N__51196\ : std_logic;
signal \N__51193\ : std_logic;
signal \N__51186\ : std_logic;
signal \N__51181\ : std_logic;
signal \N__51178\ : std_logic;
signal \N__51169\ : std_logic;
signal \N__51166\ : std_logic;
signal \N__51163\ : std_logic;
signal \N__51156\ : std_logic;
signal \N__51153\ : std_logic;
signal \N__51150\ : std_logic;
signal \N__51143\ : std_logic;
signal \N__51134\ : std_logic;
signal \N__51129\ : std_logic;
signal \N__51126\ : std_logic;
signal \N__51123\ : std_logic;
signal \N__51118\ : std_logic;
signal \N__51115\ : std_logic;
signal \N__51112\ : std_logic;
signal \N__51111\ : std_logic;
signal \N__51110\ : std_logic;
signal \N__51107\ : std_logic;
signal \N__51106\ : std_logic;
signal \N__51105\ : std_logic;
signal \N__51104\ : std_logic;
signal \N__51101\ : std_logic;
signal \N__51096\ : std_logic;
signal \N__51087\ : std_logic;
signal \N__51084\ : std_logic;
signal \N__51075\ : std_logic;
signal \N__51074\ : std_logic;
signal \N__51073\ : std_logic;
signal \N__51070\ : std_logic;
signal \N__51063\ : std_logic;
signal \N__51062\ : std_logic;
signal \N__51061\ : std_logic;
signal \N__51058\ : std_logic;
signal \N__51049\ : std_logic;
signal \N__51044\ : std_logic;
signal \N__51041\ : std_logic;
signal \N__51038\ : std_logic;
signal \N__51033\ : std_logic;
signal \N__51022\ : std_logic;
signal \N__51017\ : std_logic;
signal \N__51014\ : std_logic;
signal \N__51011\ : std_logic;
signal \N__51006\ : std_logic;
signal \N__51001\ : std_logic;
signal \N__50980\ : std_logic;
signal \N__50977\ : std_logic;
signal \N__50974\ : std_logic;
signal \N__50971\ : std_logic;
signal \N__50968\ : std_logic;
signal \N__50965\ : std_logic;
signal \N__50964\ : std_logic;
signal \N__50963\ : std_logic;
signal \N__50962\ : std_logic;
signal \N__50961\ : std_logic;
signal \N__50960\ : std_logic;
signal \N__50957\ : std_logic;
signal \N__50956\ : std_logic;
signal \N__50955\ : std_logic;
signal \N__50954\ : std_logic;
signal \N__50953\ : std_logic;
signal \N__50952\ : std_logic;
signal \N__50951\ : std_logic;
signal \N__50950\ : std_logic;
signal \N__50949\ : std_logic;
signal \N__50948\ : std_logic;
signal \N__50945\ : std_logic;
signal \N__50938\ : std_logic;
signal \N__50937\ : std_logic;
signal \N__50936\ : std_logic;
signal \N__50935\ : std_logic;
signal \N__50934\ : std_logic;
signal \N__50931\ : std_logic;
signal \N__50922\ : std_logic;
signal \N__50921\ : std_logic;
signal \N__50920\ : std_logic;
signal \N__50919\ : std_logic;
signal \N__50916\ : std_logic;
signal \N__50915\ : std_logic;
signal \N__50914\ : std_logic;
signal \N__50913\ : std_logic;
signal \N__50912\ : std_logic;
signal \N__50911\ : std_logic;
signal \N__50910\ : std_logic;
signal \N__50909\ : std_logic;
signal \N__50908\ : std_logic;
signal \N__50907\ : std_logic;
signal \N__50906\ : std_logic;
signal \N__50903\ : std_logic;
signal \N__50896\ : std_logic;
signal \N__50893\ : std_logic;
signal \N__50888\ : std_logic;
signal \N__50885\ : std_logic;
signal \N__50884\ : std_logic;
signal \N__50883\ : std_logic;
signal \N__50882\ : std_logic;
signal \N__50881\ : std_logic;
signal \N__50880\ : std_logic;
signal \N__50877\ : std_logic;
signal \N__50872\ : std_logic;
signal \N__50867\ : std_logic;
signal \N__50860\ : std_logic;
signal \N__50857\ : std_logic;
signal \N__50856\ : std_logic;
signal \N__50855\ : std_logic;
signal \N__50852\ : std_logic;
signal \N__50849\ : std_logic;
signal \N__50844\ : std_logic;
signal \N__50841\ : std_logic;
signal \N__50838\ : std_logic;
signal \N__50837\ : std_logic;
signal \N__50836\ : std_logic;
signal \N__50835\ : std_logic;
signal \N__50834\ : std_logic;
signal \N__50831\ : std_logic;
signal \N__50830\ : std_logic;
signal \N__50825\ : std_logic;
signal \N__50822\ : std_logic;
signal \N__50821\ : std_logic;
signal \N__50818\ : std_logic;
signal \N__50813\ : std_logic;
signal \N__50810\ : std_logic;
signal \N__50805\ : std_logic;
signal \N__50802\ : std_logic;
signal \N__50801\ : std_logic;
signal \N__50798\ : std_logic;
signal \N__50793\ : std_logic;
signal \N__50788\ : std_logic;
signal \N__50781\ : std_logic;
signal \N__50776\ : std_logic;
signal \N__50771\ : std_logic;
signal \N__50766\ : std_logic;
signal \N__50763\ : std_logic;
signal \N__50760\ : std_logic;
signal \N__50759\ : std_logic;
signal \N__50756\ : std_logic;
signal \N__50753\ : std_logic;
signal \N__50750\ : std_logic;
signal \N__50749\ : std_logic;
signal \N__50748\ : std_logic;
signal \N__50747\ : std_logic;
signal \N__50746\ : std_logic;
signal \N__50741\ : std_logic;
signal \N__50736\ : std_logic;
signal \N__50733\ : std_logic;
signal \N__50730\ : std_logic;
signal \N__50725\ : std_logic;
signal \N__50724\ : std_logic;
signal \N__50723\ : std_logic;
signal \N__50718\ : std_logic;
signal \N__50717\ : std_logic;
signal \N__50716\ : std_logic;
signal \N__50715\ : std_logic;
signal \N__50714\ : std_logic;
signal \N__50713\ : std_logic;
signal \N__50712\ : std_logic;
signal \N__50711\ : std_logic;
signal \N__50710\ : std_logic;
signal \N__50707\ : std_logic;
signal \N__50704\ : std_logic;
signal \N__50695\ : std_logic;
signal \N__50692\ : std_logic;
signal \N__50689\ : std_logic;
signal \N__50686\ : std_logic;
signal \N__50681\ : std_logic;
signal \N__50666\ : std_logic;
signal \N__50663\ : std_logic;
signal \N__50660\ : std_logic;
signal \N__50657\ : std_logic;
signal \N__50652\ : std_logic;
signal \N__50651\ : std_logic;
signal \N__50650\ : std_logic;
signal \N__50649\ : std_logic;
signal \N__50648\ : std_logic;
signal \N__50647\ : std_logic;
signal \N__50646\ : std_logic;
signal \N__50645\ : std_logic;
signal \N__50642\ : std_logic;
signal \N__50639\ : std_logic;
signal \N__50636\ : std_logic;
signal \N__50619\ : std_logic;
signal \N__50614\ : std_logic;
signal \N__50611\ : std_logic;
signal \N__50606\ : std_logic;
signal \N__50603\ : std_logic;
signal \N__50594\ : std_logic;
signal \N__50589\ : std_logic;
signal \N__50582\ : std_logic;
signal \N__50573\ : std_logic;
signal \N__50548\ : std_logic;
signal \N__50547\ : std_logic;
signal \N__50544\ : std_logic;
signal \N__50541\ : std_logic;
signal \N__50540\ : std_logic;
signal \N__50537\ : std_logic;
signal \N__50532\ : std_logic;
signal \N__50527\ : std_logic;
signal \N__50526\ : std_logic;
signal \N__50523\ : std_logic;
signal \N__50520\ : std_logic;
signal \N__50519\ : std_logic;
signal \N__50518\ : std_logic;
signal \N__50517\ : std_logic;
signal \N__50516\ : std_logic;
signal \N__50515\ : std_logic;
signal \N__50514\ : std_logic;
signal \N__50513\ : std_logic;
signal \N__50512\ : std_logic;
signal \N__50507\ : std_logic;
signal \N__50502\ : std_logic;
signal \N__50501\ : std_logic;
signal \N__50500\ : std_logic;
signal \N__50497\ : std_logic;
signal \N__50496\ : std_logic;
signal \N__50495\ : std_logic;
signal \N__50494\ : std_logic;
signal \N__50493\ : std_logic;
signal \N__50492\ : std_logic;
signal \N__50491\ : std_logic;
signal \N__50486\ : std_logic;
signal \N__50483\ : std_logic;
signal \N__50480\ : std_logic;
signal \N__50479\ : std_logic;
signal \N__50476\ : std_logic;
signal \N__50471\ : std_logic;
signal \N__50470\ : std_logic;
signal \N__50469\ : std_logic;
signal \N__50466\ : std_logic;
signal \N__50463\ : std_logic;
signal \N__50460\ : std_logic;
signal \N__50459\ : std_logic;
signal \N__50458\ : std_logic;
signal \N__50457\ : std_logic;
signal \N__50456\ : std_logic;
signal \N__50455\ : std_logic;
signal \N__50454\ : std_logic;
signal \N__50453\ : std_logic;
signal \N__50448\ : std_logic;
signal \N__50443\ : std_logic;
signal \N__50438\ : std_logic;
signal \N__50431\ : std_logic;
signal \N__50428\ : std_logic;
signal \N__50425\ : std_logic;
signal \N__50422\ : std_logic;
signal \N__50419\ : std_logic;
signal \N__50418\ : std_logic;
signal \N__50417\ : std_logic;
signal \N__50416\ : std_logic;
signal \N__50415\ : std_logic;
signal \N__50412\ : std_logic;
signal \N__50409\ : std_logic;
signal \N__50406\ : std_logic;
signal \N__50403\ : std_logic;
signal \N__50390\ : std_logic;
signal \N__50387\ : std_logic;
signal \N__50378\ : std_logic;
signal \N__50373\ : std_logic;
signal \N__50370\ : std_logic;
signal \N__50367\ : std_logic;
signal \N__50358\ : std_logic;
signal \N__50353\ : std_logic;
signal \N__50350\ : std_logic;
signal \N__50347\ : std_logic;
signal \N__50336\ : std_logic;
signal \N__50323\ : std_logic;
signal \N__50322\ : std_logic;
signal \N__50319\ : std_logic;
signal \N__50316\ : std_logic;
signal \N__50315\ : std_logic;
signal \N__50312\ : std_logic;
signal \N__50309\ : std_logic;
signal \N__50306\ : std_logic;
signal \N__50299\ : std_logic;
signal \N__50296\ : std_logic;
signal \N__50293\ : std_logic;
signal \N__50292\ : std_logic;
signal \N__50289\ : std_logic;
signal \N__50286\ : std_logic;
signal \N__50285\ : std_logic;
signal \N__50282\ : std_logic;
signal \N__50279\ : std_logic;
signal \N__50276\ : std_logic;
signal \N__50273\ : std_logic;
signal \N__50266\ : std_logic;
signal \N__50263\ : std_logic;
signal \N__50260\ : std_logic;
signal \N__50257\ : std_logic;
signal \N__50256\ : std_logic;
signal \N__50255\ : std_logic;
signal \N__50252\ : std_logic;
signal \N__50249\ : std_logic;
signal \N__50246\ : std_logic;
signal \N__50239\ : std_logic;
signal \N__50236\ : std_logic;
signal \N__50233\ : std_logic;
signal \N__50230\ : std_logic;
signal \N__50227\ : std_logic;
signal \N__50224\ : std_logic;
signal \N__50221\ : std_logic;
signal \N__50220\ : std_logic;
signal \N__50217\ : std_logic;
signal \N__50214\ : std_logic;
signal \N__50211\ : std_logic;
signal \N__50206\ : std_logic;
signal \N__50205\ : std_logic;
signal \N__50202\ : std_logic;
signal \N__50199\ : std_logic;
signal \N__50194\ : std_logic;
signal \N__50191\ : std_logic;
signal \N__50190\ : std_logic;
signal \N__50187\ : std_logic;
signal \N__50184\ : std_logic;
signal \N__50183\ : std_logic;
signal \N__50182\ : std_logic;
signal \N__50181\ : std_logic;
signal \N__50178\ : std_logic;
signal \N__50175\ : std_logic;
signal \N__50172\ : std_logic;
signal \N__50169\ : std_logic;
signal \N__50166\ : std_logic;
signal \N__50163\ : std_logic;
signal \N__50158\ : std_logic;
signal \N__50155\ : std_logic;
signal \N__50148\ : std_logic;
signal \N__50145\ : std_logic;
signal \N__50142\ : std_logic;
signal \N__50137\ : std_logic;
signal \N__50136\ : std_logic;
signal \N__50133\ : std_logic;
signal \N__50132\ : std_logic;
signal \N__50129\ : std_logic;
signal \N__50126\ : std_logic;
signal \N__50123\ : std_logic;
signal \N__50120\ : std_logic;
signal \N__50115\ : std_logic;
signal \N__50110\ : std_logic;
signal \N__50107\ : std_logic;
signal \N__50104\ : std_logic;
signal \N__50101\ : std_logic;
signal \N__50100\ : std_logic;
signal \N__50099\ : std_logic;
signal \N__50098\ : std_logic;
signal \N__50097\ : std_logic;
signal \N__50096\ : std_logic;
signal \N__50095\ : std_logic;
signal \N__50094\ : std_logic;
signal \N__50089\ : std_logic;
signal \N__50088\ : std_logic;
signal \N__50087\ : std_logic;
signal \N__50082\ : std_logic;
signal \N__50079\ : std_logic;
signal \N__50078\ : std_logic;
signal \N__50077\ : std_logic;
signal \N__50076\ : std_logic;
signal \N__50075\ : std_logic;
signal \N__50070\ : std_logic;
signal \N__50069\ : std_logic;
signal \N__50068\ : std_logic;
signal \N__50067\ : std_logic;
signal \N__50064\ : std_logic;
signal \N__50061\ : std_logic;
signal \N__50058\ : std_logic;
signal \N__50055\ : std_logic;
signal \N__50050\ : std_logic;
signal \N__50047\ : std_logic;
signal \N__50040\ : std_logic;
signal \N__50037\ : std_logic;
signal \N__50030\ : std_logic;
signal \N__50027\ : std_logic;
signal \N__50016\ : std_logic;
signal \N__50011\ : std_logic;
signal \N__50010\ : std_logic;
signal \N__50009\ : std_logic;
signal \N__50008\ : std_logic;
signal \N__50007\ : std_logic;
signal \N__50006\ : std_logic;
signal \N__50003\ : std_logic;
signal \N__50002\ : std_logic;
signal \N__49999\ : std_logic;
signal \N__49994\ : std_logic;
signal \N__49989\ : std_logic;
signal \N__49986\ : std_logic;
signal \N__49981\ : std_logic;
signal \N__49978\ : std_logic;
signal \N__49975\ : std_logic;
signal \N__49968\ : std_logic;
signal \N__49957\ : std_logic;
signal \N__49954\ : std_logic;
signal \N__49951\ : std_logic;
signal \N__49948\ : std_logic;
signal \N__49947\ : std_logic;
signal \N__49944\ : std_logic;
signal \N__49941\ : std_logic;
signal \N__49940\ : std_logic;
signal \N__49939\ : std_logic;
signal \N__49936\ : std_logic;
signal \N__49933\ : std_logic;
signal \N__49930\ : std_logic;
signal \N__49927\ : std_logic;
signal \N__49918\ : std_logic;
signal \N__49915\ : std_logic;
signal \N__49914\ : std_logic;
signal \N__49911\ : std_logic;
signal \N__49910\ : std_logic;
signal \N__49909\ : std_logic;
signal \N__49908\ : std_logic;
signal \N__49905\ : std_logic;
signal \N__49902\ : std_logic;
signal \N__49897\ : std_logic;
signal \N__49894\ : std_logic;
signal \N__49891\ : std_logic;
signal \N__49888\ : std_logic;
signal \N__49883\ : std_logic;
signal \N__49876\ : std_logic;
signal \N__49873\ : std_logic;
signal \N__49870\ : std_logic;
signal \N__49869\ : std_logic;
signal \N__49864\ : std_logic;
signal \N__49861\ : std_logic;
signal \N__49860\ : std_logic;
signal \N__49859\ : std_logic;
signal \N__49858\ : std_logic;
signal \N__49855\ : std_logic;
signal \N__49850\ : std_logic;
signal \N__49847\ : std_logic;
signal \N__49846\ : std_logic;
signal \N__49839\ : std_logic;
signal \N__49836\ : std_logic;
signal \N__49831\ : std_logic;
signal \N__49828\ : std_logic;
signal \N__49825\ : std_logic;
signal \N__49822\ : std_logic;
signal \N__49821\ : std_logic;
signal \N__49818\ : std_logic;
signal \N__49815\ : std_logic;
signal \N__49812\ : std_logic;
signal \N__49809\ : std_logic;
signal \N__49804\ : std_logic;
signal \N__49801\ : std_logic;
signal \N__49800\ : std_logic;
signal \N__49799\ : std_logic;
signal \N__49798\ : std_logic;
signal \N__49797\ : std_logic;
signal \N__49796\ : std_logic;
signal \N__49795\ : std_logic;
signal \N__49792\ : std_logic;
signal \N__49791\ : std_logic;
signal \N__49790\ : std_logic;
signal \N__49783\ : std_logic;
signal \N__49782\ : std_logic;
signal \N__49781\ : std_logic;
signal \N__49778\ : std_logic;
signal \N__49775\ : std_logic;
signal \N__49774\ : std_logic;
signal \N__49771\ : std_logic;
signal \N__49770\ : std_logic;
signal \N__49769\ : std_logic;
signal \N__49768\ : std_logic;
signal \N__49767\ : std_logic;
signal \N__49764\ : std_logic;
signal \N__49759\ : std_logic;
signal \N__49756\ : std_logic;
signal \N__49755\ : std_logic;
signal \N__49752\ : std_logic;
signal \N__49751\ : std_logic;
signal \N__49750\ : std_logic;
signal \N__49747\ : std_logic;
signal \N__49744\ : std_logic;
signal \N__49735\ : std_logic;
signal \N__49730\ : std_logic;
signal \N__49727\ : std_logic;
signal \N__49722\ : std_logic;
signal \N__49719\ : std_logic;
signal \N__49712\ : std_logic;
signal \N__49709\ : std_logic;
signal \N__49700\ : std_logic;
signal \N__49699\ : std_logic;
signal \N__49696\ : std_logic;
signal \N__49693\ : std_logic;
signal \N__49690\ : std_logic;
signal \N__49683\ : std_logic;
signal \N__49680\ : std_logic;
signal \N__49677\ : std_logic;
signal \N__49674\ : std_logic;
signal \N__49671\ : std_logic;
signal \N__49666\ : std_logic;
signal \N__49661\ : std_logic;
signal \N__49656\ : std_logic;
signal \N__49653\ : std_logic;
signal \N__49650\ : std_logic;
signal \N__49645\ : std_logic;
signal \N__49642\ : std_logic;
signal \N__49641\ : std_logic;
signal \N__49640\ : std_logic;
signal \N__49639\ : std_logic;
signal \N__49636\ : std_logic;
signal \N__49635\ : std_logic;
signal \N__49634\ : std_logic;
signal \N__49633\ : std_logic;
signal \N__49632\ : std_logic;
signal \N__49629\ : std_logic;
signal \N__49628\ : std_logic;
signal \N__49627\ : std_logic;
signal \N__49626\ : std_logic;
signal \N__49625\ : std_logic;
signal \N__49624\ : std_logic;
signal \N__49619\ : std_logic;
signal \N__49616\ : std_logic;
signal \N__49613\ : std_logic;
signal \N__49610\ : std_logic;
signal \N__49605\ : std_logic;
signal \N__49602\ : std_logic;
signal \N__49593\ : std_logic;
signal \N__49590\ : std_logic;
signal \N__49573\ : std_logic;
signal \N__49570\ : std_logic;
signal \N__49567\ : std_logic;
signal \N__49564\ : std_logic;
signal \N__49561\ : std_logic;
signal \N__49558\ : std_logic;
signal \N__49555\ : std_logic;
signal \N__49552\ : std_logic;
signal \N__49549\ : std_logic;
signal \N__49546\ : std_logic;
signal \N__49543\ : std_logic;
signal \N__49540\ : std_logic;
signal \N__49539\ : std_logic;
signal \N__49538\ : std_logic;
signal \N__49537\ : std_logic;
signal \N__49536\ : std_logic;
signal \N__49535\ : std_logic;
signal \N__49534\ : std_logic;
signal \N__49533\ : std_logic;
signal \N__49532\ : std_logic;
signal \N__49531\ : std_logic;
signal \N__49530\ : std_logic;
signal \N__49529\ : std_logic;
signal \N__49526\ : std_logic;
signal \N__49525\ : std_logic;
signal \N__49524\ : std_logic;
signal \N__49523\ : std_logic;
signal \N__49522\ : std_logic;
signal \N__49521\ : std_logic;
signal \N__49520\ : std_logic;
signal \N__49515\ : std_logic;
signal \N__49514\ : std_logic;
signal \N__49513\ : std_logic;
signal \N__49506\ : std_logic;
signal \N__49503\ : std_logic;
signal \N__49500\ : std_logic;
signal \N__49493\ : std_logic;
signal \N__49492\ : std_logic;
signal \N__49489\ : std_logic;
signal \N__49486\ : std_logic;
signal \N__49481\ : std_logic;
signal \N__49476\ : std_logic;
signal \N__49471\ : std_logic;
signal \N__49468\ : std_logic;
signal \N__49467\ : std_logic;
signal \N__49464\ : std_logic;
signal \N__49463\ : std_logic;
signal \N__49462\ : std_logic;
signal \N__49459\ : std_logic;
signal \N__49456\ : std_logic;
signal \N__49451\ : std_logic;
signal \N__49448\ : std_logic;
signal \N__49445\ : std_logic;
signal \N__49442\ : std_logic;
signal \N__49435\ : std_logic;
signal \N__49430\ : std_logic;
signal \N__49429\ : std_logic;
signal \N__49426\ : std_logic;
signal \N__49423\ : std_logic;
signal \N__49420\ : std_logic;
signal \N__49417\ : std_logic;
signal \N__49414\ : std_logic;
signal \N__49407\ : std_logic;
signal \N__49404\ : std_logic;
signal \N__49397\ : std_logic;
signal \N__49396\ : std_logic;
signal \N__49395\ : std_logic;
signal \N__49392\ : std_logic;
signal \N__49387\ : std_logic;
signal \N__49384\ : std_logic;
signal \N__49375\ : std_logic;
signal \N__49372\ : std_logic;
signal \N__49367\ : std_logic;
signal \N__49364\ : std_logic;
signal \N__49361\ : std_logic;
signal \N__49348\ : std_logic;
signal \N__49345\ : std_logic;
signal \N__49344\ : std_logic;
signal \N__49341\ : std_logic;
signal \N__49338\ : std_logic;
signal \N__49335\ : std_logic;
signal \N__49332\ : std_logic;
signal \N__49327\ : std_logic;
signal \N__49324\ : std_logic;
signal \N__49323\ : std_logic;
signal \N__49320\ : std_logic;
signal \N__49317\ : std_logic;
signal \N__49314\ : std_logic;
signal \N__49311\ : std_logic;
signal \N__49306\ : std_logic;
signal \N__49303\ : std_logic;
signal \N__49302\ : std_logic;
signal \N__49299\ : std_logic;
signal \N__49298\ : std_logic;
signal \N__49295\ : std_logic;
signal \N__49292\ : std_logic;
signal \N__49289\ : std_logic;
signal \N__49288\ : std_logic;
signal \N__49281\ : std_logic;
signal \N__49278\ : std_logic;
signal \N__49275\ : std_logic;
signal \N__49270\ : std_logic;
signal \N__49267\ : std_logic;
signal \N__49264\ : std_logic;
signal \N__49261\ : std_logic;
signal \N__49258\ : std_logic;
signal \N__49255\ : std_logic;
signal \N__49252\ : std_logic;
signal \N__49249\ : std_logic;
signal \N__49246\ : std_logic;
signal \N__49243\ : std_logic;
signal \N__49240\ : std_logic;
signal \N__49239\ : std_logic;
signal \N__49238\ : std_logic;
signal \N__49237\ : std_logic;
signal \N__49236\ : std_logic;
signal \N__49235\ : std_logic;
signal \N__49232\ : std_logic;
signal \N__49229\ : std_logic;
signal \N__49226\ : std_logic;
signal \N__49223\ : std_logic;
signal \N__49220\ : std_logic;
signal \N__49217\ : std_logic;
signal \N__49216\ : std_logic;
signal \N__49215\ : std_logic;
signal \N__49212\ : std_logic;
signal \N__49211\ : std_logic;
signal \N__49210\ : std_logic;
signal \N__49207\ : std_logic;
signal \N__49200\ : std_logic;
signal \N__49193\ : std_logic;
signal \N__49190\ : std_logic;
signal \N__49187\ : std_logic;
signal \N__49186\ : std_logic;
signal \N__49185\ : std_logic;
signal \N__49182\ : std_logic;
signal \N__49179\ : std_logic;
signal \N__49176\ : std_logic;
signal \N__49169\ : std_logic;
signal \N__49164\ : std_logic;
signal \N__49159\ : std_logic;
signal \N__49154\ : std_logic;
signal \N__49147\ : std_logic;
signal \N__49144\ : std_logic;
signal \N__49141\ : std_logic;
signal \N__49140\ : std_logic;
signal \N__49135\ : std_logic;
signal \N__49132\ : std_logic;
signal \N__49129\ : std_logic;
signal \N__49126\ : std_logic;
signal \N__49123\ : std_logic;
signal \N__49120\ : std_logic;
signal \N__49117\ : std_logic;
signal \N__49114\ : std_logic;
signal \N__49113\ : std_logic;
signal \N__49110\ : std_logic;
signal \N__49107\ : std_logic;
signal \N__49102\ : std_logic;
signal \N__49099\ : std_logic;
signal \N__49096\ : std_logic;
signal \N__49093\ : std_logic;
signal \N__49090\ : std_logic;
signal \N__49087\ : std_logic;
signal \N__49084\ : std_logic;
signal \N__49081\ : std_logic;
signal \N__49078\ : std_logic;
signal \N__49077\ : std_logic;
signal \N__49074\ : std_logic;
signal \N__49071\ : std_logic;
signal \N__49070\ : std_logic;
signal \N__49067\ : std_logic;
signal \N__49064\ : std_logic;
signal \N__49061\ : std_logic;
signal \N__49058\ : std_logic;
signal \N__49055\ : std_logic;
signal \N__49048\ : std_logic;
signal \N__49045\ : std_logic;
signal \N__49042\ : std_logic;
signal \N__49041\ : std_logic;
signal \N__49038\ : std_logic;
signal \N__49035\ : std_logic;
signal \N__49032\ : std_logic;
signal \N__49029\ : std_logic;
signal \N__49026\ : std_logic;
signal \N__49025\ : std_logic;
signal \N__49022\ : std_logic;
signal \N__49019\ : std_logic;
signal \N__49016\ : std_logic;
signal \N__49009\ : std_logic;
signal \N__49008\ : std_logic;
signal \N__49005\ : std_logic;
signal \N__49004\ : std_logic;
signal \N__49001\ : std_logic;
signal \N__49000\ : std_logic;
signal \N__48999\ : std_logic;
signal \N__48998\ : std_logic;
signal \N__48997\ : std_logic;
signal \N__48994\ : std_logic;
signal \N__48991\ : std_logic;
signal \N__48990\ : std_logic;
signal \N__48987\ : std_logic;
signal \N__48984\ : std_logic;
signal \N__48979\ : std_logic;
signal \N__48976\ : std_logic;
signal \N__48975\ : std_logic;
signal \N__48970\ : std_logic;
signal \N__48969\ : std_logic;
signal \N__48968\ : std_logic;
signal \N__48967\ : std_logic;
signal \N__48966\ : std_logic;
signal \N__48963\ : std_logic;
signal \N__48962\ : std_logic;
signal \N__48961\ : std_logic;
signal \N__48960\ : std_logic;
signal \N__48959\ : std_logic;
signal \N__48954\ : std_logic;
signal \N__48953\ : std_logic;
signal \N__48948\ : std_logic;
signal \N__48945\ : std_logic;
signal \N__48942\ : std_logic;
signal \N__48939\ : std_logic;
signal \N__48936\ : std_logic;
signal \N__48931\ : std_logic;
signal \N__48928\ : std_logic;
signal \N__48923\ : std_logic;
signal \N__48918\ : std_logic;
signal \N__48915\ : std_logic;
signal \N__48912\ : std_logic;
signal \N__48911\ : std_logic;
signal \N__48910\ : std_logic;
signal \N__48905\ : std_logic;
signal \N__48898\ : std_logic;
signal \N__48895\ : std_logic;
signal \N__48894\ : std_logic;
signal \N__48893\ : std_logic;
signal \N__48892\ : std_logic;
signal \N__48887\ : std_logic;
signal \N__48884\ : std_logic;
signal \N__48879\ : std_logic;
signal \N__48874\ : std_logic;
signal \N__48873\ : std_logic;
signal \N__48870\ : std_logic;
signal \N__48867\ : std_logic;
signal \N__48864\ : std_logic;
signal \N__48859\ : std_logic;
signal \N__48856\ : std_logic;
signal \N__48847\ : std_logic;
signal \N__48844\ : std_logic;
signal \N__48829\ : std_logic;
signal \N__48828\ : std_logic;
signal \N__48825\ : std_logic;
signal \N__48822\ : std_logic;
signal \N__48821\ : std_logic;
signal \N__48818\ : std_logic;
signal \N__48815\ : std_logic;
signal \N__48812\ : std_logic;
signal \N__48809\ : std_logic;
signal \N__48806\ : std_logic;
signal \N__48799\ : std_logic;
signal \N__48798\ : std_logic;
signal \N__48795\ : std_logic;
signal \N__48792\ : std_logic;
signal \N__48789\ : std_logic;
signal \N__48786\ : std_logic;
signal \N__48785\ : std_logic;
signal \N__48782\ : std_logic;
signal \N__48779\ : std_logic;
signal \N__48776\ : std_logic;
signal \N__48769\ : std_logic;
signal \N__48766\ : std_logic;
signal \N__48763\ : std_logic;
signal \N__48760\ : std_logic;
signal \N__48757\ : std_logic;
signal \N__48754\ : std_logic;
signal \N__48751\ : std_logic;
signal \N__48748\ : std_logic;
signal \N__48745\ : std_logic;
signal \N__48744\ : std_logic;
signal \N__48741\ : std_logic;
signal \N__48738\ : std_logic;
signal \N__48737\ : std_logic;
signal \N__48734\ : std_logic;
signal \N__48731\ : std_logic;
signal \N__48728\ : std_logic;
signal \N__48725\ : std_logic;
signal \N__48720\ : std_logic;
signal \N__48717\ : std_logic;
signal \N__48714\ : std_logic;
signal \N__48709\ : std_logic;
signal \N__48706\ : std_logic;
signal \N__48703\ : std_logic;
signal \N__48700\ : std_logic;
signal \N__48699\ : std_logic;
signal \N__48696\ : std_logic;
signal \N__48693\ : std_logic;
signal \N__48688\ : std_logic;
signal \N__48685\ : std_logic;
signal \N__48682\ : std_logic;
signal \N__48681\ : std_logic;
signal \N__48678\ : std_logic;
signal \N__48675\ : std_logic;
signal \N__48672\ : std_logic;
signal \N__48667\ : std_logic;
signal \N__48664\ : std_logic;
signal \N__48663\ : std_logic;
signal \N__48662\ : std_logic;
signal \N__48659\ : std_logic;
signal \N__48656\ : std_logic;
signal \N__48655\ : std_logic;
signal \N__48652\ : std_logic;
signal \N__48649\ : std_logic;
signal \N__48646\ : std_logic;
signal \N__48643\ : std_logic;
signal \N__48640\ : std_logic;
signal \N__48635\ : std_logic;
signal \N__48632\ : std_logic;
signal \N__48631\ : std_logic;
signal \N__48628\ : std_logic;
signal \N__48623\ : std_logic;
signal \N__48620\ : std_logic;
signal \N__48617\ : std_logic;
signal \N__48614\ : std_logic;
signal \N__48611\ : std_logic;
signal \N__48604\ : std_logic;
signal \N__48603\ : std_logic;
signal \N__48600\ : std_logic;
signal \N__48597\ : std_logic;
signal \N__48596\ : std_logic;
signal \N__48593\ : std_logic;
signal \N__48590\ : std_logic;
signal \N__48587\ : std_logic;
signal \N__48586\ : std_logic;
signal \N__48583\ : std_logic;
signal \N__48580\ : std_logic;
signal \N__48577\ : std_logic;
signal \N__48574\ : std_logic;
signal \N__48565\ : std_logic;
signal \N__48564\ : std_logic;
signal \N__48561\ : std_logic;
signal \N__48558\ : std_logic;
signal \N__48557\ : std_logic;
signal \N__48554\ : std_logic;
signal \N__48551\ : std_logic;
signal \N__48548\ : std_logic;
signal \N__48545\ : std_logic;
signal \N__48542\ : std_logic;
signal \N__48535\ : std_logic;
signal \N__48534\ : std_logic;
signal \N__48533\ : std_logic;
signal \N__48530\ : std_logic;
signal \N__48527\ : std_logic;
signal \N__48526\ : std_logic;
signal \N__48525\ : std_logic;
signal \N__48524\ : std_logic;
signal \N__48521\ : std_logic;
signal \N__48518\ : std_logic;
signal \N__48515\ : std_logic;
signal \N__48512\ : std_logic;
signal \N__48511\ : std_logic;
signal \N__48510\ : std_logic;
signal \N__48509\ : std_logic;
signal \N__48508\ : std_logic;
signal \N__48507\ : std_logic;
signal \N__48506\ : std_logic;
signal \N__48505\ : std_logic;
signal \N__48504\ : std_logic;
signal \N__48499\ : std_logic;
signal \N__48496\ : std_logic;
signal \N__48495\ : std_logic;
signal \N__48494\ : std_logic;
signal \N__48493\ : std_logic;
signal \N__48492\ : std_logic;
signal \N__48489\ : std_logic;
signal \N__48484\ : std_logic;
signal \N__48481\ : std_logic;
signal \N__48480\ : std_logic;
signal \N__48479\ : std_logic;
signal \N__48478\ : std_logic;
signal \N__48469\ : std_logic;
signal \N__48464\ : std_logic;
signal \N__48461\ : std_logic;
signal \N__48456\ : std_logic;
signal \N__48453\ : std_logic;
signal \N__48448\ : std_logic;
signal \N__48445\ : std_logic;
signal \N__48440\ : std_logic;
signal \N__48439\ : std_logic;
signal \N__48438\ : std_logic;
signal \N__48437\ : std_logic;
signal \N__48432\ : std_logic;
signal \N__48427\ : std_logic;
signal \N__48422\ : std_logic;
signal \N__48419\ : std_logic;
signal \N__48416\ : std_logic;
signal \N__48413\ : std_logic;
signal \N__48408\ : std_logic;
signal \N__48405\ : std_logic;
signal \N__48402\ : std_logic;
signal \N__48399\ : std_logic;
signal \N__48396\ : std_logic;
signal \N__48389\ : std_logic;
signal \N__48386\ : std_logic;
signal \N__48383\ : std_logic;
signal \N__48378\ : std_logic;
signal \N__48375\ : std_logic;
signal \N__48358\ : std_logic;
signal \N__48355\ : std_logic;
signal \N__48352\ : std_logic;
signal \N__48351\ : std_logic;
signal \N__48350\ : std_logic;
signal \N__48349\ : std_logic;
signal \N__48348\ : std_logic;
signal \N__48347\ : std_logic;
signal \N__48346\ : std_logic;
signal \N__48343\ : std_logic;
signal \N__48336\ : std_logic;
signal \N__48335\ : std_logic;
signal \N__48332\ : std_logic;
signal \N__48329\ : std_logic;
signal \N__48326\ : std_logic;
signal \N__48325\ : std_logic;
signal \N__48324\ : std_logic;
signal \N__48323\ : std_logic;
signal \N__48322\ : std_logic;
signal \N__48321\ : std_logic;
signal \N__48320\ : std_logic;
signal \N__48319\ : std_logic;
signal \N__48316\ : std_logic;
signal \N__48315\ : std_logic;
signal \N__48314\ : std_logic;
signal \N__48311\ : std_logic;
signal \N__48308\ : std_logic;
signal \N__48305\ : std_logic;
signal \N__48302\ : std_logic;
signal \N__48293\ : std_logic;
signal \N__48288\ : std_logic;
signal \N__48287\ : std_logic;
signal \N__48286\ : std_logic;
signal \N__48285\ : std_logic;
signal \N__48284\ : std_logic;
signal \N__48283\ : std_logic;
signal \N__48282\ : std_logic;
signal \N__48281\ : std_logic;
signal \N__48280\ : std_logic;
signal \N__48275\ : std_logic;
signal \N__48272\ : std_logic;
signal \N__48269\ : std_logic;
signal \N__48266\ : std_logic;
signal \N__48265\ : std_logic;
signal \N__48264\ : std_logic;
signal \N__48263\ : std_logic;
signal \N__48262\ : std_logic;
signal \N__48259\ : std_logic;
signal \N__48256\ : std_logic;
signal \N__48251\ : std_logic;
signal \N__48248\ : std_logic;
signal \N__48245\ : std_logic;
signal \N__48242\ : std_logic;
signal \N__48235\ : std_logic;
signal \N__48232\ : std_logic;
signal \N__48229\ : std_logic;
signal \N__48226\ : std_logic;
signal \N__48225\ : std_logic;
signal \N__48224\ : std_logic;
signal \N__48223\ : std_logic;
signal \N__48220\ : std_logic;
signal \N__48219\ : std_logic;
signal \N__48218\ : std_logic;
signal \N__48217\ : std_logic;
signal \N__48216\ : std_logic;
signal \N__48209\ : std_logic;
signal \N__48206\ : std_logic;
signal \N__48205\ : std_logic;
signal \N__48204\ : std_logic;
signal \N__48203\ : std_logic;
signal \N__48202\ : std_logic;
signal \N__48199\ : std_logic;
signal \N__48198\ : std_logic;
signal \N__48197\ : std_logic;
signal \N__48196\ : std_logic;
signal \N__48195\ : std_logic;
signal \N__48194\ : std_logic;
signal \N__48191\ : std_logic;
signal \N__48188\ : std_logic;
signal \N__48185\ : std_logic;
signal \N__48184\ : std_logic;
signal \N__48183\ : std_logic;
signal \N__48182\ : std_logic;
signal \N__48181\ : std_logic;
signal \N__48180\ : std_logic;
signal \N__48179\ : std_logic;
signal \N__48178\ : std_logic;
signal \N__48177\ : std_logic;
signal \N__48176\ : std_logic;
signal \N__48175\ : std_logic;
signal \N__48174\ : std_logic;
signal \N__48173\ : std_logic;
signal \N__48166\ : std_logic;
signal \N__48157\ : std_logic;
signal \N__48144\ : std_logic;
signal \N__48139\ : std_logic;
signal \N__48136\ : std_logic;
signal \N__48131\ : std_logic;
signal \N__48128\ : std_logic;
signal \N__48125\ : std_logic;
signal \N__48118\ : std_logic;
signal \N__48117\ : std_logic;
signal \N__48114\ : std_logic;
signal \N__48113\ : std_logic;
signal \N__48112\ : std_logic;
signal \N__48109\ : std_logic;
signal \N__48098\ : std_logic;
signal \N__48081\ : std_logic;
signal \N__48076\ : std_logic;
signal \N__48065\ : std_logic;
signal \N__48060\ : std_logic;
signal \N__48051\ : std_logic;
signal \N__48048\ : std_logic;
signal \N__48043\ : std_logic;
signal \N__48042\ : std_logic;
signal \N__48041\ : std_logic;
signal \N__48040\ : std_logic;
signal \N__48039\ : std_logic;
signal \N__48038\ : std_logic;
signal \N__48037\ : std_logic;
signal \N__48036\ : std_logic;
signal \N__48035\ : std_logic;
signal \N__48032\ : std_logic;
signal \N__48025\ : std_logic;
signal \N__48018\ : std_logic;
signal \N__48013\ : std_logic;
signal \N__48010\ : std_logic;
signal \N__48003\ : std_logic;
signal \N__47994\ : std_logic;
signal \N__47985\ : std_logic;
signal \N__47968\ : std_logic;
signal \N__47967\ : std_logic;
signal \N__47964\ : std_logic;
signal \N__47961\ : std_logic;
signal \N__47958\ : std_logic;
signal \N__47955\ : std_logic;
signal \N__47952\ : std_logic;
signal \N__47949\ : std_logic;
signal \N__47948\ : std_logic;
signal \N__47945\ : std_logic;
signal \N__47942\ : std_logic;
signal \N__47939\ : std_logic;
signal \N__47932\ : std_logic;
signal \N__47929\ : std_logic;
signal \N__47928\ : std_logic;
signal \N__47925\ : std_logic;
signal \N__47924\ : std_logic;
signal \N__47921\ : std_logic;
signal \N__47918\ : std_logic;
signal \N__47915\ : std_logic;
signal \N__47908\ : std_logic;
signal \N__47905\ : std_logic;
signal \N__47902\ : std_logic;
signal \N__47899\ : std_logic;
signal \N__47898\ : std_logic;
signal \N__47895\ : std_logic;
signal \N__47892\ : std_logic;
signal \N__47889\ : std_logic;
signal \N__47886\ : std_logic;
signal \N__47881\ : std_logic;
signal \N__47880\ : std_logic;
signal \N__47877\ : std_logic;
signal \N__47874\ : std_logic;
signal \N__47873\ : std_logic;
signal \N__47870\ : std_logic;
signal \N__47867\ : std_logic;
signal \N__47864\ : std_logic;
signal \N__47861\ : std_logic;
signal \N__47854\ : std_logic;
signal \N__47851\ : std_logic;
signal \N__47850\ : std_logic;
signal \N__47849\ : std_logic;
signal \N__47848\ : std_logic;
signal \N__47847\ : std_logic;
signal \N__47846\ : std_logic;
signal \N__47845\ : std_logic;
signal \N__47844\ : std_logic;
signal \N__47843\ : std_logic;
signal \N__47840\ : std_logic;
signal \N__47837\ : std_logic;
signal \N__47836\ : std_logic;
signal \N__47835\ : std_logic;
signal \N__47834\ : std_logic;
signal \N__47833\ : std_logic;
signal \N__47832\ : std_logic;
signal \N__47831\ : std_logic;
signal \N__47830\ : std_logic;
signal \N__47829\ : std_logic;
signal \N__47826\ : std_logic;
signal \N__47825\ : std_logic;
signal \N__47824\ : std_logic;
signal \N__47823\ : std_logic;
signal \N__47822\ : std_logic;
signal \N__47821\ : std_logic;
signal \N__47820\ : std_logic;
signal \N__47817\ : std_logic;
signal \N__47814\ : std_logic;
signal \N__47811\ : std_logic;
signal \N__47806\ : std_logic;
signal \N__47803\ : std_logic;
signal \N__47800\ : std_logic;
signal \N__47797\ : std_logic;
signal \N__47794\ : std_logic;
signal \N__47791\ : std_logic;
signal \N__47790\ : std_logic;
signal \N__47789\ : std_logic;
signal \N__47788\ : std_logic;
signal \N__47787\ : std_logic;
signal \N__47786\ : std_logic;
signal \N__47785\ : std_logic;
signal \N__47784\ : std_logic;
signal \N__47783\ : std_logic;
signal \N__47782\ : std_logic;
signal \N__47781\ : std_logic;
signal \N__47780\ : std_logic;
signal \N__47779\ : std_logic;
signal \N__47778\ : std_logic;
signal \N__47775\ : std_logic;
signal \N__47774\ : std_logic;
signal \N__47771\ : std_logic;
signal \N__47768\ : std_logic;
signal \N__47763\ : std_logic;
signal \N__47758\ : std_logic;
signal \N__47755\ : std_logic;
signal \N__47754\ : std_logic;
signal \N__47753\ : std_logic;
signal \N__47752\ : std_logic;
signal \N__47749\ : std_logic;
signal \N__47748\ : std_logic;
signal \N__47747\ : std_logic;
signal \N__47746\ : std_logic;
signal \N__47745\ : std_logic;
signal \N__47744\ : std_logic;
signal \N__47743\ : std_logic;
signal \N__47742\ : std_logic;
signal \N__47741\ : std_logic;
signal \N__47738\ : std_logic;
signal \N__47737\ : std_logic;
signal \N__47734\ : std_logic;
signal \N__47731\ : std_logic;
signal \N__47728\ : std_logic;
signal \N__47727\ : std_logic;
signal \N__47726\ : std_logic;
signal \N__47721\ : std_logic;
signal \N__47718\ : std_logic;
signal \N__47705\ : std_logic;
signal \N__47702\ : std_logic;
signal \N__47701\ : std_logic;
signal \N__47700\ : std_logic;
signal \N__47699\ : std_logic;
signal \N__47698\ : std_logic;
signal \N__47697\ : std_logic;
signal \N__47696\ : std_logic;
signal \N__47695\ : std_logic;
signal \N__47694\ : std_logic;
signal \N__47691\ : std_logic;
signal \N__47688\ : std_logic;
signal \N__47683\ : std_logic;
signal \N__47674\ : std_logic;
signal \N__47665\ : std_logic;
signal \N__47662\ : std_logic;
signal \N__47659\ : std_logic;
signal \N__47654\ : std_logic;
signal \N__47649\ : std_logic;
signal \N__47646\ : std_logic;
signal \N__47643\ : std_logic;
signal \N__47640\ : std_logic;
signal \N__47637\ : std_logic;
signal \N__47634\ : std_logic;
signal \N__47631\ : std_logic;
signal \N__47628\ : std_logic;
signal \N__47623\ : std_logic;
signal \N__47618\ : std_logic;
signal \N__47615\ : std_logic;
signal \N__47612\ : std_logic;
signal \N__47609\ : std_logic;
signal \N__47606\ : std_logic;
signal \N__47601\ : std_logic;
signal \N__47598\ : std_logic;
signal \N__47593\ : std_logic;
signal \N__47584\ : std_logic;
signal \N__47581\ : std_logic;
signal \N__47580\ : std_logic;
signal \N__47579\ : std_logic;
signal \N__47578\ : std_logic;
signal \N__47573\ : std_logic;
signal \N__47568\ : std_logic;
signal \N__47565\ : std_logic;
signal \N__47562\ : std_logic;
signal \N__47559\ : std_logic;
signal \N__47556\ : std_logic;
signal \N__47545\ : std_logic;
signal \N__47542\ : std_logic;
signal \N__47533\ : std_logic;
signal \N__47520\ : std_logic;
signal \N__47509\ : std_logic;
signal \N__47508\ : std_logic;
signal \N__47503\ : std_logic;
signal \N__47498\ : std_logic;
signal \N__47495\ : std_logic;
signal \N__47488\ : std_logic;
signal \N__47479\ : std_logic;
signal \N__47464\ : std_logic;
signal \N__47461\ : std_logic;
signal \N__47456\ : std_logic;
signal \N__47443\ : std_logic;
signal \N__47440\ : std_logic;
signal \N__47437\ : std_logic;
signal \N__47434\ : std_logic;
signal \N__47431\ : std_logic;
signal \N__47428\ : std_logic;
signal \N__47425\ : std_logic;
signal \N__47422\ : std_logic;
signal \N__47419\ : std_logic;
signal \N__47416\ : std_logic;
signal \N__47413\ : std_logic;
signal \N__47412\ : std_logic;
signal \N__47409\ : std_logic;
signal \N__47406\ : std_logic;
signal \N__47403\ : std_logic;
signal \N__47402\ : std_logic;
signal \N__47399\ : std_logic;
signal \N__47396\ : std_logic;
signal \N__47393\ : std_logic;
signal \N__47390\ : std_logic;
signal \N__47387\ : std_logic;
signal \N__47380\ : std_logic;
signal \N__47377\ : std_logic;
signal \N__47376\ : std_logic;
signal \N__47373\ : std_logic;
signal \N__47370\ : std_logic;
signal \N__47369\ : std_logic;
signal \N__47366\ : std_logic;
signal \N__47363\ : std_logic;
signal \N__47360\ : std_logic;
signal \N__47357\ : std_logic;
signal \N__47354\ : std_logic;
signal \N__47347\ : std_logic;
signal \N__47344\ : std_logic;
signal \N__47343\ : std_logic;
signal \N__47340\ : std_logic;
signal \N__47337\ : std_logic;
signal \N__47336\ : std_logic;
signal \N__47333\ : std_logic;
signal \N__47330\ : std_logic;
signal \N__47327\ : std_logic;
signal \N__47324\ : std_logic;
signal \N__47321\ : std_logic;
signal \N__47314\ : std_logic;
signal \N__47311\ : std_logic;
signal \N__47308\ : std_logic;
signal \N__47307\ : std_logic;
signal \N__47304\ : std_logic;
signal \N__47301\ : std_logic;
signal \N__47298\ : std_logic;
signal \N__47297\ : std_logic;
signal \N__47292\ : std_logic;
signal \N__47289\ : std_logic;
signal \N__47286\ : std_logic;
signal \N__47281\ : std_logic;
signal \N__47278\ : std_logic;
signal \N__47275\ : std_logic;
signal \N__47274\ : std_logic;
signal \N__47271\ : std_logic;
signal \N__47268\ : std_logic;
signal \N__47267\ : std_logic;
signal \N__47264\ : std_logic;
signal \N__47261\ : std_logic;
signal \N__47258\ : std_logic;
signal \N__47255\ : std_logic;
signal \N__47252\ : std_logic;
signal \N__47245\ : std_logic;
signal \N__47242\ : std_logic;
signal \N__47241\ : std_logic;
signal \N__47240\ : std_logic;
signal \N__47237\ : std_logic;
signal \N__47234\ : std_logic;
signal \N__47231\ : std_logic;
signal \N__47224\ : std_logic;
signal \N__47221\ : std_logic;
signal \N__47218\ : std_logic;
signal \N__47217\ : std_logic;
signal \N__47214\ : std_logic;
signal \N__47211\ : std_logic;
signal \N__47208\ : std_logic;
signal \N__47203\ : std_logic;
signal \N__47200\ : std_logic;
signal \N__47197\ : std_logic;
signal \N__47196\ : std_logic;
signal \N__47193\ : std_logic;
signal \N__47190\ : std_logic;
signal \N__47187\ : std_logic;
signal \N__47182\ : std_logic;
signal \N__47179\ : std_logic;
signal \N__47176\ : std_logic;
signal \N__47173\ : std_logic;
signal \N__47172\ : std_logic;
signal \N__47169\ : std_logic;
signal \N__47166\ : std_logic;
signal \N__47163\ : std_logic;
signal \N__47158\ : std_logic;
signal \N__47155\ : std_logic;
signal \N__47152\ : std_logic;
signal \N__47149\ : std_logic;
signal \N__47146\ : std_logic;
signal \N__47143\ : std_logic;
signal \N__47140\ : std_logic;
signal \N__47137\ : std_logic;
signal \N__47136\ : std_logic;
signal \N__47135\ : std_logic;
signal \N__47132\ : std_logic;
signal \N__47129\ : std_logic;
signal \N__47128\ : std_logic;
signal \N__47125\ : std_logic;
signal \N__47124\ : std_logic;
signal \N__47119\ : std_logic;
signal \N__47116\ : std_logic;
signal \N__47113\ : std_logic;
signal \N__47110\ : std_logic;
signal \N__47105\ : std_logic;
signal \N__47104\ : std_logic;
signal \N__47101\ : std_logic;
signal \N__47098\ : std_logic;
signal \N__47095\ : std_logic;
signal \N__47092\ : std_logic;
signal \N__47085\ : std_logic;
signal \N__47082\ : std_logic;
signal \N__47081\ : std_logic;
signal \N__47078\ : std_logic;
signal \N__47075\ : std_logic;
signal \N__47072\ : std_logic;
signal \N__47065\ : std_logic;
signal \N__47062\ : std_logic;
signal \N__47061\ : std_logic;
signal \N__47058\ : std_logic;
signal \N__47057\ : std_logic;
signal \N__47056\ : std_logic;
signal \N__47053\ : std_logic;
signal \N__47052\ : std_logic;
signal \N__47049\ : std_logic;
signal \N__47048\ : std_logic;
signal \N__47045\ : std_logic;
signal \N__47042\ : std_logic;
signal \N__47039\ : std_logic;
signal \N__47036\ : std_logic;
signal \N__47033\ : std_logic;
signal \N__47030\ : std_logic;
signal \N__47027\ : std_logic;
signal \N__47024\ : std_logic;
signal \N__47019\ : std_logic;
signal \N__47014\ : std_logic;
signal \N__47011\ : std_logic;
signal \N__47006\ : std_logic;
signal \N__47003\ : std_logic;
signal \N__46996\ : std_logic;
signal \N__46993\ : std_logic;
signal \N__46990\ : std_logic;
signal \N__46987\ : std_logic;
signal \N__46986\ : std_logic;
signal \N__46983\ : std_logic;
signal \N__46980\ : std_logic;
signal \N__46977\ : std_logic;
signal \N__46976\ : std_logic;
signal \N__46975\ : std_logic;
signal \N__46972\ : std_logic;
signal \N__46969\ : std_logic;
signal \N__46968\ : std_logic;
signal \N__46963\ : std_logic;
signal \N__46960\ : std_logic;
signal \N__46957\ : std_logic;
signal \N__46956\ : std_logic;
signal \N__46953\ : std_logic;
signal \N__46946\ : std_logic;
signal \N__46943\ : std_logic;
signal \N__46936\ : std_logic;
signal \N__46935\ : std_logic;
signal \N__46932\ : std_logic;
signal \N__46929\ : std_logic;
signal \N__46928\ : std_logic;
signal \N__46923\ : std_logic;
signal \N__46920\ : std_logic;
signal \N__46917\ : std_logic;
signal \N__46912\ : std_logic;
signal \N__46909\ : std_logic;
signal \N__46908\ : std_logic;
signal \N__46907\ : std_logic;
signal \N__46904\ : std_logic;
signal \N__46901\ : std_logic;
signal \N__46898\ : std_logic;
signal \N__46895\ : std_logic;
signal \N__46892\ : std_logic;
signal \N__46885\ : std_logic;
signal \N__46882\ : std_logic;
signal \N__46881\ : std_logic;
signal \N__46878\ : std_logic;
signal \N__46875\ : std_logic;
signal \N__46872\ : std_logic;
signal \N__46871\ : std_logic;
signal \N__46866\ : std_logic;
signal \N__46863\ : std_logic;
signal \N__46860\ : std_logic;
signal \N__46855\ : std_logic;
signal \N__46852\ : std_logic;
signal \N__46851\ : std_logic;
signal \N__46848\ : std_logic;
signal \N__46845\ : std_logic;
signal \N__46842\ : std_logic;
signal \N__46839\ : std_logic;
signal \N__46838\ : std_logic;
signal \N__46835\ : std_logic;
signal \N__46832\ : std_logic;
signal \N__46829\ : std_logic;
signal \N__46826\ : std_logic;
signal \N__46823\ : std_logic;
signal \N__46816\ : std_logic;
signal \N__46813\ : std_logic;
signal \N__46812\ : std_logic;
signal \N__46809\ : std_logic;
signal \N__46806\ : std_logic;
signal \N__46803\ : std_logic;
signal \N__46802\ : std_logic;
signal \N__46797\ : std_logic;
signal \N__46794\ : std_logic;
signal \N__46791\ : std_logic;
signal \N__46786\ : std_logic;
signal \N__46783\ : std_logic;
signal \N__46782\ : std_logic;
signal \N__46779\ : std_logic;
signal \N__46776\ : std_logic;
signal \N__46773\ : std_logic;
signal \N__46772\ : std_logic;
signal \N__46767\ : std_logic;
signal \N__46764\ : std_logic;
signal \N__46761\ : std_logic;
signal \N__46756\ : std_logic;
signal \N__46753\ : std_logic;
signal \N__46750\ : std_logic;
signal \N__46747\ : std_logic;
signal \N__46744\ : std_logic;
signal \N__46741\ : std_logic;
signal \N__46738\ : std_logic;
signal \N__46735\ : std_logic;
signal \N__46734\ : std_logic;
signal \N__46731\ : std_logic;
signal \N__46728\ : std_logic;
signal \N__46725\ : std_logic;
signal \N__46720\ : std_logic;
signal \N__46717\ : std_logic;
signal \N__46714\ : std_logic;
signal \N__46711\ : std_logic;
signal \N__46708\ : std_logic;
signal \N__46707\ : std_logic;
signal \N__46704\ : std_logic;
signal \N__46701\ : std_logic;
signal \N__46700\ : std_logic;
signal \N__46697\ : std_logic;
signal \N__46694\ : std_logic;
signal \N__46691\ : std_logic;
signal \N__46688\ : std_logic;
signal \N__46683\ : std_logic;
signal \N__46680\ : std_logic;
signal \N__46677\ : std_logic;
signal \N__46674\ : std_logic;
signal \N__46671\ : std_logic;
signal \N__46666\ : std_logic;
signal \N__46665\ : std_logic;
signal \N__46664\ : std_logic;
signal \N__46661\ : std_logic;
signal \N__46658\ : std_logic;
signal \N__46655\ : std_logic;
signal \N__46654\ : std_logic;
signal \N__46651\ : std_logic;
signal \N__46648\ : std_logic;
signal \N__46647\ : std_logic;
signal \N__46646\ : std_logic;
signal \N__46643\ : std_logic;
signal \N__46640\ : std_logic;
signal \N__46637\ : std_logic;
signal \N__46634\ : std_logic;
signal \N__46631\ : std_logic;
signal \N__46628\ : std_logic;
signal \N__46625\ : std_logic;
signal \N__46622\ : std_logic;
signal \N__46619\ : std_logic;
signal \N__46614\ : std_logic;
signal \N__46611\ : std_logic;
signal \N__46606\ : std_logic;
signal \N__46597\ : std_logic;
signal \N__46594\ : std_logic;
signal \N__46591\ : std_logic;
signal \N__46588\ : std_logic;
signal \N__46585\ : std_logic;
signal \N__46582\ : std_logic;
signal \N__46581\ : std_logic;
signal \N__46578\ : std_logic;
signal \N__46575\ : std_logic;
signal \N__46570\ : std_logic;
signal \N__46567\ : std_logic;
signal \N__46564\ : std_logic;
signal \N__46561\ : std_logic;
signal \N__46558\ : std_logic;
signal \N__46555\ : std_logic;
signal \N__46552\ : std_logic;
signal \N__46549\ : std_logic;
signal \N__46546\ : std_logic;
signal \N__46543\ : std_logic;
signal \N__46540\ : std_logic;
signal \N__46537\ : std_logic;
signal \N__46534\ : std_logic;
signal \N__46531\ : std_logic;
signal \N__46528\ : std_logic;
signal \N__46525\ : std_logic;
signal \N__46522\ : std_logic;
signal \N__46519\ : std_logic;
signal \N__46516\ : std_logic;
signal \N__46513\ : std_logic;
signal \N__46510\ : std_logic;
signal \N__46507\ : std_logic;
signal \N__46504\ : std_logic;
signal \N__46501\ : std_logic;
signal \N__46500\ : std_logic;
signal \N__46497\ : std_logic;
signal \N__46494\ : std_logic;
signal \N__46491\ : std_logic;
signal \N__46488\ : std_logic;
signal \N__46483\ : std_logic;
signal \N__46480\ : std_logic;
signal \N__46477\ : std_logic;
signal \N__46474\ : std_logic;
signal \N__46471\ : std_logic;
signal \N__46468\ : std_logic;
signal \N__46467\ : std_logic;
signal \N__46462\ : std_logic;
signal \N__46459\ : std_logic;
signal \N__46456\ : std_logic;
signal \N__46453\ : std_logic;
signal \N__46450\ : std_logic;
signal \N__46447\ : std_logic;
signal \N__46444\ : std_logic;
signal \N__46441\ : std_logic;
signal \N__46438\ : std_logic;
signal \N__46435\ : std_logic;
signal \N__46432\ : std_logic;
signal \N__46429\ : std_logic;
signal \N__46426\ : std_logic;
signal \N__46423\ : std_logic;
signal \N__46422\ : std_logic;
signal \N__46419\ : std_logic;
signal \N__46416\ : std_logic;
signal \N__46413\ : std_logic;
signal \N__46408\ : std_logic;
signal \N__46405\ : std_logic;
signal \N__46402\ : std_logic;
signal \N__46399\ : std_logic;
signal \N__46398\ : std_logic;
signal \N__46395\ : std_logic;
signal \N__46392\ : std_logic;
signal \N__46387\ : std_logic;
signal \N__46384\ : std_logic;
signal \N__46381\ : std_logic;
signal \N__46378\ : std_logic;
signal \N__46377\ : std_logic;
signal \N__46376\ : std_logic;
signal \N__46375\ : std_logic;
signal \N__46374\ : std_logic;
signal \N__46373\ : std_logic;
signal \N__46372\ : std_logic;
signal \N__46371\ : std_logic;
signal \N__46370\ : std_logic;
signal \N__46367\ : std_logic;
signal \N__46364\ : std_logic;
signal \N__46349\ : std_logic;
signal \N__46342\ : std_logic;
signal \N__46339\ : std_logic;
signal \N__46336\ : std_logic;
signal \N__46333\ : std_logic;
signal \N__46332\ : std_logic;
signal \N__46331\ : std_logic;
signal \N__46330\ : std_logic;
signal \N__46329\ : std_logic;
signal \N__46328\ : std_logic;
signal \N__46327\ : std_logic;
signal \N__46326\ : std_logic;
signal \N__46323\ : std_logic;
signal \N__46308\ : std_logic;
signal \N__46303\ : std_logic;
signal \N__46300\ : std_logic;
signal \N__46297\ : std_logic;
signal \N__46294\ : std_logic;
signal \N__46293\ : std_logic;
signal \N__46290\ : std_logic;
signal \N__46287\ : std_logic;
signal \N__46282\ : std_logic;
signal \N__46279\ : std_logic;
signal \N__46276\ : std_logic;
signal \N__46273\ : std_logic;
signal \N__46270\ : std_logic;
signal \N__46269\ : std_logic;
signal \N__46266\ : std_logic;
signal \N__46263\ : std_logic;
signal \N__46258\ : std_logic;
signal \N__46257\ : std_logic;
signal \N__46254\ : std_logic;
signal \N__46251\ : std_logic;
signal \N__46246\ : std_logic;
signal \N__46243\ : std_logic;
signal \N__46242\ : std_logic;
signal \N__46239\ : std_logic;
signal \N__46236\ : std_logic;
signal \N__46231\ : std_logic;
signal \N__46228\ : std_logic;
signal \N__46227\ : std_logic;
signal \N__46224\ : std_logic;
signal \N__46221\ : std_logic;
signal \N__46216\ : std_logic;
signal \N__46213\ : std_logic;
signal \N__46210\ : std_logic;
signal \N__46207\ : std_logic;
signal \N__46206\ : std_logic;
signal \N__46203\ : std_logic;
signal \N__46200\ : std_logic;
signal \N__46195\ : std_logic;
signal \N__46192\ : std_logic;
signal \N__46191\ : std_logic;
signal \N__46188\ : std_logic;
signal \N__46185\ : std_logic;
signal \N__46180\ : std_logic;
signal \N__46179\ : std_logic;
signal \N__46176\ : std_logic;
signal \N__46173\ : std_logic;
signal \N__46168\ : std_logic;
signal \N__46165\ : std_logic;
signal \N__46162\ : std_logic;
signal \N__46159\ : std_logic;
signal \N__46156\ : std_logic;
signal \N__46155\ : std_logic;
signal \N__46152\ : std_logic;
signal \N__46149\ : std_logic;
signal \N__46146\ : std_logic;
signal \N__46143\ : std_logic;
signal \N__46138\ : std_logic;
signal \N__46137\ : std_logic;
signal \N__46134\ : std_logic;
signal \N__46131\ : std_logic;
signal \N__46128\ : std_logic;
signal \N__46125\ : std_logic;
signal \N__46120\ : std_logic;
signal \N__46117\ : std_logic;
signal \N__46114\ : std_logic;
signal \N__46111\ : std_logic;
signal \N__46108\ : std_logic;
signal \N__46105\ : std_logic;
signal \N__46102\ : std_logic;
signal \N__46099\ : std_logic;
signal \N__46096\ : std_logic;
signal \N__46093\ : std_logic;
signal \N__46090\ : std_logic;
signal \N__46087\ : std_logic;
signal \N__46084\ : std_logic;
signal \N__46081\ : std_logic;
signal \N__46078\ : std_logic;
signal \N__46077\ : std_logic;
signal \N__46074\ : std_logic;
signal \N__46071\ : std_logic;
signal \N__46066\ : std_logic;
signal \N__46063\ : std_logic;
signal \N__46060\ : std_logic;
signal \N__46057\ : std_logic;
signal \N__46054\ : std_logic;
signal \N__46053\ : std_logic;
signal \N__46050\ : std_logic;
signal \N__46047\ : std_logic;
signal \N__46042\ : std_logic;
signal \N__46039\ : std_logic;
signal \N__46038\ : std_logic;
signal \N__46037\ : std_logic;
signal \N__46034\ : std_logic;
signal \N__46031\ : std_logic;
signal \N__46028\ : std_logic;
signal \N__46021\ : std_logic;
signal \N__46020\ : std_logic;
signal \N__46019\ : std_logic;
signal \N__46018\ : std_logic;
signal \N__46017\ : std_logic;
signal \N__46016\ : std_logic;
signal \N__46015\ : std_logic;
signal \N__46014\ : std_logic;
signal \N__46013\ : std_logic;
signal \N__46010\ : std_logic;
signal \N__46007\ : std_logic;
signal \N__46006\ : std_logic;
signal \N__46005\ : std_logic;
signal \N__45994\ : std_logic;
signal \N__45991\ : std_logic;
signal \N__45988\ : std_logic;
signal \N__45987\ : std_logic;
signal \N__45982\ : std_logic;
signal \N__45977\ : std_logic;
signal \N__45974\ : std_logic;
signal \N__45969\ : std_logic;
signal \N__45966\ : std_logic;
signal \N__45965\ : std_logic;
signal \N__45960\ : std_logic;
signal \N__45953\ : std_logic;
signal \N__45950\ : std_logic;
signal \N__45947\ : std_logic;
signal \N__45942\ : std_logic;
signal \N__45937\ : std_logic;
signal \N__45934\ : std_logic;
signal \N__45933\ : std_logic;
signal \N__45930\ : std_logic;
signal \N__45927\ : std_logic;
signal \N__45924\ : std_logic;
signal \N__45921\ : std_logic;
signal \N__45916\ : std_logic;
signal \N__45915\ : std_logic;
signal \N__45914\ : std_logic;
signal \N__45913\ : std_logic;
signal \N__45912\ : std_logic;
signal \N__45911\ : std_logic;
signal \N__45908\ : std_logic;
signal \N__45905\ : std_logic;
signal \N__45902\ : std_logic;
signal \N__45901\ : std_logic;
signal \N__45900\ : std_logic;
signal \N__45897\ : std_logic;
signal \N__45896\ : std_logic;
signal \N__45895\ : std_logic;
signal \N__45892\ : std_logic;
signal \N__45891\ : std_logic;
signal \N__45888\ : std_logic;
signal \N__45877\ : std_logic;
signal \N__45876\ : std_logic;
signal \N__45871\ : std_logic;
signal \N__45868\ : std_logic;
signal \N__45865\ : std_logic;
signal \N__45862\ : std_logic;
signal \N__45859\ : std_logic;
signal \N__45856\ : std_logic;
signal \N__45853\ : std_logic;
signal \N__45850\ : std_logic;
signal \N__45847\ : std_logic;
signal \N__45844\ : std_logic;
signal \N__45841\ : std_logic;
signal \N__45840\ : std_logic;
signal \N__45839\ : std_logic;
signal \N__45838\ : std_logic;
signal \N__45835\ : std_logic;
signal \N__45830\ : std_logic;
signal \N__45829\ : std_logic;
signal \N__45822\ : std_logic;
signal \N__45819\ : std_logic;
signal \N__45816\ : std_logic;
signal \N__45811\ : std_logic;
signal \N__45810\ : std_logic;
signal \N__45807\ : std_logic;
signal \N__45804\ : std_logic;
signal \N__45801\ : std_logic;
signal \N__45798\ : std_logic;
signal \N__45795\ : std_logic;
signal \N__45790\ : std_logic;
signal \N__45787\ : std_logic;
signal \N__45772\ : std_logic;
signal \N__45769\ : std_logic;
signal \N__45768\ : std_logic;
signal \N__45767\ : std_logic;
signal \N__45766\ : std_logic;
signal \N__45765\ : std_logic;
signal \N__45762\ : std_logic;
signal \N__45759\ : std_logic;
signal \N__45756\ : std_logic;
signal \N__45753\ : std_logic;
signal \N__45750\ : std_logic;
signal \N__45747\ : std_logic;
signal \N__45744\ : std_logic;
signal \N__45741\ : std_logic;
signal \N__45738\ : std_logic;
signal \N__45735\ : std_logic;
signal \N__45728\ : std_logic;
signal \N__45727\ : std_logic;
signal \N__45724\ : std_logic;
signal \N__45721\ : std_logic;
signal \N__45718\ : std_logic;
signal \N__45715\ : std_logic;
signal \N__45712\ : std_logic;
signal \N__45709\ : std_logic;
signal \N__45706\ : std_logic;
signal \N__45697\ : std_logic;
signal \N__45696\ : std_logic;
signal \N__45695\ : std_logic;
signal \N__45694\ : std_logic;
signal \N__45693\ : std_logic;
signal \N__45692\ : std_logic;
signal \N__45691\ : std_logic;
signal \N__45688\ : std_logic;
signal \N__45681\ : std_logic;
signal \N__45678\ : std_logic;
signal \N__45677\ : std_logic;
signal \N__45676\ : std_logic;
signal \N__45675\ : std_logic;
signal \N__45674\ : std_logic;
signal \N__45673\ : std_logic;
signal \N__45668\ : std_logic;
signal \N__45661\ : std_logic;
signal \N__45658\ : std_logic;
signal \N__45657\ : std_logic;
signal \N__45656\ : std_logic;
signal \N__45655\ : std_logic;
signal \N__45650\ : std_logic;
signal \N__45647\ : std_logic;
signal \N__45644\ : std_logic;
signal \N__45641\ : std_logic;
signal \N__45638\ : std_logic;
signal \N__45635\ : std_logic;
signal \N__45632\ : std_logic;
signal \N__45629\ : std_logic;
signal \N__45626\ : std_logic;
signal \N__45621\ : std_logic;
signal \N__45616\ : std_logic;
signal \N__45611\ : std_logic;
signal \N__45608\ : std_logic;
signal \N__45595\ : std_logic;
signal \N__45592\ : std_logic;
signal \N__45591\ : std_logic;
signal \N__45588\ : std_logic;
signal \N__45585\ : std_logic;
signal \N__45582\ : std_logic;
signal \N__45581\ : std_logic;
signal \N__45578\ : std_logic;
signal \N__45575\ : std_logic;
signal \N__45572\ : std_logic;
signal \N__45567\ : std_logic;
signal \N__45562\ : std_logic;
signal \N__45561\ : std_logic;
signal \N__45558\ : std_logic;
signal \N__45555\ : std_logic;
signal \N__45552\ : std_logic;
signal \N__45549\ : std_logic;
signal \N__45546\ : std_logic;
signal \N__45543\ : std_logic;
signal \N__45538\ : std_logic;
signal \N__45535\ : std_logic;
signal \N__45534\ : std_logic;
signal \N__45531\ : std_logic;
signal \N__45528\ : std_logic;
signal \N__45525\ : std_logic;
signal \N__45522\ : std_logic;
signal \N__45519\ : std_logic;
signal \N__45516\ : std_logic;
signal \N__45511\ : std_logic;
signal \N__45510\ : std_logic;
signal \N__45507\ : std_logic;
signal \N__45504\ : std_logic;
signal \N__45501\ : std_logic;
signal \N__45498\ : std_logic;
signal \N__45497\ : std_logic;
signal \N__45494\ : std_logic;
signal \N__45491\ : std_logic;
signal \N__45488\ : std_logic;
signal \N__45483\ : std_logic;
signal \N__45478\ : std_logic;
signal \N__45477\ : std_logic;
signal \N__45474\ : std_logic;
signal \N__45471\ : std_logic;
signal \N__45470\ : std_logic;
signal \N__45467\ : std_logic;
signal \N__45464\ : std_logic;
signal \N__45461\ : std_logic;
signal \N__45456\ : std_logic;
signal \N__45451\ : std_logic;
signal \N__45448\ : std_logic;
signal \N__45445\ : std_logic;
signal \N__45442\ : std_logic;
signal \N__45439\ : std_logic;
signal \N__45436\ : std_logic;
signal \N__45433\ : std_logic;
signal \N__45432\ : std_logic;
signal \N__45431\ : std_logic;
signal \N__45428\ : std_logic;
signal \N__45425\ : std_logic;
signal \N__45422\ : std_logic;
signal \N__45419\ : std_logic;
signal \N__45414\ : std_logic;
signal \N__45411\ : std_logic;
signal \N__45408\ : std_logic;
signal \N__45403\ : std_logic;
signal \N__45400\ : std_logic;
signal \N__45397\ : std_logic;
signal \N__45394\ : std_logic;
signal \N__45391\ : std_logic;
signal \N__45388\ : std_logic;
signal \N__45385\ : std_logic;
signal \N__45382\ : std_logic;
signal \N__45381\ : std_logic;
signal \N__45380\ : std_logic;
signal \N__45377\ : std_logic;
signal \N__45376\ : std_logic;
signal \N__45373\ : std_logic;
signal \N__45370\ : std_logic;
signal \N__45367\ : std_logic;
signal \N__45364\ : std_logic;
signal \N__45361\ : std_logic;
signal \N__45356\ : std_logic;
signal \N__45353\ : std_logic;
signal \N__45350\ : std_logic;
signal \N__45347\ : std_logic;
signal \N__45344\ : std_logic;
signal \N__45341\ : std_logic;
signal \N__45338\ : std_logic;
signal \N__45331\ : std_logic;
signal \N__45330\ : std_logic;
signal \N__45329\ : std_logic;
signal \N__45328\ : std_logic;
signal \N__45327\ : std_logic;
signal \N__45324\ : std_logic;
signal \N__45317\ : std_logic;
signal \N__45314\ : std_logic;
signal \N__45311\ : std_logic;
signal \N__45310\ : std_logic;
signal \N__45307\ : std_logic;
signal \N__45304\ : std_logic;
signal \N__45301\ : std_logic;
signal \N__45298\ : std_logic;
signal \N__45293\ : std_logic;
signal \N__45292\ : std_logic;
signal \N__45289\ : std_logic;
signal \N__45286\ : std_logic;
signal \N__45283\ : std_logic;
signal \N__45280\ : std_logic;
signal \N__45279\ : std_logic;
signal \N__45276\ : std_logic;
signal \N__45273\ : std_logic;
signal \N__45268\ : std_logic;
signal \N__45265\ : std_logic;
signal \N__45256\ : std_logic;
signal \N__45255\ : std_logic;
signal \N__45254\ : std_logic;
signal \N__45251\ : std_logic;
signal \N__45248\ : std_logic;
signal \N__45245\ : std_logic;
signal \N__45242\ : std_logic;
signal \N__45235\ : std_logic;
signal \N__45232\ : std_logic;
signal \N__45231\ : std_logic;
signal \N__45228\ : std_logic;
signal \N__45227\ : std_logic;
signal \N__45224\ : std_logic;
signal \N__45221\ : std_logic;
signal \N__45218\ : std_logic;
signal \N__45211\ : std_logic;
signal \N__45208\ : std_logic;
signal \N__45205\ : std_logic;
signal \N__45202\ : std_logic;
signal \N__45201\ : std_logic;
signal \N__45198\ : std_logic;
signal \N__45195\ : std_logic;
signal \N__45192\ : std_logic;
signal \N__45189\ : std_logic;
signal \N__45186\ : std_logic;
signal \N__45183\ : std_logic;
signal \N__45180\ : std_logic;
signal \N__45179\ : std_logic;
signal \N__45176\ : std_logic;
signal \N__45173\ : std_logic;
signal \N__45170\ : std_logic;
signal \N__45163\ : std_logic;
signal \N__45160\ : std_logic;
signal \N__45159\ : std_logic;
signal \N__45156\ : std_logic;
signal \N__45155\ : std_logic;
signal \N__45152\ : std_logic;
signal \N__45149\ : std_logic;
signal \N__45144\ : std_logic;
signal \N__45139\ : std_logic;
signal \N__45138\ : std_logic;
signal \N__45135\ : std_logic;
signal \N__45132\ : std_logic;
signal \N__45129\ : std_logic;
signal \N__45126\ : std_logic;
signal \N__45123\ : std_logic;
signal \N__45120\ : std_logic;
signal \N__45117\ : std_logic;
signal \N__45114\ : std_logic;
signal \N__45113\ : std_logic;
signal \N__45110\ : std_logic;
signal \N__45107\ : std_logic;
signal \N__45104\ : std_logic;
signal \N__45101\ : std_logic;
signal \N__45098\ : std_logic;
signal \N__45091\ : std_logic;
signal \N__45088\ : std_logic;
signal \N__45087\ : std_logic;
signal \N__45086\ : std_logic;
signal \N__45083\ : std_logic;
signal \N__45080\ : std_logic;
signal \N__45077\ : std_logic;
signal \N__45074\ : std_logic;
signal \N__45067\ : std_logic;
signal \N__45064\ : std_logic;
signal \N__45061\ : std_logic;
signal \N__45058\ : std_logic;
signal \N__45055\ : std_logic;
signal \N__45052\ : std_logic;
signal \N__45049\ : std_logic;
signal \N__45046\ : std_logic;
signal \N__45043\ : std_logic;
signal \N__45040\ : std_logic;
signal \N__45039\ : std_logic;
signal \N__45034\ : std_logic;
signal \N__45031\ : std_logic;
signal \N__45028\ : std_logic;
signal \N__45025\ : std_logic;
signal \N__45022\ : std_logic;
signal \N__45019\ : std_logic;
signal \N__45016\ : std_logic;
signal \N__45013\ : std_logic;
signal \N__45010\ : std_logic;
signal \N__45007\ : std_logic;
signal \N__45004\ : std_logic;
signal \N__45001\ : std_logic;
signal \N__44998\ : std_logic;
signal \N__44995\ : std_logic;
signal \N__44992\ : std_logic;
signal \N__44989\ : std_logic;
signal \N__44988\ : std_logic;
signal \N__44985\ : std_logic;
signal \N__44982\ : std_logic;
signal \N__44979\ : std_logic;
signal \N__44974\ : std_logic;
signal \N__44971\ : std_logic;
signal \N__44968\ : std_logic;
signal \N__44967\ : std_logic;
signal \N__44964\ : std_logic;
signal \N__44961\ : std_logic;
signal \N__44956\ : std_logic;
signal \N__44953\ : std_logic;
signal \N__44952\ : std_logic;
signal \N__44949\ : std_logic;
signal \N__44946\ : std_logic;
signal \N__44943\ : std_logic;
signal \N__44938\ : std_logic;
signal \N__44935\ : std_logic;
signal \N__44932\ : std_logic;
signal \N__44931\ : std_logic;
signal \N__44928\ : std_logic;
signal \N__44925\ : std_logic;
signal \N__44920\ : std_logic;
signal \N__44917\ : std_logic;
signal \N__44914\ : std_logic;
signal \N__44911\ : std_logic;
signal \N__44910\ : std_logic;
signal \N__44907\ : std_logic;
signal \N__44906\ : std_logic;
signal \N__44903\ : std_logic;
signal \N__44902\ : std_logic;
signal \N__44899\ : std_logic;
signal \N__44896\ : std_logic;
signal \N__44893\ : std_logic;
signal \N__44890\ : std_logic;
signal \N__44887\ : std_logic;
signal \N__44884\ : std_logic;
signal \N__44879\ : std_logic;
signal \N__44872\ : std_logic;
signal \N__44871\ : std_logic;
signal \N__44868\ : std_logic;
signal \N__44865\ : std_logic;
signal \N__44862\ : std_logic;
signal \N__44857\ : std_logic;
signal \N__44854\ : std_logic;
signal \N__44851\ : std_logic;
signal \N__44850\ : std_logic;
signal \N__44849\ : std_logic;
signal \N__44848\ : std_logic;
signal \N__44847\ : std_logic;
signal \N__44846\ : std_logic;
signal \N__44843\ : std_logic;
signal \N__44840\ : std_logic;
signal \N__44837\ : std_logic;
signal \N__44834\ : std_logic;
signal \N__44831\ : std_logic;
signal \N__44828\ : std_logic;
signal \N__44825\ : std_logic;
signal \N__44822\ : std_logic;
signal \N__44819\ : std_logic;
signal \N__44812\ : std_logic;
signal \N__44809\ : std_logic;
signal \N__44806\ : std_logic;
signal \N__44801\ : std_logic;
signal \N__44800\ : std_logic;
signal \N__44799\ : std_logic;
signal \N__44796\ : std_logic;
signal \N__44793\ : std_logic;
signal \N__44790\ : std_logic;
signal \N__44785\ : std_logic;
signal \N__44782\ : std_logic;
signal \N__44779\ : std_logic;
signal \N__44776\ : std_logic;
signal \N__44767\ : std_logic;
signal \N__44764\ : std_logic;
signal \N__44761\ : std_logic;
signal \N__44758\ : std_logic;
signal \N__44755\ : std_logic;
signal \N__44754\ : std_logic;
signal \N__44751\ : std_logic;
signal \N__44748\ : std_logic;
signal \N__44745\ : std_logic;
signal \N__44744\ : std_logic;
signal \N__44741\ : std_logic;
signal \N__44738\ : std_logic;
signal \N__44735\ : std_logic;
signal \N__44732\ : std_logic;
signal \N__44725\ : std_logic;
signal \N__44722\ : std_logic;
signal \N__44719\ : std_logic;
signal \N__44718\ : std_logic;
signal \N__44717\ : std_logic;
signal \N__44714\ : std_logic;
signal \N__44709\ : std_logic;
signal \N__44704\ : std_logic;
signal \N__44703\ : std_logic;
signal \N__44700\ : std_logic;
signal \N__44697\ : std_logic;
signal \N__44692\ : std_logic;
signal \N__44689\ : std_logic;
signal \N__44688\ : std_logic;
signal \N__44685\ : std_logic;
signal \N__44682\ : std_logic;
signal \N__44679\ : std_logic;
signal \N__44674\ : std_logic;
signal \N__44671\ : std_logic;
signal \N__44670\ : std_logic;
signal \N__44667\ : std_logic;
signal \N__44664\ : std_logic;
signal \N__44661\ : std_logic;
signal \N__44656\ : std_logic;
signal \N__44653\ : std_logic;
signal \N__44650\ : std_logic;
signal \N__44649\ : std_logic;
signal \N__44646\ : std_logic;
signal \N__44643\ : std_logic;
signal \N__44640\ : std_logic;
signal \N__44635\ : std_logic;
signal \N__44632\ : std_logic;
signal \N__44631\ : std_logic;
signal \N__44628\ : std_logic;
signal \N__44625\ : std_logic;
signal \N__44620\ : std_logic;
signal \N__44617\ : std_logic;
signal \N__44616\ : std_logic;
signal \N__44613\ : std_logic;
signal \N__44610\ : std_logic;
signal \N__44605\ : std_logic;
signal \N__44602\ : std_logic;
signal \N__44601\ : std_logic;
signal \N__44598\ : std_logic;
signal \N__44595\ : std_logic;
signal \N__44590\ : std_logic;
signal \N__44587\ : std_logic;
signal \N__44586\ : std_logic;
signal \N__44583\ : std_logic;
signal \N__44580\ : std_logic;
signal \N__44575\ : std_logic;
signal \N__44572\ : std_logic;
signal \N__44571\ : std_logic;
signal \N__44568\ : std_logic;
signal \N__44565\ : std_logic;
signal \N__44562\ : std_logic;
signal \N__44557\ : std_logic;
signal \N__44554\ : std_logic;
signal \N__44553\ : std_logic;
signal \N__44550\ : std_logic;
signal \N__44547\ : std_logic;
signal \N__44542\ : std_logic;
signal \N__44539\ : std_logic;
signal \N__44536\ : std_logic;
signal \N__44535\ : std_logic;
signal \N__44532\ : std_logic;
signal \N__44529\ : std_logic;
signal \N__44524\ : std_logic;
signal \N__44521\ : std_logic;
signal \N__44520\ : std_logic;
signal \N__44517\ : std_logic;
signal \N__44514\ : std_logic;
signal \N__44509\ : std_logic;
signal \N__44506\ : std_logic;
signal \N__44505\ : std_logic;
signal \N__44502\ : std_logic;
signal \N__44499\ : std_logic;
signal \N__44496\ : std_logic;
signal \N__44491\ : std_logic;
signal \N__44488\ : std_logic;
signal \N__44487\ : std_logic;
signal \N__44484\ : std_logic;
signal \N__44481\ : std_logic;
signal \N__44476\ : std_logic;
signal \N__44473\ : std_logic;
signal \N__44472\ : std_logic;
signal \N__44469\ : std_logic;
signal \N__44466\ : std_logic;
signal \N__44463\ : std_logic;
signal \N__44458\ : std_logic;
signal \N__44455\ : std_logic;
signal \N__44454\ : std_logic;
signal \N__44451\ : std_logic;
signal \N__44448\ : std_logic;
signal \N__44443\ : std_logic;
signal \N__44440\ : std_logic;
signal \N__44437\ : std_logic;
signal \N__44434\ : std_logic;
signal \N__44431\ : std_logic;
signal \N__44428\ : std_logic;
signal \N__44425\ : std_logic;
signal \N__44422\ : std_logic;
signal \N__44419\ : std_logic;
signal \N__44418\ : std_logic;
signal \N__44415\ : std_logic;
signal \N__44412\ : std_logic;
signal \N__44411\ : std_logic;
signal \N__44408\ : std_logic;
signal \N__44405\ : std_logic;
signal \N__44402\ : std_logic;
signal \N__44401\ : std_logic;
signal \N__44400\ : std_logic;
signal \N__44397\ : std_logic;
signal \N__44392\ : std_logic;
signal \N__44389\ : std_logic;
signal \N__44386\ : std_logic;
signal \N__44379\ : std_logic;
signal \N__44374\ : std_logic;
signal \N__44371\ : std_logic;
signal \N__44368\ : std_logic;
signal \N__44365\ : std_logic;
signal \N__44362\ : std_logic;
signal \N__44359\ : std_logic;
signal \N__44356\ : std_logic;
signal \N__44353\ : std_logic;
signal \N__44350\ : std_logic;
signal \N__44347\ : std_logic;
signal \N__44344\ : std_logic;
signal \N__44341\ : std_logic;
signal \N__44338\ : std_logic;
signal \N__44335\ : std_logic;
signal \N__44332\ : std_logic;
signal \N__44329\ : std_logic;
signal \N__44326\ : std_logic;
signal \N__44323\ : std_logic;
signal \N__44322\ : std_logic;
signal \N__44319\ : std_logic;
signal \N__44316\ : std_logic;
signal \N__44311\ : std_logic;
signal \N__44310\ : std_logic;
signal \N__44307\ : std_logic;
signal \N__44304\ : std_logic;
signal \N__44301\ : std_logic;
signal \N__44298\ : std_logic;
signal \N__44295\ : std_logic;
signal \N__44292\ : std_logic;
signal \N__44287\ : std_logic;
signal \N__44284\ : std_logic;
signal \N__44283\ : std_logic;
signal \N__44282\ : std_logic;
signal \N__44279\ : std_logic;
signal \N__44276\ : std_logic;
signal \N__44273\ : std_logic;
signal \N__44272\ : std_logic;
signal \N__44271\ : std_logic;
signal \N__44270\ : std_logic;
signal \N__44263\ : std_logic;
signal \N__44260\ : std_logic;
signal \N__44257\ : std_logic;
signal \N__44254\ : std_logic;
signal \N__44251\ : std_logic;
signal \N__44242\ : std_logic;
signal \N__44239\ : std_logic;
signal \N__44236\ : std_logic;
signal \N__44233\ : std_logic;
signal \N__44232\ : std_logic;
signal \N__44231\ : std_logic;
signal \N__44228\ : std_logic;
signal \N__44225\ : std_logic;
signal \N__44222\ : std_logic;
signal \N__44219\ : std_logic;
signal \N__44216\ : std_logic;
signal \N__44213\ : std_logic;
signal \N__44210\ : std_logic;
signal \N__44207\ : std_logic;
signal \N__44204\ : std_logic;
signal \N__44197\ : std_logic;
signal \N__44194\ : std_logic;
signal \N__44191\ : std_logic;
signal \N__44188\ : std_logic;
signal \N__44185\ : std_logic;
signal \N__44182\ : std_logic;
signal \N__44179\ : std_logic;
signal \N__44176\ : std_logic;
signal \N__44173\ : std_logic;
signal \N__44170\ : std_logic;
signal \N__44167\ : std_logic;
signal \N__44164\ : std_logic;
signal \N__44161\ : std_logic;
signal \N__44158\ : std_logic;
signal \N__44155\ : std_logic;
signal \N__44152\ : std_logic;
signal \N__44149\ : std_logic;
signal \N__44148\ : std_logic;
signal \N__44147\ : std_logic;
signal \N__44146\ : std_logic;
signal \N__44143\ : std_logic;
signal \N__44140\ : std_logic;
signal \N__44137\ : std_logic;
signal \N__44134\ : std_logic;
signal \N__44131\ : std_logic;
signal \N__44128\ : std_logic;
signal \N__44127\ : std_logic;
signal \N__44124\ : std_logic;
signal \N__44121\ : std_logic;
signal \N__44116\ : std_logic;
signal \N__44113\ : std_logic;
signal \N__44112\ : std_logic;
signal \N__44109\ : std_logic;
signal \N__44108\ : std_logic;
signal \N__44107\ : std_logic;
signal \N__44104\ : std_logic;
signal \N__44101\ : std_logic;
signal \N__44098\ : std_logic;
signal \N__44095\ : std_logic;
signal \N__44092\ : std_logic;
signal \N__44089\ : std_logic;
signal \N__44086\ : std_logic;
signal \N__44085\ : std_logic;
signal \N__44084\ : std_logic;
signal \N__44081\ : std_logic;
signal \N__44076\ : std_logic;
signal \N__44073\ : std_logic;
signal \N__44066\ : std_logic;
signal \N__44061\ : std_logic;
signal \N__44058\ : std_logic;
signal \N__44053\ : std_logic;
signal \N__44050\ : std_logic;
signal \N__44047\ : std_logic;
signal \N__44040\ : std_logic;
signal \N__44035\ : std_logic;
signal \N__44032\ : std_logic;
signal \N__44031\ : std_logic;
signal \N__44028\ : std_logic;
signal \N__44025\ : std_logic;
signal \N__44022\ : std_logic;
signal \N__44019\ : std_logic;
signal \N__44016\ : std_logic;
signal \N__44013\ : std_logic;
signal \N__44010\ : std_logic;
signal \N__44009\ : std_logic;
signal \N__44006\ : std_logic;
signal \N__44003\ : std_logic;
signal \N__44000\ : std_logic;
signal \N__43997\ : std_logic;
signal \N__43990\ : std_logic;
signal \N__43987\ : std_logic;
signal \N__43984\ : std_logic;
signal \N__43981\ : std_logic;
signal \N__43980\ : std_logic;
signal \N__43977\ : std_logic;
signal \N__43974\ : std_logic;
signal \N__43969\ : std_logic;
signal \N__43966\ : std_logic;
signal \N__43963\ : std_logic;
signal \N__43960\ : std_logic;
signal \N__43957\ : std_logic;
signal \N__43954\ : std_logic;
signal \N__43951\ : std_logic;
signal \N__43948\ : std_logic;
signal \N__43945\ : std_logic;
signal \N__43942\ : std_logic;
signal \N__43939\ : std_logic;
signal \N__43936\ : std_logic;
signal \N__43933\ : std_logic;
signal \N__43930\ : std_logic;
signal \N__43927\ : std_logic;
signal \N__43924\ : std_logic;
signal \N__43923\ : std_logic;
signal \N__43920\ : std_logic;
signal \N__43917\ : std_logic;
signal \N__43914\ : std_logic;
signal \N__43911\ : std_logic;
signal \N__43908\ : std_logic;
signal \N__43905\ : std_logic;
signal \N__43902\ : std_logic;
signal \N__43899\ : std_logic;
signal \N__43896\ : std_logic;
signal \N__43893\ : std_logic;
signal \N__43890\ : std_logic;
signal \N__43887\ : std_logic;
signal \N__43884\ : std_logic;
signal \N__43881\ : std_logic;
signal \N__43878\ : std_logic;
signal \N__43873\ : std_logic;
signal \N__43872\ : std_logic;
signal \N__43871\ : std_logic;
signal \N__43866\ : std_logic;
signal \N__43865\ : std_logic;
signal \N__43864\ : std_logic;
signal \N__43861\ : std_logic;
signal \N__43858\ : std_logic;
signal \N__43855\ : std_logic;
signal \N__43852\ : std_logic;
signal \N__43849\ : std_logic;
signal \N__43848\ : std_logic;
signal \N__43847\ : std_logic;
signal \N__43842\ : std_logic;
signal \N__43837\ : std_logic;
signal \N__43834\ : std_logic;
signal \N__43831\ : std_logic;
signal \N__43822\ : std_logic;
signal \N__43821\ : std_logic;
signal \N__43818\ : std_logic;
signal \N__43817\ : std_logic;
signal \N__43816\ : std_logic;
signal \N__43813\ : std_logic;
signal \N__43810\ : std_logic;
signal \N__43807\ : std_logic;
signal \N__43806\ : std_logic;
signal \N__43803\ : std_logic;
signal \N__43802\ : std_logic;
signal \N__43797\ : std_logic;
signal \N__43796\ : std_logic;
signal \N__43793\ : std_logic;
signal \N__43790\ : std_logic;
signal \N__43787\ : std_logic;
signal \N__43784\ : std_logic;
signal \N__43781\ : std_logic;
signal \N__43778\ : std_logic;
signal \N__43775\ : std_logic;
signal \N__43772\ : std_logic;
signal \N__43769\ : std_logic;
signal \N__43768\ : std_logic;
signal \N__43761\ : std_logic;
signal \N__43760\ : std_logic;
signal \N__43755\ : std_logic;
signal \N__43752\ : std_logic;
signal \N__43749\ : std_logic;
signal \N__43746\ : std_logic;
signal \N__43743\ : std_logic;
signal \N__43740\ : std_logic;
signal \N__43735\ : std_logic;
signal \N__43732\ : std_logic;
signal \N__43729\ : std_logic;
signal \N__43726\ : std_logic;
signal \N__43723\ : std_logic;
signal \N__43720\ : std_logic;
signal \N__43711\ : std_logic;
signal \N__43710\ : std_logic;
signal \N__43707\ : std_logic;
signal \N__43704\ : std_logic;
signal \N__43701\ : std_logic;
signal \N__43698\ : std_logic;
signal \N__43695\ : std_logic;
signal \N__43692\ : std_logic;
signal \N__43687\ : std_logic;
signal \N__43686\ : std_logic;
signal \N__43685\ : std_logic;
signal \N__43678\ : std_logic;
signal \N__43677\ : std_logic;
signal \N__43674\ : std_logic;
signal \N__43673\ : std_logic;
signal \N__43670\ : std_logic;
signal \N__43667\ : std_logic;
signal \N__43664\ : std_logic;
signal \N__43661\ : std_logic;
signal \N__43658\ : std_logic;
signal \N__43655\ : std_logic;
signal \N__43652\ : std_logic;
signal \N__43645\ : std_logic;
signal \N__43642\ : std_logic;
signal \N__43641\ : std_logic;
signal \N__43638\ : std_logic;
signal \N__43635\ : std_logic;
signal \N__43630\ : std_logic;
signal \N__43627\ : std_logic;
signal \N__43624\ : std_logic;
signal \N__43621\ : std_logic;
signal \N__43618\ : std_logic;
signal \N__43615\ : std_logic;
signal \N__43612\ : std_logic;
signal \N__43609\ : std_logic;
signal \N__43606\ : std_logic;
signal \N__43603\ : std_logic;
signal \N__43600\ : std_logic;
signal \N__43597\ : std_logic;
signal \N__43594\ : std_logic;
signal \N__43591\ : std_logic;
signal \N__43588\ : std_logic;
signal \N__43585\ : std_logic;
signal \N__43582\ : std_logic;
signal \N__43579\ : std_logic;
signal \N__43576\ : std_logic;
signal \N__43573\ : std_logic;
signal \N__43570\ : std_logic;
signal \N__43569\ : std_logic;
signal \N__43566\ : std_logic;
signal \N__43563\ : std_logic;
signal \N__43562\ : std_logic;
signal \N__43559\ : std_logic;
signal \N__43556\ : std_logic;
signal \N__43553\ : std_logic;
signal \N__43546\ : std_logic;
signal \N__43545\ : std_logic;
signal \N__43542\ : std_logic;
signal \N__43539\ : std_logic;
signal \N__43534\ : std_logic;
signal \N__43533\ : std_logic;
signal \N__43532\ : std_logic;
signal \N__43529\ : std_logic;
signal \N__43526\ : std_logic;
signal \N__43525\ : std_logic;
signal \N__43524\ : std_logic;
signal \N__43521\ : std_logic;
signal \N__43520\ : std_logic;
signal \N__43517\ : std_logic;
signal \N__43514\ : std_logic;
signal \N__43511\ : std_logic;
signal \N__43508\ : std_logic;
signal \N__43505\ : std_logic;
signal \N__43504\ : std_logic;
signal \N__43501\ : std_logic;
signal \N__43496\ : std_logic;
signal \N__43493\ : std_logic;
signal \N__43488\ : std_logic;
signal \N__43487\ : std_logic;
signal \N__43484\ : std_logic;
signal \N__43481\ : std_logic;
signal \N__43478\ : std_logic;
signal \N__43475\ : std_logic;
signal \N__43474\ : std_logic;
signal \N__43471\ : std_logic;
signal \N__43468\ : std_logic;
signal \N__43465\ : std_logic;
signal \N__43462\ : std_logic;
signal \N__43461\ : std_logic;
signal \N__43456\ : std_logic;
signal \N__43453\ : std_logic;
signal \N__43450\ : std_logic;
signal \N__43447\ : std_logic;
signal \N__43444\ : std_logic;
signal \N__43441\ : std_logic;
signal \N__43438\ : std_logic;
signal \N__43435\ : std_logic;
signal \N__43428\ : std_logic;
signal \N__43417\ : std_logic;
signal \N__43414\ : std_logic;
signal \N__43413\ : std_logic;
signal \N__43410\ : std_logic;
signal \N__43409\ : std_logic;
signal \N__43406\ : std_logic;
signal \N__43403\ : std_logic;
signal \N__43400\ : std_logic;
signal \N__43397\ : std_logic;
signal \N__43390\ : std_logic;
signal \N__43387\ : std_logic;
signal \N__43384\ : std_logic;
signal \N__43383\ : std_logic;
signal \N__43382\ : std_logic;
signal \N__43379\ : std_logic;
signal \N__43376\ : std_logic;
signal \N__43375\ : std_logic;
signal \N__43374\ : std_logic;
signal \N__43371\ : std_logic;
signal \N__43366\ : std_logic;
signal \N__43363\ : std_logic;
signal \N__43360\ : std_logic;
signal \N__43357\ : std_logic;
signal \N__43354\ : std_logic;
signal \N__43351\ : std_logic;
signal \N__43348\ : std_logic;
signal \N__43347\ : std_logic;
signal \N__43344\ : std_logic;
signal \N__43339\ : std_logic;
signal \N__43336\ : std_logic;
signal \N__43333\ : std_logic;
signal \N__43328\ : std_logic;
signal \N__43321\ : std_logic;
signal \N__43320\ : std_logic;
signal \N__43319\ : std_logic;
signal \N__43316\ : std_logic;
signal \N__43313\ : std_logic;
signal \N__43310\ : std_logic;
signal \N__43305\ : std_logic;
signal \N__43300\ : std_logic;
signal \N__43299\ : std_logic;
signal \N__43296\ : std_logic;
signal \N__43295\ : std_logic;
signal \N__43292\ : std_logic;
signal \N__43291\ : std_logic;
signal \N__43288\ : std_logic;
signal \N__43285\ : std_logic;
signal \N__43284\ : std_logic;
signal \N__43281\ : std_logic;
signal \N__43278\ : std_logic;
signal \N__43277\ : std_logic;
signal \N__43276\ : std_logic;
signal \N__43275\ : std_logic;
signal \N__43274\ : std_logic;
signal \N__43273\ : std_logic;
signal \N__43268\ : std_logic;
signal \N__43265\ : std_logic;
signal \N__43260\ : std_logic;
signal \N__43257\ : std_logic;
signal \N__43254\ : std_logic;
signal \N__43249\ : std_logic;
signal \N__43246\ : std_logic;
signal \N__43243\ : std_logic;
signal \N__43228\ : std_logic;
signal \N__43225\ : std_logic;
signal \N__43222\ : std_logic;
signal \N__43219\ : std_logic;
signal \N__43218\ : std_logic;
signal \N__43213\ : std_logic;
signal \N__43210\ : std_logic;
signal \N__43207\ : std_logic;
signal \N__43204\ : std_logic;
signal \N__43201\ : std_logic;
signal \N__43198\ : std_logic;
signal \N__43195\ : std_logic;
signal \N__43192\ : std_logic;
signal \N__43189\ : std_logic;
signal \N__43186\ : std_logic;
signal \N__43183\ : std_logic;
signal \N__43180\ : std_logic;
signal \N__43177\ : std_logic;
signal \N__43174\ : std_logic;
signal \N__43171\ : std_logic;
signal \N__43168\ : std_logic;
signal \N__43165\ : std_logic;
signal \N__43162\ : std_logic;
signal \N__43159\ : std_logic;
signal \N__43158\ : std_logic;
signal \N__43155\ : std_logic;
signal \N__43152\ : std_logic;
signal \N__43149\ : std_logic;
signal \N__43146\ : std_logic;
signal \N__43143\ : std_logic;
signal \N__43140\ : std_logic;
signal \N__43137\ : std_logic;
signal \N__43134\ : std_logic;
signal \N__43131\ : std_logic;
signal \N__43128\ : std_logic;
signal \N__43125\ : std_logic;
signal \N__43122\ : std_logic;
signal \N__43119\ : std_logic;
signal \N__43116\ : std_logic;
signal \N__43113\ : std_logic;
signal \N__43108\ : std_logic;
signal \N__43105\ : std_logic;
signal \N__43104\ : std_logic;
signal \N__43101\ : std_logic;
signal \N__43098\ : std_logic;
signal \N__43097\ : std_logic;
signal \N__43094\ : std_logic;
signal \N__43091\ : std_logic;
signal \N__43088\ : std_logic;
signal \N__43085\ : std_logic;
signal \N__43082\ : std_logic;
signal \N__43079\ : std_logic;
signal \N__43076\ : std_logic;
signal \N__43073\ : std_logic;
signal \N__43066\ : std_logic;
signal \N__43065\ : std_logic;
signal \N__43062\ : std_logic;
signal \N__43059\ : std_logic;
signal \N__43056\ : std_logic;
signal \N__43055\ : std_logic;
signal \N__43050\ : std_logic;
signal \N__43047\ : std_logic;
signal \N__43044\ : std_logic;
signal \N__43039\ : std_logic;
signal \N__43038\ : std_logic;
signal \N__43035\ : std_logic;
signal \N__43032\ : std_logic;
signal \N__43029\ : std_logic;
signal \N__43024\ : std_logic;
signal \N__43023\ : std_logic;
signal \N__43020\ : std_logic;
signal \N__43017\ : std_logic;
signal \N__43014\ : std_logic;
signal \N__43009\ : std_logic;
signal \N__43006\ : std_logic;
signal \N__43003\ : std_logic;
signal \N__43000\ : std_logic;
signal \N__42997\ : std_logic;
signal \N__42994\ : std_logic;
signal \N__42991\ : std_logic;
signal \N__42988\ : std_logic;
signal \N__42985\ : std_logic;
signal \N__42982\ : std_logic;
signal \N__42979\ : std_logic;
signal \N__42976\ : std_logic;
signal \N__42973\ : std_logic;
signal \N__42970\ : std_logic;
signal \N__42967\ : std_logic;
signal \N__42966\ : std_logic;
signal \N__42963\ : std_logic;
signal \N__42960\ : std_logic;
signal \N__42957\ : std_logic;
signal \N__42954\ : std_logic;
signal \N__42951\ : std_logic;
signal \N__42948\ : std_logic;
signal \N__42945\ : std_logic;
signal \N__42942\ : std_logic;
signal \N__42939\ : std_logic;
signal \N__42936\ : std_logic;
signal \N__42933\ : std_logic;
signal \N__42930\ : std_logic;
signal \N__42927\ : std_logic;
signal \N__42924\ : std_logic;
signal \N__42921\ : std_logic;
signal \N__42916\ : std_logic;
signal \N__42915\ : std_logic;
signal \N__42912\ : std_logic;
signal \N__42909\ : std_logic;
signal \N__42906\ : std_logic;
signal \N__42901\ : std_logic;
signal \N__42898\ : std_logic;
signal \N__42895\ : std_logic;
signal \N__42892\ : std_logic;
signal \N__42889\ : std_logic;
signal \N__42886\ : std_logic;
signal \N__42885\ : std_logic;
signal \N__42882\ : std_logic;
signal \N__42879\ : std_logic;
signal \N__42874\ : std_logic;
signal \N__42873\ : std_logic;
signal \N__42870\ : std_logic;
signal \N__42867\ : std_logic;
signal \N__42864\ : std_logic;
signal \N__42859\ : std_logic;
signal \N__42856\ : std_logic;
signal \N__42855\ : std_logic;
signal \N__42852\ : std_logic;
signal \N__42849\ : std_logic;
signal \N__42846\ : std_logic;
signal \N__42841\ : std_logic;
signal \N__42840\ : std_logic;
signal \N__42839\ : std_logic;
signal \N__42836\ : std_logic;
signal \N__42833\ : std_logic;
signal \N__42830\ : std_logic;
signal \N__42823\ : std_logic;
signal \N__42822\ : std_logic;
signal \N__42819\ : std_logic;
signal \N__42816\ : std_logic;
signal \N__42815\ : std_logic;
signal \N__42812\ : std_logic;
signal \N__42809\ : std_logic;
signal \N__42808\ : std_logic;
signal \N__42805\ : std_logic;
signal \N__42804\ : std_logic;
signal \N__42801\ : std_logic;
signal \N__42798\ : std_logic;
signal \N__42795\ : std_logic;
signal \N__42792\ : std_logic;
signal \N__42789\ : std_logic;
signal \N__42788\ : std_logic;
signal \N__42785\ : std_logic;
signal \N__42782\ : std_logic;
signal \N__42779\ : std_logic;
signal \N__42774\ : std_logic;
signal \N__42771\ : std_logic;
signal \N__42768\ : std_logic;
signal \N__42759\ : std_logic;
signal \N__42754\ : std_logic;
signal \N__42753\ : std_logic;
signal \N__42750\ : std_logic;
signal \N__42747\ : std_logic;
signal \N__42746\ : std_logic;
signal \N__42743\ : std_logic;
signal \N__42740\ : std_logic;
signal \N__42737\ : std_logic;
signal \N__42732\ : std_logic;
signal \N__42727\ : std_logic;
signal \N__42726\ : std_logic;
signal \N__42725\ : std_logic;
signal \N__42720\ : std_logic;
signal \N__42717\ : std_logic;
signal \N__42712\ : std_logic;
signal \N__42711\ : std_logic;
signal \N__42708\ : std_logic;
signal \N__42705\ : std_logic;
signal \N__42702\ : std_logic;
signal \N__42701\ : std_logic;
signal \N__42698\ : std_logic;
signal \N__42695\ : std_logic;
signal \N__42692\ : std_logic;
signal \N__42689\ : std_logic;
signal \N__42682\ : std_logic;
signal \N__42679\ : std_logic;
signal \N__42678\ : std_logic;
signal \N__42677\ : std_logic;
signal \N__42674\ : std_logic;
signal \N__42671\ : std_logic;
signal \N__42668\ : std_logic;
signal \N__42663\ : std_logic;
signal \N__42658\ : std_logic;
signal \N__42655\ : std_logic;
signal \N__42654\ : std_logic;
signal \N__42651\ : std_logic;
signal \N__42648\ : std_logic;
signal \N__42645\ : std_logic;
signal \N__42644\ : std_logic;
signal \N__42641\ : std_logic;
signal \N__42638\ : std_logic;
signal \N__42635\ : std_logic;
signal \N__42632\ : std_logic;
signal \N__42625\ : std_logic;
signal \N__42624\ : std_logic;
signal \N__42623\ : std_logic;
signal \N__42620\ : std_logic;
signal \N__42619\ : std_logic;
signal \N__42616\ : std_logic;
signal \N__42615\ : std_logic;
signal \N__42612\ : std_logic;
signal \N__42609\ : std_logic;
signal \N__42606\ : std_logic;
signal \N__42603\ : std_logic;
signal \N__42600\ : std_logic;
signal \N__42597\ : std_logic;
signal \N__42596\ : std_logic;
signal \N__42593\ : std_logic;
signal \N__42590\ : std_logic;
signal \N__42587\ : std_logic;
signal \N__42584\ : std_logic;
signal \N__42581\ : std_logic;
signal \N__42578\ : std_logic;
signal \N__42575\ : std_logic;
signal \N__42570\ : std_logic;
signal \N__42567\ : std_logic;
signal \N__42562\ : std_logic;
signal \N__42559\ : std_logic;
signal \N__42556\ : std_logic;
signal \N__42551\ : std_logic;
signal \N__42544\ : std_logic;
signal \N__42543\ : std_logic;
signal \N__42540\ : std_logic;
signal \N__42537\ : std_logic;
signal \N__42534\ : std_logic;
signal \N__42531\ : std_logic;
signal \N__42530\ : std_logic;
signal \N__42527\ : std_logic;
signal \N__42524\ : std_logic;
signal \N__42521\ : std_logic;
signal \N__42518\ : std_logic;
signal \N__42515\ : std_logic;
signal \N__42508\ : std_logic;
signal \N__42507\ : std_logic;
signal \N__42506\ : std_logic;
signal \N__42503\ : std_logic;
signal \N__42500\ : std_logic;
signal \N__42497\ : std_logic;
signal \N__42490\ : std_logic;
signal \N__42489\ : std_logic;
signal \N__42484\ : std_logic;
signal \N__42481\ : std_logic;
signal \N__42478\ : std_logic;
signal \N__42475\ : std_logic;
signal \N__42472\ : std_logic;
signal \N__42471\ : std_logic;
signal \N__42468\ : std_logic;
signal \N__42465\ : std_logic;
signal \N__42460\ : std_logic;
signal \N__42459\ : std_logic;
signal \N__42456\ : std_logic;
signal \N__42453\ : std_logic;
signal \N__42450\ : std_logic;
signal \N__42447\ : std_logic;
signal \N__42444\ : std_logic;
signal \N__42439\ : std_logic;
signal \N__42436\ : std_logic;
signal \N__42435\ : std_logic;
signal \N__42432\ : std_logic;
signal \N__42429\ : std_logic;
signal \N__42426\ : std_logic;
signal \N__42423\ : std_logic;
signal \N__42420\ : std_logic;
signal \N__42417\ : std_logic;
signal \N__42412\ : std_logic;
signal \N__42409\ : std_logic;
signal \N__42408\ : std_logic;
signal \N__42405\ : std_logic;
signal \N__42402\ : std_logic;
signal \N__42397\ : std_logic;
signal \N__42396\ : std_logic;
signal \N__42393\ : std_logic;
signal \N__42390\ : std_logic;
signal \N__42387\ : std_logic;
signal \N__42382\ : std_logic;
signal \N__42381\ : std_logic;
signal \N__42376\ : std_logic;
signal \N__42373\ : std_logic;
signal \N__42370\ : std_logic;
signal \N__42367\ : std_logic;
signal \N__42364\ : std_logic;
signal \N__42361\ : std_logic;
signal \N__42358\ : std_logic;
signal \N__42357\ : std_logic;
signal \N__42354\ : std_logic;
signal \N__42353\ : std_logic;
signal \N__42350\ : std_logic;
signal \N__42347\ : std_logic;
signal \N__42346\ : std_logic;
signal \N__42345\ : std_logic;
signal \N__42344\ : std_logic;
signal \N__42343\ : std_logic;
signal \N__42342\ : std_logic;
signal \N__42341\ : std_logic;
signal \N__42340\ : std_logic;
signal \N__42339\ : std_logic;
signal \N__42336\ : std_logic;
signal \N__42333\ : std_logic;
signal \N__42330\ : std_logic;
signal \N__42327\ : std_logic;
signal \N__42324\ : std_logic;
signal \N__42321\ : std_logic;
signal \N__42318\ : std_logic;
signal \N__42315\ : std_logic;
signal \N__42312\ : std_logic;
signal \N__42309\ : std_logic;
signal \N__42306\ : std_logic;
signal \N__42303\ : std_logic;
signal \N__42300\ : std_logic;
signal \N__42297\ : std_logic;
signal \N__42288\ : std_logic;
signal \N__42279\ : std_logic;
signal \N__42268\ : std_logic;
signal \N__42265\ : std_logic;
signal \N__42262\ : std_logic;
signal \N__42259\ : std_logic;
signal \N__42256\ : std_logic;
signal \N__42253\ : std_logic;
signal \N__42250\ : std_logic;
signal \N__42247\ : std_logic;
signal \N__42244\ : std_logic;
signal \N__42241\ : std_logic;
signal \N__42238\ : std_logic;
signal \N__42235\ : std_logic;
signal \N__42232\ : std_logic;
signal \N__42229\ : std_logic;
signal \N__42226\ : std_logic;
signal \N__42223\ : std_logic;
signal \N__42220\ : std_logic;
signal \N__42217\ : std_logic;
signal \N__42216\ : std_logic;
signal \N__42213\ : std_logic;
signal \N__42210\ : std_logic;
signal \N__42207\ : std_logic;
signal \N__42204\ : std_logic;
signal \N__42201\ : std_logic;
signal \N__42198\ : std_logic;
signal \N__42195\ : std_logic;
signal \N__42192\ : std_logic;
signal \N__42189\ : std_logic;
signal \N__42186\ : std_logic;
signal \N__42183\ : std_logic;
signal \N__42180\ : std_logic;
signal \N__42177\ : std_logic;
signal \N__42172\ : std_logic;
signal \N__42169\ : std_logic;
signal \N__42166\ : std_logic;
signal \N__42163\ : std_logic;
signal \N__42160\ : std_logic;
signal \N__42157\ : std_logic;
signal \N__42154\ : std_logic;
signal \N__42151\ : std_logic;
signal \N__42148\ : std_logic;
signal \N__42145\ : std_logic;
signal \N__42144\ : std_logic;
signal \N__42143\ : std_logic;
signal \N__42140\ : std_logic;
signal \N__42139\ : std_logic;
signal \N__42136\ : std_logic;
signal \N__42135\ : std_logic;
signal \N__42132\ : std_logic;
signal \N__42127\ : std_logic;
signal \N__42126\ : std_logic;
signal \N__42123\ : std_logic;
signal \N__42120\ : std_logic;
signal \N__42119\ : std_logic;
signal \N__42116\ : std_logic;
signal \N__42113\ : std_logic;
signal \N__42110\ : std_logic;
signal \N__42105\ : std_logic;
signal \N__42102\ : std_logic;
signal \N__42095\ : std_logic;
signal \N__42090\ : std_logic;
signal \N__42087\ : std_logic;
signal \N__42084\ : std_logic;
signal \N__42081\ : std_logic;
signal \N__42076\ : std_logic;
signal \N__42075\ : std_logic;
signal \N__42074\ : std_logic;
signal \N__42071\ : std_logic;
signal \N__42068\ : std_logic;
signal \N__42065\ : std_logic;
signal \N__42062\ : std_logic;
signal \N__42057\ : std_logic;
signal \N__42054\ : std_logic;
signal \N__42051\ : std_logic;
signal \N__42046\ : std_logic;
signal \N__42045\ : std_logic;
signal \N__42044\ : std_logic;
signal \N__42041\ : std_logic;
signal \N__42038\ : std_logic;
signal \N__42035\ : std_logic;
signal \N__42030\ : std_logic;
signal \N__42025\ : std_logic;
signal \N__42024\ : std_logic;
signal \N__42021\ : std_logic;
signal \N__42020\ : std_logic;
signal \N__42019\ : std_logic;
signal \N__42016\ : std_logic;
signal \N__42009\ : std_logic;
signal \N__42008\ : std_logic;
signal \N__42007\ : std_logic;
signal \N__42006\ : std_logic;
signal \N__42005\ : std_logic;
signal \N__42004\ : std_logic;
signal \N__42001\ : std_logic;
signal \N__41998\ : std_logic;
signal \N__41993\ : std_logic;
signal \N__41992\ : std_logic;
signal \N__41991\ : std_logic;
signal \N__41990\ : std_logic;
signal \N__41989\ : std_logic;
signal \N__41988\ : std_logic;
signal \N__41987\ : std_logic;
signal \N__41980\ : std_logic;
signal \N__41973\ : std_logic;
signal \N__41968\ : std_logic;
signal \N__41959\ : std_logic;
signal \N__41950\ : std_logic;
signal \N__41947\ : std_logic;
signal \N__41944\ : std_logic;
signal \N__41943\ : std_logic;
signal \N__41940\ : std_logic;
signal \N__41937\ : std_logic;
signal \N__41932\ : std_logic;
signal \N__41929\ : std_logic;
signal \N__41926\ : std_logic;
signal \N__41923\ : std_logic;
signal \N__41920\ : std_logic;
signal \N__41917\ : std_logic;
signal \N__41914\ : std_logic;
signal \N__41913\ : std_logic;
signal \N__41912\ : std_logic;
signal \N__41909\ : std_logic;
signal \N__41904\ : std_logic;
signal \N__41899\ : std_logic;
signal \N__41896\ : std_logic;
signal \N__41895\ : std_logic;
signal \N__41892\ : std_logic;
signal \N__41891\ : std_logic;
signal \N__41888\ : std_logic;
signal \N__41885\ : std_logic;
signal \N__41882\ : std_logic;
signal \N__41875\ : std_logic;
signal \N__41872\ : std_logic;
signal \N__41869\ : std_logic;
signal \N__41866\ : std_logic;
signal \N__41863\ : std_logic;
signal \N__41862\ : std_logic;
signal \N__41861\ : std_logic;
signal \N__41858\ : std_logic;
signal \N__41855\ : std_logic;
signal \N__41852\ : std_logic;
signal \N__41847\ : std_logic;
signal \N__41842\ : std_logic;
signal \N__41841\ : std_logic;
signal \N__41836\ : std_logic;
signal \N__41833\ : std_logic;
signal \N__41830\ : std_logic;
signal \N__41827\ : std_logic;
signal \N__41826\ : std_logic;
signal \N__41825\ : std_logic;
signal \N__41822\ : std_logic;
signal \N__41819\ : std_logic;
signal \N__41816\ : std_logic;
signal \N__41813\ : std_logic;
signal \N__41808\ : std_logic;
signal \N__41805\ : std_logic;
signal \N__41802\ : std_logic;
signal \N__41797\ : std_logic;
signal \N__41796\ : std_logic;
signal \N__41791\ : std_logic;
signal \N__41788\ : std_logic;
signal \N__41785\ : std_logic;
signal \N__41782\ : std_logic;
signal \N__41781\ : std_logic;
signal \N__41778\ : std_logic;
signal \N__41775\ : std_logic;
signal \N__41772\ : std_logic;
signal \N__41769\ : std_logic;
signal \N__41766\ : std_logic;
signal \N__41763\ : std_logic;
signal \N__41760\ : std_logic;
signal \N__41757\ : std_logic;
signal \N__41752\ : std_logic;
signal \N__41751\ : std_logic;
signal \N__41748\ : std_logic;
signal \N__41745\ : std_logic;
signal \N__41744\ : std_logic;
signal \N__41741\ : std_logic;
signal \N__41738\ : std_logic;
signal \N__41735\ : std_logic;
signal \N__41732\ : std_logic;
signal \N__41729\ : std_logic;
signal \N__41722\ : std_logic;
signal \N__41719\ : std_logic;
signal \N__41718\ : std_logic;
signal \N__41715\ : std_logic;
signal \N__41714\ : std_logic;
signal \N__41711\ : std_logic;
signal \N__41708\ : std_logic;
signal \N__41705\ : std_logic;
signal \N__41698\ : std_logic;
signal \N__41695\ : std_logic;
signal \N__41692\ : std_logic;
signal \N__41691\ : std_logic;
signal \N__41688\ : std_logic;
signal \N__41685\ : std_logic;
signal \N__41684\ : std_logic;
signal \N__41681\ : std_logic;
signal \N__41678\ : std_logic;
signal \N__41675\ : std_logic;
signal \N__41672\ : std_logic;
signal \N__41669\ : std_logic;
signal \N__41664\ : std_logic;
signal \N__41661\ : std_logic;
signal \N__41656\ : std_logic;
signal \N__41653\ : std_logic;
signal \N__41650\ : std_logic;
signal \N__41647\ : std_logic;
signal \N__41646\ : std_logic;
signal \N__41643\ : std_logic;
signal \N__41642\ : std_logic;
signal \N__41639\ : std_logic;
signal \N__41636\ : std_logic;
signal \N__41633\ : std_logic;
signal \N__41626\ : std_logic;
signal \N__41623\ : std_logic;
signal \N__41622\ : std_logic;
signal \N__41619\ : std_logic;
signal \N__41616\ : std_logic;
signal \N__41615\ : std_logic;
signal \N__41614\ : std_logic;
signal \N__41609\ : std_logic;
signal \N__41606\ : std_logic;
signal \N__41603\ : std_logic;
signal \N__41596\ : std_logic;
signal \N__41593\ : std_logic;
signal \N__41592\ : std_logic;
signal \N__41591\ : std_logic;
signal \N__41588\ : std_logic;
signal \N__41585\ : std_logic;
signal \N__41582\ : std_logic;
signal \N__41579\ : std_logic;
signal \N__41576\ : std_logic;
signal \N__41569\ : std_logic;
signal \N__41566\ : std_logic;
signal \N__41565\ : std_logic;
signal \N__41562\ : std_logic;
signal \N__41561\ : std_logic;
signal \N__41558\ : std_logic;
signal \N__41555\ : std_logic;
signal \N__41552\ : std_logic;
signal \N__41545\ : std_logic;
signal \N__41544\ : std_logic;
signal \N__41541\ : std_logic;
signal \N__41536\ : std_logic;
signal \N__41535\ : std_logic;
signal \N__41532\ : std_logic;
signal \N__41529\ : std_logic;
signal \N__41528\ : std_logic;
signal \N__41527\ : std_logic;
signal \N__41526\ : std_logic;
signal \N__41523\ : std_logic;
signal \N__41518\ : std_logic;
signal \N__41515\ : std_logic;
signal \N__41512\ : std_logic;
signal \N__41507\ : std_logic;
signal \N__41506\ : std_logic;
signal \N__41503\ : std_logic;
signal \N__41500\ : std_logic;
signal \N__41497\ : std_logic;
signal \N__41494\ : std_logic;
signal \N__41491\ : std_logic;
signal \N__41488\ : std_logic;
signal \N__41485\ : std_logic;
signal \N__41482\ : std_logic;
signal \N__41477\ : std_logic;
signal \N__41470\ : std_logic;
signal \N__41469\ : std_logic;
signal \N__41466\ : std_logic;
signal \N__41463\ : std_logic;
signal \N__41460\ : std_logic;
signal \N__41457\ : std_logic;
signal \N__41452\ : std_logic;
signal \N__41449\ : std_logic;
signal \N__41446\ : std_logic;
signal \N__41443\ : std_logic;
signal \N__41440\ : std_logic;
signal \N__41437\ : std_logic;
signal \N__41436\ : std_logic;
signal \N__41433\ : std_logic;
signal \N__41430\ : std_logic;
signal \N__41427\ : std_logic;
signal \N__41426\ : std_logic;
signal \N__41425\ : std_logic;
signal \N__41422\ : std_logic;
signal \N__41419\ : std_logic;
signal \N__41416\ : std_logic;
signal \N__41413\ : std_logic;
signal \N__41410\ : std_logic;
signal \N__41405\ : std_logic;
signal \N__41402\ : std_logic;
signal \N__41399\ : std_logic;
signal \N__41396\ : std_logic;
signal \N__41393\ : std_logic;
signal \N__41390\ : std_logic;
signal \N__41387\ : std_logic;
signal \N__41386\ : std_logic;
signal \N__41383\ : std_logic;
signal \N__41378\ : std_logic;
signal \N__41375\ : std_logic;
signal \N__41372\ : std_logic;
signal \N__41365\ : std_logic;
signal \N__41364\ : std_logic;
signal \N__41363\ : std_logic;
signal \N__41360\ : std_logic;
signal \N__41357\ : std_logic;
signal \N__41356\ : std_logic;
signal \N__41355\ : std_logic;
signal \N__41354\ : std_logic;
signal \N__41351\ : std_logic;
signal \N__41348\ : std_logic;
signal \N__41347\ : std_logic;
signal \N__41342\ : std_logic;
signal \N__41339\ : std_logic;
signal \N__41336\ : std_logic;
signal \N__41333\ : std_logic;
signal \N__41330\ : std_logic;
signal \N__41327\ : std_logic;
signal \N__41324\ : std_logic;
signal \N__41321\ : std_logic;
signal \N__41318\ : std_logic;
signal \N__41315\ : std_logic;
signal \N__41312\ : std_logic;
signal \N__41309\ : std_logic;
signal \N__41306\ : std_logic;
signal \N__41303\ : std_logic;
signal \N__41300\ : std_logic;
signal \N__41293\ : std_logic;
signal \N__41284\ : std_logic;
signal \N__41283\ : std_logic;
signal \N__41280\ : std_logic;
signal \N__41277\ : std_logic;
signal \N__41274\ : std_logic;
signal \N__41269\ : std_logic;
signal \N__41266\ : std_logic;
signal \N__41263\ : std_logic;
signal \N__41260\ : std_logic;
signal \N__41259\ : std_logic;
signal \N__41256\ : std_logic;
signal \N__41253\ : std_logic;
signal \N__41248\ : std_logic;
signal \N__41245\ : std_logic;
signal \N__41242\ : std_logic;
signal \N__41239\ : std_logic;
signal \N__41236\ : std_logic;
signal \N__41233\ : std_logic;
signal \N__41230\ : std_logic;
signal \N__41227\ : std_logic;
signal \N__41224\ : std_logic;
signal \N__41221\ : std_logic;
signal \N__41218\ : std_logic;
signal \N__41215\ : std_logic;
signal \N__41212\ : std_logic;
signal \N__41209\ : std_logic;
signal \N__41206\ : std_logic;
signal \N__41203\ : std_logic;
signal \N__41200\ : std_logic;
signal \N__41197\ : std_logic;
signal \N__41196\ : std_logic;
signal \N__41193\ : std_logic;
signal \N__41190\ : std_logic;
signal \N__41189\ : std_logic;
signal \N__41186\ : std_logic;
signal \N__41183\ : std_logic;
signal \N__41180\ : std_logic;
signal \N__41177\ : std_logic;
signal \N__41170\ : std_logic;
signal \N__41169\ : std_logic;
signal \N__41166\ : std_logic;
signal \N__41165\ : std_logic;
signal \N__41164\ : std_logic;
signal \N__41161\ : std_logic;
signal \N__41158\ : std_logic;
signal \N__41153\ : std_logic;
signal \N__41150\ : std_logic;
signal \N__41143\ : std_logic;
signal \N__41142\ : std_logic;
signal \N__41141\ : std_logic;
signal \N__41138\ : std_logic;
signal \N__41135\ : std_logic;
signal \N__41134\ : std_logic;
signal \N__41133\ : std_logic;
signal \N__41132\ : std_logic;
signal \N__41131\ : std_logic;
signal \N__41130\ : std_logic;
signal \N__41129\ : std_logic;
signal \N__41126\ : std_logic;
signal \N__41123\ : std_logic;
signal \N__41120\ : std_logic;
signal \N__41117\ : std_logic;
signal \N__41116\ : std_logic;
signal \N__41115\ : std_logic;
signal \N__41112\ : std_logic;
signal \N__41109\ : std_logic;
signal \N__41106\ : std_logic;
signal \N__41103\ : std_logic;
signal \N__41100\ : std_logic;
signal \N__41099\ : std_logic;
signal \N__41098\ : std_logic;
signal \N__41097\ : std_logic;
signal \N__41094\ : std_logic;
signal \N__41087\ : std_logic;
signal \N__41084\ : std_logic;
signal \N__41083\ : std_logic;
signal \N__41082\ : std_logic;
signal \N__41081\ : std_logic;
signal \N__41080\ : std_logic;
signal \N__41079\ : std_logic;
signal \N__41076\ : std_logic;
signal \N__41073\ : std_logic;
signal \N__41070\ : std_logic;
signal \N__41067\ : std_logic;
signal \N__41062\ : std_logic;
signal \N__41059\ : std_logic;
signal \N__41056\ : std_logic;
signal \N__41053\ : std_logic;
signal \N__41046\ : std_logic;
signal \N__41043\ : std_logic;
signal \N__41040\ : std_logic;
signal \N__41037\ : std_logic;
signal \N__41034\ : std_logic;
signal \N__41031\ : std_logic;
signal \N__41026\ : std_logic;
signal \N__41017\ : std_logic;
signal \N__41012\ : std_logic;
signal \N__41009\ : std_logic;
signal \N__41006\ : std_logic;
signal \N__41003\ : std_logic;
signal \N__41000\ : std_logic;
signal \N__40997\ : std_logic;
signal \N__40994\ : std_logic;
signal \N__40987\ : std_logic;
signal \N__40984\ : std_logic;
signal \N__40979\ : std_logic;
signal \N__40970\ : std_logic;
signal \N__40967\ : std_logic;
signal \N__40962\ : std_logic;
signal \N__40961\ : std_logic;
signal \N__40958\ : std_logic;
signal \N__40955\ : std_logic;
signal \N__40952\ : std_logic;
signal \N__40945\ : std_logic;
signal \N__40942\ : std_logic;
signal \N__40939\ : std_logic;
signal \N__40938\ : std_logic;
signal \N__40935\ : std_logic;
signal \N__40932\ : std_logic;
signal \N__40929\ : std_logic;
signal \N__40928\ : std_logic;
signal \N__40925\ : std_logic;
signal \N__40922\ : std_logic;
signal \N__40919\ : std_logic;
signal \N__40916\ : std_logic;
signal \N__40913\ : std_logic;
signal \N__40910\ : std_logic;
signal \N__40907\ : std_logic;
signal \N__40906\ : std_logic;
signal \N__40901\ : std_logic;
signal \N__40898\ : std_logic;
signal \N__40895\ : std_logic;
signal \N__40888\ : std_logic;
signal \N__40885\ : std_logic;
signal \N__40882\ : std_logic;
signal \N__40881\ : std_logic;
signal \N__40878\ : std_logic;
signal \N__40875\ : std_logic;
signal \N__40872\ : std_logic;
signal \N__40869\ : std_logic;
signal \N__40864\ : std_logic;
signal \N__40861\ : std_logic;
signal \N__40860\ : std_logic;
signal \N__40857\ : std_logic;
signal \N__40854\ : std_logic;
signal \N__40853\ : std_logic;
signal \N__40850\ : std_logic;
signal \N__40847\ : std_logic;
signal \N__40844\ : std_logic;
signal \N__40841\ : std_logic;
signal \N__40838\ : std_logic;
signal \N__40831\ : std_logic;
signal \N__40828\ : std_logic;
signal \N__40825\ : std_logic;
signal \N__40822\ : std_logic;
signal \N__40819\ : std_logic;
signal \N__40816\ : std_logic;
signal \N__40813\ : std_logic;
signal \N__40810\ : std_logic;
signal \N__40807\ : std_logic;
signal \N__40804\ : std_logic;
signal \N__40801\ : std_logic;
signal \N__40798\ : std_logic;
signal \N__40795\ : std_logic;
signal \N__40792\ : std_logic;
signal \N__40789\ : std_logic;
signal \N__40786\ : std_logic;
signal \N__40785\ : std_logic;
signal \N__40784\ : std_logic;
signal \N__40781\ : std_logic;
signal \N__40778\ : std_logic;
signal \N__40775\ : std_logic;
signal \N__40772\ : std_logic;
signal \N__40769\ : std_logic;
signal \N__40766\ : std_logic;
signal \N__40763\ : std_logic;
signal \N__40760\ : std_logic;
signal \N__40757\ : std_logic;
signal \N__40750\ : std_logic;
signal \N__40747\ : std_logic;
signal \N__40744\ : std_logic;
signal \N__40741\ : std_logic;
signal \N__40738\ : std_logic;
signal \N__40735\ : std_logic;
signal \N__40732\ : std_logic;
signal \N__40729\ : std_logic;
signal \N__40726\ : std_logic;
signal \N__40723\ : std_logic;
signal \N__40720\ : std_logic;
signal \N__40717\ : std_logic;
signal \N__40714\ : std_logic;
signal \N__40711\ : std_logic;
signal \N__40708\ : std_logic;
signal \N__40705\ : std_logic;
signal \N__40702\ : std_logic;
signal \N__40699\ : std_logic;
signal \N__40696\ : std_logic;
signal \N__40693\ : std_logic;
signal \N__40690\ : std_logic;
signal \N__40687\ : std_logic;
signal \N__40684\ : std_logic;
signal \N__40683\ : std_logic;
signal \N__40680\ : std_logic;
signal \N__40677\ : std_logic;
signal \N__40674\ : std_logic;
signal \N__40671\ : std_logic;
signal \N__40668\ : std_logic;
signal \N__40665\ : std_logic;
signal \N__40660\ : std_logic;
signal \N__40657\ : std_logic;
signal \N__40654\ : std_logic;
signal \N__40651\ : std_logic;
signal \N__40648\ : std_logic;
signal \N__40645\ : std_logic;
signal \N__40642\ : std_logic;
signal \N__40641\ : std_logic;
signal \N__40638\ : std_logic;
signal \N__40635\ : std_logic;
signal \N__40632\ : std_logic;
signal \N__40629\ : std_logic;
signal \N__40626\ : std_logic;
signal \N__40621\ : std_logic;
signal \N__40618\ : std_logic;
signal \N__40615\ : std_logic;
signal \N__40612\ : std_logic;
signal \N__40609\ : std_logic;
signal \N__40606\ : std_logic;
signal \N__40603\ : std_logic;
signal \N__40600\ : std_logic;
signal \N__40597\ : std_logic;
signal \N__40594\ : std_logic;
signal \N__40591\ : std_logic;
signal \N__40588\ : std_logic;
signal \N__40585\ : std_logic;
signal \N__40582\ : std_logic;
signal \N__40579\ : std_logic;
signal \N__40576\ : std_logic;
signal \N__40573\ : std_logic;
signal \N__40570\ : std_logic;
signal \N__40567\ : std_logic;
signal \N__40564\ : std_logic;
signal \N__40561\ : std_logic;
signal \N__40558\ : std_logic;
signal \N__40555\ : std_logic;
signal \N__40552\ : std_logic;
signal \N__40551\ : std_logic;
signal \N__40548\ : std_logic;
signal \N__40545\ : std_logic;
signal \N__40542\ : std_logic;
signal \N__40539\ : std_logic;
signal \N__40536\ : std_logic;
signal \N__40533\ : std_logic;
signal \N__40530\ : std_logic;
signal \N__40527\ : std_logic;
signal \N__40524\ : std_logic;
signal \N__40523\ : std_logic;
signal \N__40520\ : std_logic;
signal \N__40517\ : std_logic;
signal \N__40514\ : std_logic;
signal \N__40511\ : std_logic;
signal \N__40508\ : std_logic;
signal \N__40501\ : std_logic;
signal \N__40498\ : std_logic;
signal \N__40495\ : std_logic;
signal \N__40492\ : std_logic;
signal \N__40489\ : std_logic;
signal \N__40486\ : std_logic;
signal \N__40483\ : std_logic;
signal \N__40480\ : std_logic;
signal \N__40477\ : std_logic;
signal \N__40474\ : std_logic;
signal \N__40471\ : std_logic;
signal \N__40468\ : std_logic;
signal \N__40465\ : std_logic;
signal \N__40462\ : std_logic;
signal \N__40459\ : std_logic;
signal \N__40456\ : std_logic;
signal \N__40453\ : std_logic;
signal \N__40450\ : std_logic;
signal \N__40447\ : std_logic;
signal \N__40446\ : std_logic;
signal \N__40443\ : std_logic;
signal \N__40440\ : std_logic;
signal \N__40437\ : std_logic;
signal \N__40434\ : std_logic;
signal \N__40431\ : std_logic;
signal \N__40428\ : std_logic;
signal \N__40425\ : std_logic;
signal \N__40422\ : std_logic;
signal \N__40419\ : std_logic;
signal \N__40416\ : std_logic;
signal \N__40413\ : std_logic;
signal \N__40412\ : std_logic;
signal \N__40409\ : std_logic;
signal \N__40406\ : std_logic;
signal \N__40403\ : std_logic;
signal \N__40400\ : std_logic;
signal \N__40397\ : std_logic;
signal \N__40390\ : std_logic;
signal \N__40387\ : std_logic;
signal \N__40384\ : std_logic;
signal \N__40381\ : std_logic;
signal \N__40378\ : std_logic;
signal \N__40375\ : std_logic;
signal \N__40374\ : std_logic;
signal \N__40373\ : std_logic;
signal \N__40370\ : std_logic;
signal \N__40367\ : std_logic;
signal \N__40364\ : std_logic;
signal \N__40361\ : std_logic;
signal \N__40358\ : std_logic;
signal \N__40355\ : std_logic;
signal \N__40352\ : std_logic;
signal \N__40349\ : std_logic;
signal \N__40342\ : std_logic;
signal \N__40339\ : std_logic;
signal \N__40336\ : std_logic;
signal \N__40333\ : std_logic;
signal \N__40330\ : std_logic;
signal \N__40329\ : std_logic;
signal \N__40326\ : std_logic;
signal \N__40323\ : std_logic;
signal \N__40320\ : std_logic;
signal \N__40317\ : std_logic;
signal \N__40316\ : std_logic;
signal \N__40315\ : std_logic;
signal \N__40314\ : std_logic;
signal \N__40311\ : std_logic;
signal \N__40308\ : std_logic;
signal \N__40305\ : std_logic;
signal \N__40302\ : std_logic;
signal \N__40299\ : std_logic;
signal \N__40288\ : std_logic;
signal \N__40285\ : std_logic;
signal \N__40282\ : std_logic;
signal \N__40279\ : std_logic;
signal \N__40276\ : std_logic;
signal \N__40275\ : std_logic;
signal \N__40274\ : std_logic;
signal \N__40271\ : std_logic;
signal \N__40266\ : std_logic;
signal \N__40261\ : std_logic;
signal \N__40260\ : std_logic;
signal \N__40257\ : std_logic;
signal \N__40256\ : std_logic;
signal \N__40253\ : std_logic;
signal \N__40250\ : std_logic;
signal \N__40247\ : std_logic;
signal \N__40242\ : std_logic;
signal \N__40239\ : std_logic;
signal \N__40234\ : std_logic;
signal \N__40231\ : std_logic;
signal \N__40230\ : std_logic;
signal \N__40229\ : std_logic;
signal \N__40226\ : std_logic;
signal \N__40223\ : std_logic;
signal \N__40220\ : std_logic;
signal \N__40213\ : std_logic;
signal \N__40210\ : std_logic;
signal \N__40209\ : std_logic;
signal \N__40206\ : std_logic;
signal \N__40203\ : std_logic;
signal \N__40200\ : std_logic;
signal \N__40197\ : std_logic;
signal \N__40192\ : std_logic;
signal \N__40189\ : std_logic;
signal \N__40186\ : std_logic;
signal \N__40185\ : std_logic;
signal \N__40182\ : std_logic;
signal \N__40179\ : std_logic;
signal \N__40174\ : std_logic;
signal \N__40171\ : std_logic;
signal \N__40168\ : std_logic;
signal \N__40165\ : std_logic;
signal \N__40162\ : std_logic;
signal \N__40159\ : std_logic;
signal \N__40156\ : std_logic;
signal \N__40153\ : std_logic;
signal \N__40150\ : std_logic;
signal \N__40147\ : std_logic;
signal \N__40144\ : std_logic;
signal \N__40141\ : std_logic;
signal \N__40138\ : std_logic;
signal \N__40135\ : std_logic;
signal \N__40132\ : std_logic;
signal \N__40129\ : std_logic;
signal \N__40126\ : std_logic;
signal \N__40125\ : std_logic;
signal \N__40122\ : std_logic;
signal \N__40119\ : std_logic;
signal \N__40116\ : std_logic;
signal \N__40113\ : std_logic;
signal \N__40110\ : std_logic;
signal \N__40107\ : std_logic;
signal \N__40104\ : std_logic;
signal \N__40101\ : std_logic;
signal \N__40098\ : std_logic;
signal \N__40097\ : std_logic;
signal \N__40094\ : std_logic;
signal \N__40091\ : std_logic;
signal \N__40088\ : std_logic;
signal \N__40085\ : std_logic;
signal \N__40082\ : std_logic;
signal \N__40079\ : std_logic;
signal \N__40074\ : std_logic;
signal \N__40069\ : std_logic;
signal \N__40066\ : std_logic;
signal \N__40063\ : std_logic;
signal \N__40060\ : std_logic;
signal \N__40057\ : std_logic;
signal \N__40054\ : std_logic;
signal \N__40051\ : std_logic;
signal \N__40048\ : std_logic;
signal \N__40045\ : std_logic;
signal \N__40042\ : std_logic;
signal \N__40039\ : std_logic;
signal \N__40036\ : std_logic;
signal \N__40033\ : std_logic;
signal \N__40030\ : std_logic;
signal \N__40027\ : std_logic;
signal \N__40024\ : std_logic;
signal \N__40021\ : std_logic;
signal \N__40020\ : std_logic;
signal \N__40017\ : std_logic;
signal \N__40014\ : std_logic;
signal \N__40011\ : std_logic;
signal \N__40008\ : std_logic;
signal \N__40005\ : std_logic;
signal \N__40002\ : std_logic;
signal \N__39999\ : std_logic;
signal \N__39996\ : std_logic;
signal \N__39993\ : std_logic;
signal \N__39990\ : std_logic;
signal \N__39987\ : std_logic;
signal \N__39986\ : std_logic;
signal \N__39983\ : std_logic;
signal \N__39980\ : std_logic;
signal \N__39977\ : std_logic;
signal \N__39972\ : std_logic;
signal \N__39967\ : std_logic;
signal \N__39964\ : std_logic;
signal \N__39961\ : std_logic;
signal \N__39958\ : std_logic;
signal \N__39955\ : std_logic;
signal \N__39952\ : std_logic;
signal \N__39949\ : std_logic;
signal \N__39946\ : std_logic;
signal \N__39943\ : std_logic;
signal \N__39940\ : std_logic;
signal \N__39937\ : std_logic;
signal \N__39934\ : std_logic;
signal \N__39931\ : std_logic;
signal \N__39928\ : std_logic;
signal \N__39925\ : std_logic;
signal \N__39922\ : std_logic;
signal \N__39919\ : std_logic;
signal \N__39916\ : std_logic;
signal \N__39915\ : std_logic;
signal \N__39912\ : std_logic;
signal \N__39909\ : std_logic;
signal \N__39906\ : std_logic;
signal \N__39903\ : std_logic;
signal \N__39900\ : std_logic;
signal \N__39897\ : std_logic;
signal \N__39894\ : std_logic;
signal \N__39891\ : std_logic;
signal \N__39888\ : std_logic;
signal \N__39885\ : std_logic;
signal \N__39882\ : std_logic;
signal \N__39881\ : std_logic;
signal \N__39878\ : std_logic;
signal \N__39875\ : std_logic;
signal \N__39872\ : std_logic;
signal \N__39869\ : std_logic;
signal \N__39866\ : std_logic;
signal \N__39859\ : std_logic;
signal \N__39856\ : std_logic;
signal \N__39853\ : std_logic;
signal \N__39850\ : std_logic;
signal \N__39847\ : std_logic;
signal \N__39844\ : std_logic;
signal \N__39841\ : std_logic;
signal \N__39838\ : std_logic;
signal \N__39835\ : std_logic;
signal \N__39832\ : std_logic;
signal \N__39829\ : std_logic;
signal \N__39826\ : std_logic;
signal \N__39823\ : std_logic;
signal \N__39820\ : std_logic;
signal \N__39817\ : std_logic;
signal \N__39814\ : std_logic;
signal \N__39813\ : std_logic;
signal \N__39810\ : std_logic;
signal \N__39807\ : std_logic;
signal \N__39804\ : std_logic;
signal \N__39801\ : std_logic;
signal \N__39798\ : std_logic;
signal \N__39795\ : std_logic;
signal \N__39792\ : std_logic;
signal \N__39789\ : std_logic;
signal \N__39786\ : std_logic;
signal \N__39783\ : std_logic;
signal \N__39780\ : std_logic;
signal \N__39779\ : std_logic;
signal \N__39776\ : std_logic;
signal \N__39773\ : std_logic;
signal \N__39770\ : std_logic;
signal \N__39767\ : std_logic;
signal \N__39764\ : std_logic;
signal \N__39757\ : std_logic;
signal \N__39754\ : std_logic;
signal \N__39751\ : std_logic;
signal \N__39748\ : std_logic;
signal \N__39745\ : std_logic;
signal \N__39742\ : std_logic;
signal \N__39739\ : std_logic;
signal \N__39736\ : std_logic;
signal \N__39733\ : std_logic;
signal \N__39730\ : std_logic;
signal \N__39727\ : std_logic;
signal \N__39724\ : std_logic;
signal \N__39721\ : std_logic;
signal \N__39718\ : std_logic;
signal \N__39715\ : std_logic;
signal \N__39712\ : std_logic;
signal \N__39709\ : std_logic;
signal \N__39706\ : std_logic;
signal \N__39705\ : std_logic;
signal \N__39702\ : std_logic;
signal \N__39699\ : std_logic;
signal \N__39696\ : std_logic;
signal \N__39693\ : std_logic;
signal \N__39690\ : std_logic;
signal \N__39687\ : std_logic;
signal \N__39684\ : std_logic;
signal \N__39681\ : std_logic;
signal \N__39678\ : std_logic;
signal \N__39675\ : std_logic;
signal \N__39672\ : std_logic;
signal \N__39671\ : std_logic;
signal \N__39668\ : std_logic;
signal \N__39665\ : std_logic;
signal \N__39662\ : std_logic;
signal \N__39659\ : std_logic;
signal \N__39656\ : std_logic;
signal \N__39649\ : std_logic;
signal \N__39646\ : std_logic;
signal \N__39643\ : std_logic;
signal \N__39640\ : std_logic;
signal \N__39637\ : std_logic;
signal \N__39634\ : std_logic;
signal \N__39631\ : std_logic;
signal \N__39628\ : std_logic;
signal \N__39625\ : std_logic;
signal \N__39622\ : std_logic;
signal \N__39619\ : std_logic;
signal \N__39616\ : std_logic;
signal \N__39613\ : std_logic;
signal \N__39610\ : std_logic;
signal \N__39607\ : std_logic;
signal \N__39604\ : std_logic;
signal \N__39601\ : std_logic;
signal \N__39598\ : std_logic;
signal \N__39597\ : std_logic;
signal \N__39594\ : std_logic;
signal \N__39591\ : std_logic;
signal \N__39588\ : std_logic;
signal \N__39585\ : std_logic;
signal \N__39582\ : std_logic;
signal \N__39579\ : std_logic;
signal \N__39576\ : std_logic;
signal \N__39573\ : std_logic;
signal \N__39570\ : std_logic;
signal \N__39567\ : std_logic;
signal \N__39564\ : std_logic;
signal \N__39563\ : std_logic;
signal \N__39560\ : std_logic;
signal \N__39557\ : std_logic;
signal \N__39554\ : std_logic;
signal \N__39551\ : std_logic;
signal \N__39548\ : std_logic;
signal \N__39541\ : std_logic;
signal \N__39538\ : std_logic;
signal \N__39535\ : std_logic;
signal \N__39532\ : std_logic;
signal \N__39529\ : std_logic;
signal \N__39526\ : std_logic;
signal \N__39523\ : std_logic;
signal \N__39520\ : std_logic;
signal \N__39517\ : std_logic;
signal \N__39514\ : std_logic;
signal \N__39511\ : std_logic;
signal \N__39508\ : std_logic;
signal \N__39505\ : std_logic;
signal \N__39502\ : std_logic;
signal \N__39499\ : std_logic;
signal \N__39496\ : std_logic;
signal \N__39493\ : std_logic;
signal \N__39492\ : std_logic;
signal \N__39489\ : std_logic;
signal \N__39486\ : std_logic;
signal \N__39483\ : std_logic;
signal \N__39480\ : std_logic;
signal \N__39477\ : std_logic;
signal \N__39474\ : std_logic;
signal \N__39471\ : std_logic;
signal \N__39468\ : std_logic;
signal \N__39465\ : std_logic;
signal \N__39462\ : std_logic;
signal \N__39459\ : std_logic;
signal \N__39458\ : std_logic;
signal \N__39455\ : std_logic;
signal \N__39452\ : std_logic;
signal \N__39449\ : std_logic;
signal \N__39446\ : std_logic;
signal \N__39443\ : std_logic;
signal \N__39436\ : std_logic;
signal \N__39433\ : std_logic;
signal \N__39430\ : std_logic;
signal \N__39427\ : std_logic;
signal \N__39424\ : std_logic;
signal \N__39421\ : std_logic;
signal \N__39418\ : std_logic;
signal \N__39415\ : std_logic;
signal \N__39412\ : std_logic;
signal \N__39409\ : std_logic;
signal \N__39406\ : std_logic;
signal \N__39403\ : std_logic;
signal \N__39400\ : std_logic;
signal \N__39397\ : std_logic;
signal \N__39394\ : std_logic;
signal \N__39391\ : std_logic;
signal \N__39390\ : std_logic;
signal \N__39387\ : std_logic;
signal \N__39384\ : std_logic;
signal \N__39381\ : std_logic;
signal \N__39378\ : std_logic;
signal \N__39375\ : std_logic;
signal \N__39372\ : std_logic;
signal \N__39369\ : std_logic;
signal \N__39366\ : std_logic;
signal \N__39363\ : std_logic;
signal \N__39360\ : std_logic;
signal \N__39357\ : std_logic;
signal \N__39356\ : std_logic;
signal \N__39353\ : std_logic;
signal \N__39350\ : std_logic;
signal \N__39347\ : std_logic;
signal \N__39344\ : std_logic;
signal \N__39341\ : std_logic;
signal \N__39334\ : std_logic;
signal \N__39331\ : std_logic;
signal \N__39330\ : std_logic;
signal \N__39329\ : std_logic;
signal \N__39328\ : std_logic;
signal \N__39327\ : std_logic;
signal \N__39324\ : std_logic;
signal \N__39323\ : std_logic;
signal \N__39318\ : std_logic;
signal \N__39317\ : std_logic;
signal \N__39316\ : std_logic;
signal \N__39315\ : std_logic;
signal \N__39314\ : std_logic;
signal \N__39313\ : std_logic;
signal \N__39308\ : std_logic;
signal \N__39303\ : std_logic;
signal \N__39300\ : std_logic;
signal \N__39293\ : std_logic;
signal \N__39288\ : std_logic;
signal \N__39287\ : std_logic;
signal \N__39286\ : std_logic;
signal \N__39285\ : std_logic;
signal \N__39280\ : std_logic;
signal \N__39277\ : std_logic;
signal \N__39274\ : std_logic;
signal \N__39273\ : std_logic;
signal \N__39272\ : std_logic;
signal \N__39269\ : std_logic;
signal \N__39262\ : std_logic;
signal \N__39255\ : std_logic;
signal \N__39250\ : std_logic;
signal \N__39241\ : std_logic;
signal \N__39240\ : std_logic;
signal \N__39239\ : std_logic;
signal \N__39238\ : std_logic;
signal \N__39237\ : std_logic;
signal \N__39236\ : std_logic;
signal \N__39233\ : std_logic;
signal \N__39226\ : std_logic;
signal \N__39223\ : std_logic;
signal \N__39220\ : std_logic;
signal \N__39219\ : std_logic;
signal \N__39212\ : std_logic;
signal \N__39209\ : std_logic;
signal \N__39206\ : std_logic;
signal \N__39205\ : std_logic;
signal \N__39198\ : std_logic;
signal \N__39195\ : std_logic;
signal \N__39190\ : std_logic;
signal \N__39187\ : std_logic;
signal \N__39184\ : std_logic;
signal \N__39183\ : std_logic;
signal \N__39180\ : std_logic;
signal \N__39177\ : std_logic;
signal \N__39174\ : std_logic;
signal \N__39171\ : std_logic;
signal \N__39168\ : std_logic;
signal \N__39165\ : std_logic;
signal \N__39160\ : std_logic;
signal \N__39157\ : std_logic;
signal \N__39156\ : std_logic;
signal \N__39153\ : std_logic;
signal \N__39152\ : std_logic;
signal \N__39151\ : std_logic;
signal \N__39150\ : std_logic;
signal \N__39143\ : std_logic;
signal \N__39142\ : std_logic;
signal \N__39141\ : std_logic;
signal \N__39138\ : std_logic;
signal \N__39137\ : std_logic;
signal \N__39134\ : std_logic;
signal \N__39131\ : std_logic;
signal \N__39128\ : std_logic;
signal \N__39123\ : std_logic;
signal \N__39122\ : std_logic;
signal \N__39119\ : std_logic;
signal \N__39116\ : std_logic;
signal \N__39109\ : std_logic;
signal \N__39108\ : std_logic;
signal \N__39107\ : std_logic;
signal \N__39106\ : std_logic;
signal \N__39105\ : std_logic;
signal \N__39102\ : std_logic;
signal \N__39099\ : std_logic;
signal \N__39094\ : std_logic;
signal \N__39089\ : std_logic;
signal \N__39086\ : std_logic;
signal \N__39081\ : std_logic;
signal \N__39076\ : std_logic;
signal \N__39073\ : std_logic;
signal \N__39064\ : std_logic;
signal \N__39063\ : std_logic;
signal \N__39058\ : std_logic;
signal \N__39057\ : std_logic;
signal \N__39054\ : std_logic;
signal \N__39051\ : std_logic;
signal \N__39048\ : std_logic;
signal \N__39043\ : std_logic;
signal \N__39040\ : std_logic;
signal \N__39037\ : std_logic;
signal \N__39034\ : std_logic;
signal \N__39031\ : std_logic;
signal \N__39028\ : std_logic;
signal \N__39025\ : std_logic;
signal \N__39022\ : std_logic;
signal \N__39019\ : std_logic;
signal \N__39016\ : std_logic;
signal \N__39013\ : std_logic;
signal \N__39010\ : std_logic;
signal \N__39007\ : std_logic;
signal \N__39004\ : std_logic;
signal \N__39001\ : std_logic;
signal \N__38998\ : std_logic;
signal \N__38995\ : std_logic;
signal \N__38992\ : std_logic;
signal \N__38991\ : std_logic;
signal \N__38988\ : std_logic;
signal \N__38985\ : std_logic;
signal \N__38982\ : std_logic;
signal \N__38979\ : std_logic;
signal \N__38976\ : std_logic;
signal \N__38973\ : std_logic;
signal \N__38970\ : std_logic;
signal \N__38967\ : std_logic;
signal \N__38964\ : std_logic;
signal \N__38961\ : std_logic;
signal \N__38958\ : std_logic;
signal \N__38955\ : std_logic;
signal \N__38952\ : std_logic;
signal \N__38949\ : std_logic;
signal \N__38946\ : std_logic;
signal \N__38941\ : std_logic;
signal \N__38938\ : std_logic;
signal \N__38937\ : std_logic;
signal \N__38936\ : std_logic;
signal \N__38935\ : std_logic;
signal \N__38932\ : std_logic;
signal \N__38929\ : std_logic;
signal \N__38926\ : std_logic;
signal \N__38923\ : std_logic;
signal \N__38920\ : std_logic;
signal \N__38917\ : std_logic;
signal \N__38914\ : std_logic;
signal \N__38907\ : std_logic;
signal \N__38902\ : std_logic;
signal \N__38899\ : std_logic;
signal \N__38898\ : std_logic;
signal \N__38897\ : std_logic;
signal \N__38894\ : std_logic;
signal \N__38891\ : std_logic;
signal \N__38888\ : std_logic;
signal \N__38885\ : std_logic;
signal \N__38882\ : std_logic;
signal \N__38879\ : std_logic;
signal \N__38874\ : std_logic;
signal \N__38869\ : std_logic;
signal \N__38866\ : std_logic;
signal \N__38865\ : std_logic;
signal \N__38862\ : std_logic;
signal \N__38859\ : std_logic;
signal \N__38856\ : std_logic;
signal \N__38855\ : std_logic;
signal \N__38852\ : std_logic;
signal \N__38849\ : std_logic;
signal \N__38846\ : std_logic;
signal \N__38843\ : std_logic;
signal \N__38838\ : std_logic;
signal \N__38833\ : std_logic;
signal \N__38830\ : std_logic;
signal \N__38827\ : std_logic;
signal \N__38826\ : std_logic;
signal \N__38825\ : std_logic;
signal \N__38822\ : std_logic;
signal \N__38817\ : std_logic;
signal \N__38812\ : std_logic;
signal \N__38809\ : std_logic;
signal \N__38808\ : std_logic;
signal \N__38805\ : std_logic;
signal \N__38802\ : std_logic;
signal \N__38799\ : std_logic;
signal \N__38794\ : std_logic;
signal \N__38791\ : std_logic;
signal \N__38790\ : std_logic;
signal \N__38787\ : std_logic;
signal \N__38784\ : std_logic;
signal \N__38781\ : std_logic;
signal \N__38776\ : std_logic;
signal \N__38773\ : std_logic;
signal \N__38770\ : std_logic;
signal \N__38767\ : std_logic;
signal \N__38764\ : std_logic;
signal \N__38763\ : std_logic;
signal \N__38760\ : std_logic;
signal \N__38759\ : std_logic;
signal \N__38756\ : std_logic;
signal \N__38753\ : std_logic;
signal \N__38750\ : std_logic;
signal \N__38747\ : std_logic;
signal \N__38744\ : std_logic;
signal \N__38741\ : std_logic;
signal \N__38734\ : std_logic;
signal \N__38733\ : std_logic;
signal \N__38732\ : std_logic;
signal \N__38731\ : std_logic;
signal \N__38730\ : std_logic;
signal \N__38729\ : std_logic;
signal \N__38726\ : std_logic;
signal \N__38723\ : std_logic;
signal \N__38720\ : std_logic;
signal \N__38719\ : std_logic;
signal \N__38716\ : std_logic;
signal \N__38713\ : std_logic;
signal \N__38712\ : std_logic;
signal \N__38709\ : std_logic;
signal \N__38706\ : std_logic;
signal \N__38703\ : std_logic;
signal \N__38700\ : std_logic;
signal \N__38697\ : std_logic;
signal \N__38694\ : std_logic;
signal \N__38691\ : std_logic;
signal \N__38688\ : std_logic;
signal \N__38685\ : std_logic;
signal \N__38682\ : std_logic;
signal \N__38679\ : std_logic;
signal \N__38676\ : std_logic;
signal \N__38673\ : std_logic;
signal \N__38668\ : std_logic;
signal \N__38665\ : std_logic;
signal \N__38662\ : std_logic;
signal \N__38659\ : std_logic;
signal \N__38654\ : std_logic;
signal \N__38651\ : std_logic;
signal \N__38650\ : std_logic;
signal \N__38645\ : std_logic;
signal \N__38640\ : std_logic;
signal \N__38635\ : std_logic;
signal \N__38632\ : std_logic;
signal \N__38623\ : std_logic;
signal \N__38620\ : std_logic;
signal \N__38617\ : std_logic;
signal \N__38614\ : std_logic;
signal \N__38613\ : std_logic;
signal \N__38612\ : std_logic;
signal \N__38609\ : std_logic;
signal \N__38606\ : std_logic;
signal \N__38603\ : std_logic;
signal \N__38600\ : std_logic;
signal \N__38597\ : std_logic;
signal \N__38590\ : std_logic;
signal \N__38587\ : std_logic;
signal \N__38584\ : std_logic;
signal \N__38581\ : std_logic;
signal \N__38580\ : std_logic;
signal \N__38577\ : std_logic;
signal \N__38574\ : std_logic;
signal \N__38571\ : std_logic;
signal \N__38568\ : std_logic;
signal \N__38565\ : std_logic;
signal \N__38562\ : std_logic;
signal \N__38557\ : std_logic;
signal \N__38554\ : std_logic;
signal \N__38551\ : std_logic;
signal \N__38550\ : std_logic;
signal \N__38547\ : std_logic;
signal \N__38546\ : std_logic;
signal \N__38545\ : std_logic;
signal \N__38544\ : std_logic;
signal \N__38541\ : std_logic;
signal \N__38540\ : std_logic;
signal \N__38537\ : std_logic;
signal \N__38534\ : std_logic;
signal \N__38533\ : std_logic;
signal \N__38530\ : std_logic;
signal \N__38527\ : std_logic;
signal \N__38524\ : std_logic;
signal \N__38523\ : std_logic;
signal \N__38520\ : std_logic;
signal \N__38515\ : std_logic;
signal \N__38512\ : std_logic;
signal \N__38509\ : std_logic;
signal \N__38504\ : std_logic;
signal \N__38501\ : std_logic;
signal \N__38498\ : std_logic;
signal \N__38497\ : std_logic;
signal \N__38494\ : std_logic;
signal \N__38487\ : std_logic;
signal \N__38482\ : std_logic;
signal \N__38479\ : std_logic;
signal \N__38470\ : std_logic;
signal \N__38469\ : std_logic;
signal \N__38466\ : std_logic;
signal \N__38463\ : std_logic;
signal \N__38460\ : std_logic;
signal \N__38457\ : std_logic;
signal \N__38454\ : std_logic;
signal \N__38451\ : std_logic;
signal \N__38446\ : std_logic;
signal \N__38443\ : std_logic;
signal \N__38442\ : std_logic;
signal \N__38439\ : std_logic;
signal \N__38436\ : std_logic;
signal \N__38433\ : std_logic;
signal \N__38430\ : std_logic;
signal \N__38427\ : std_logic;
signal \N__38422\ : std_logic;
signal \N__38419\ : std_logic;
signal \N__38418\ : std_logic;
signal \N__38417\ : std_logic;
signal \N__38414\ : std_logic;
signal \N__38411\ : std_logic;
signal \N__38408\ : std_logic;
signal \N__38405\ : std_logic;
signal \N__38402\ : std_logic;
signal \N__38395\ : std_logic;
signal \N__38394\ : std_logic;
signal \N__38391\ : std_logic;
signal \N__38390\ : std_logic;
signal \N__38387\ : std_logic;
signal \N__38384\ : std_logic;
signal \N__38379\ : std_logic;
signal \N__38374\ : std_logic;
signal \N__38373\ : std_logic;
signal \N__38372\ : std_logic;
signal \N__38369\ : std_logic;
signal \N__38364\ : std_logic;
signal \N__38359\ : std_logic;
signal \N__38356\ : std_logic;
signal \N__38353\ : std_logic;
signal \N__38350\ : std_logic;
signal \N__38347\ : std_logic;
signal \N__38346\ : std_logic;
signal \N__38343\ : std_logic;
signal \N__38340\ : std_logic;
signal \N__38337\ : std_logic;
signal \N__38334\ : std_logic;
signal \N__38329\ : std_logic;
signal \N__38326\ : std_logic;
signal \N__38323\ : std_logic;
signal \N__38320\ : std_logic;
signal \N__38319\ : std_logic;
signal \N__38316\ : std_logic;
signal \N__38313\ : std_logic;
signal \N__38308\ : std_logic;
signal \N__38305\ : std_logic;
signal \N__38304\ : std_logic;
signal \N__38303\ : std_logic;
signal \N__38300\ : std_logic;
signal \N__38297\ : std_logic;
signal \N__38294\ : std_logic;
signal \N__38291\ : std_logic;
signal \N__38288\ : std_logic;
signal \N__38285\ : std_logic;
signal \N__38282\ : std_logic;
signal \N__38275\ : std_logic;
signal \N__38272\ : std_logic;
signal \N__38269\ : std_logic;
signal \N__38266\ : std_logic;
signal \N__38263\ : std_logic;
signal \N__38260\ : std_logic;
signal \N__38259\ : std_logic;
signal \N__38256\ : std_logic;
signal \N__38253\ : std_logic;
signal \N__38250\ : std_logic;
signal \N__38245\ : std_logic;
signal \N__38242\ : std_logic;
signal \N__38239\ : std_logic;
signal \N__38236\ : std_logic;
signal \N__38233\ : std_logic;
signal \N__38230\ : std_logic;
signal \N__38227\ : std_logic;
signal \N__38224\ : std_logic;
signal \N__38221\ : std_logic;
signal \N__38218\ : std_logic;
signal \N__38215\ : std_logic;
signal \N__38212\ : std_logic;
signal \N__38209\ : std_logic;
signal \N__38208\ : std_logic;
signal \N__38203\ : std_logic;
signal \N__38202\ : std_logic;
signal \N__38201\ : std_logic;
signal \N__38198\ : std_logic;
signal \N__38193\ : std_logic;
signal \N__38190\ : std_logic;
signal \N__38185\ : std_logic;
signal \N__38182\ : std_logic;
signal \N__38179\ : std_logic;
signal \N__38176\ : std_logic;
signal \N__38175\ : std_logic;
signal \N__38172\ : std_logic;
signal \N__38169\ : std_logic;
signal \N__38166\ : std_logic;
signal \N__38163\ : std_logic;
signal \N__38162\ : std_logic;
signal \N__38159\ : std_logic;
signal \N__38156\ : std_logic;
signal \N__38153\ : std_logic;
signal \N__38148\ : std_logic;
signal \N__38143\ : std_logic;
signal \N__38140\ : std_logic;
signal \N__38137\ : std_logic;
signal \N__38134\ : std_logic;
signal \N__38131\ : std_logic;
signal \N__38128\ : std_logic;
signal \N__38125\ : std_logic;
signal \N__38122\ : std_logic;
signal \N__38119\ : std_logic;
signal \N__38116\ : std_logic;
signal \N__38113\ : std_logic;
signal \N__38110\ : std_logic;
signal \N__38107\ : std_logic;
signal \N__38104\ : std_logic;
signal \N__38101\ : std_logic;
signal \N__38098\ : std_logic;
signal \N__38095\ : std_logic;
signal \N__38092\ : std_logic;
signal \N__38089\ : std_logic;
signal \N__38086\ : std_logic;
signal \N__38083\ : std_logic;
signal \N__38080\ : std_logic;
signal \N__38077\ : std_logic;
signal \N__38076\ : std_logic;
signal \N__38073\ : std_logic;
signal \N__38070\ : std_logic;
signal \N__38067\ : std_logic;
signal \N__38064\ : std_logic;
signal \N__38061\ : std_logic;
signal \N__38056\ : std_logic;
signal \N__38053\ : std_logic;
signal \N__38050\ : std_logic;
signal \N__38047\ : std_logic;
signal \N__38044\ : std_logic;
signal \N__38041\ : std_logic;
signal \N__38038\ : std_logic;
signal \N__38035\ : std_logic;
signal \N__38032\ : std_logic;
signal \N__38029\ : std_logic;
signal \N__38026\ : std_logic;
signal \N__38023\ : std_logic;
signal \N__38022\ : std_logic;
signal \N__38019\ : std_logic;
signal \N__38018\ : std_logic;
signal \N__38017\ : std_logic;
signal \N__38016\ : std_logic;
signal \N__38013\ : std_logic;
signal \N__38010\ : std_logic;
signal \N__38007\ : std_logic;
signal \N__38004\ : std_logic;
signal \N__38001\ : std_logic;
signal \N__37996\ : std_logic;
signal \N__37995\ : std_logic;
signal \N__37994\ : std_logic;
signal \N__37991\ : std_logic;
signal \N__37988\ : std_logic;
signal \N__37985\ : std_logic;
signal \N__37982\ : std_logic;
signal \N__37981\ : std_logic;
signal \N__37978\ : std_logic;
signal \N__37975\ : std_logic;
signal \N__37972\ : std_logic;
signal \N__37969\ : std_logic;
signal \N__37966\ : std_logic;
signal \N__37963\ : std_logic;
signal \N__37960\ : std_logic;
signal \N__37957\ : std_logic;
signal \N__37954\ : std_logic;
signal \N__37953\ : std_logic;
signal \N__37948\ : std_logic;
signal \N__37941\ : std_logic;
signal \N__37938\ : std_logic;
signal \N__37935\ : std_logic;
signal \N__37932\ : std_logic;
signal \N__37921\ : std_logic;
signal \N__37920\ : std_logic;
signal \N__37917\ : std_logic;
signal \N__37914\ : std_logic;
signal \N__37909\ : std_logic;
signal \N__37906\ : std_logic;
signal \N__37905\ : std_logic;
signal \N__37902\ : std_logic;
signal \N__37899\ : std_logic;
signal \N__37894\ : std_logic;
signal \N__37891\ : std_logic;
signal \N__37888\ : std_logic;
signal \N__37885\ : std_logic;
signal \N__37884\ : std_logic;
signal \N__37879\ : std_logic;
signal \N__37878\ : std_logic;
signal \N__37877\ : std_logic;
signal \N__37876\ : std_logic;
signal \N__37875\ : std_logic;
signal \N__37874\ : std_logic;
signal \N__37873\ : std_logic;
signal \N__37872\ : std_logic;
signal \N__37871\ : std_logic;
signal \N__37870\ : std_logic;
signal \N__37869\ : std_logic;
signal \N__37868\ : std_logic;
signal \N__37865\ : std_logic;
signal \N__37860\ : std_logic;
signal \N__37851\ : std_logic;
signal \N__37848\ : std_logic;
signal \N__37845\ : std_logic;
signal \N__37844\ : std_logic;
signal \N__37841\ : std_logic;
signal \N__37840\ : std_logic;
signal \N__37839\ : std_logic;
signal \N__37838\ : std_logic;
signal \N__37837\ : std_logic;
signal \N__37836\ : std_logic;
signal \N__37835\ : std_logic;
signal \N__37834\ : std_logic;
signal \N__37833\ : std_logic;
signal \N__37832\ : std_logic;
signal \N__37827\ : std_logic;
signal \N__37824\ : std_logic;
signal \N__37817\ : std_logic;
signal \N__37814\ : std_logic;
signal \N__37811\ : std_logic;
signal \N__37808\ : std_logic;
signal \N__37801\ : std_logic;
signal \N__37788\ : std_logic;
signal \N__37787\ : std_logic;
signal \N__37786\ : std_logic;
signal \N__37785\ : std_logic;
signal \N__37784\ : std_logic;
signal \N__37783\ : std_logic;
signal \N__37782\ : std_logic;
signal \N__37781\ : std_logic;
signal \N__37780\ : std_logic;
signal \N__37779\ : std_logic;
signal \N__37776\ : std_logic;
signal \N__37771\ : std_logic;
signal \N__37766\ : std_logic;
signal \N__37759\ : std_logic;
signal \N__37752\ : std_logic;
signal \N__37739\ : std_logic;
signal \N__37726\ : std_logic;
signal \N__37723\ : std_logic;
signal \N__37720\ : std_logic;
signal \N__37719\ : std_logic;
signal \N__37718\ : std_logic;
signal \N__37715\ : std_logic;
signal \N__37712\ : std_logic;
signal \N__37709\ : std_logic;
signal \N__37702\ : std_logic;
signal \N__37699\ : std_logic;
signal \N__37696\ : std_logic;
signal \N__37693\ : std_logic;
signal \N__37690\ : std_logic;
signal \N__37689\ : std_logic;
signal \N__37686\ : std_logic;
signal \N__37683\ : std_logic;
signal \N__37678\ : std_logic;
signal \N__37675\ : std_logic;
signal \N__37672\ : std_logic;
signal \N__37669\ : std_logic;
signal \N__37666\ : std_logic;
signal \N__37663\ : std_logic;
signal \N__37662\ : std_logic;
signal \N__37659\ : std_logic;
signal \N__37656\ : std_logic;
signal \N__37653\ : std_logic;
signal \N__37650\ : std_logic;
signal \N__37645\ : std_logic;
signal \N__37642\ : std_logic;
signal \N__37639\ : std_logic;
signal \N__37636\ : std_logic;
signal \N__37633\ : std_logic;
signal \N__37630\ : std_logic;
signal \N__37629\ : std_logic;
signal \N__37628\ : std_logic;
signal \N__37625\ : std_logic;
signal \N__37620\ : std_logic;
signal \N__37617\ : std_logic;
signal \N__37614\ : std_logic;
signal \N__37609\ : std_logic;
signal \N__37606\ : std_logic;
signal \N__37605\ : std_logic;
signal \N__37604\ : std_logic;
signal \N__37603\ : std_logic;
signal \N__37602\ : std_logic;
signal \N__37599\ : std_logic;
signal \N__37596\ : std_logic;
signal \N__37595\ : std_logic;
signal \N__37594\ : std_logic;
signal \N__37593\ : std_logic;
signal \N__37590\ : std_logic;
signal \N__37587\ : std_logic;
signal \N__37584\ : std_logic;
signal \N__37583\ : std_logic;
signal \N__37582\ : std_logic;
signal \N__37581\ : std_logic;
signal \N__37580\ : std_logic;
signal \N__37577\ : std_logic;
signal \N__37574\ : std_logic;
signal \N__37569\ : std_logic;
signal \N__37566\ : std_logic;
signal \N__37559\ : std_logic;
signal \N__37550\ : std_logic;
signal \N__37547\ : std_logic;
signal \N__37540\ : std_logic;
signal \N__37537\ : std_logic;
signal \N__37528\ : std_logic;
signal \N__37525\ : std_logic;
signal \N__37522\ : std_logic;
signal \N__37519\ : std_logic;
signal \N__37516\ : std_logic;
signal \N__37515\ : std_logic;
signal \N__37512\ : std_logic;
signal \N__37509\ : std_logic;
signal \N__37506\ : std_logic;
signal \N__37501\ : std_logic;
signal \N__37498\ : std_logic;
signal \N__37497\ : std_logic;
signal \N__37494\ : std_logic;
signal \N__37491\ : std_logic;
signal \N__37488\ : std_logic;
signal \N__37483\ : std_logic;
signal \N__37482\ : std_logic;
signal \N__37479\ : std_logic;
signal \N__37476\ : std_logic;
signal \N__37473\ : std_logic;
signal \N__37470\ : std_logic;
signal \N__37467\ : std_logic;
signal \N__37464\ : std_logic;
signal \N__37459\ : std_logic;
signal \N__37456\ : std_logic;
signal \N__37453\ : std_logic;
signal \N__37452\ : std_logic;
signal \N__37449\ : std_logic;
signal \N__37446\ : std_logic;
signal \N__37445\ : std_logic;
signal \N__37444\ : std_logic;
signal \N__37439\ : std_logic;
signal \N__37436\ : std_logic;
signal \N__37433\ : std_logic;
signal \N__37426\ : std_logic;
signal \N__37425\ : std_logic;
signal \N__37424\ : std_logic;
signal \N__37421\ : std_logic;
signal \N__37418\ : std_logic;
signal \N__37415\ : std_logic;
signal \N__37412\ : std_logic;
signal \N__37407\ : std_logic;
signal \N__37404\ : std_logic;
signal \N__37401\ : std_logic;
signal \N__37396\ : std_logic;
signal \N__37395\ : std_logic;
signal \N__37392\ : std_logic;
signal \N__37391\ : std_logic;
signal \N__37388\ : std_logic;
signal \N__37383\ : std_logic;
signal \N__37378\ : std_logic;
signal \N__37377\ : std_logic;
signal \N__37376\ : std_logic;
signal \N__37369\ : std_logic;
signal \N__37366\ : std_logic;
signal \N__37363\ : std_logic;
signal \N__37360\ : std_logic;
signal \N__37357\ : std_logic;
signal \N__37356\ : std_logic;
signal \N__37355\ : std_logic;
signal \N__37350\ : std_logic;
signal \N__37347\ : std_logic;
signal \N__37346\ : std_logic;
signal \N__37343\ : std_logic;
signal \N__37342\ : std_logic;
signal \N__37339\ : std_logic;
signal \N__37336\ : std_logic;
signal \N__37333\ : std_logic;
signal \N__37330\ : std_logic;
signal \N__37325\ : std_logic;
signal \N__37322\ : std_logic;
signal \N__37317\ : std_logic;
signal \N__37314\ : std_logic;
signal \N__37311\ : std_logic;
signal \N__37308\ : std_logic;
signal \N__37305\ : std_logic;
signal \N__37300\ : std_logic;
signal \N__37297\ : std_logic;
signal \N__37294\ : std_logic;
signal \N__37291\ : std_logic;
signal \N__37288\ : std_logic;
signal \N__37287\ : std_logic;
signal \N__37284\ : std_logic;
signal \N__37281\ : std_logic;
signal \N__37278\ : std_logic;
signal \N__37273\ : std_logic;
signal \N__37270\ : std_logic;
signal \N__37269\ : std_logic;
signal \N__37266\ : std_logic;
signal \N__37263\ : std_logic;
signal \N__37258\ : std_logic;
signal \N__37255\ : std_logic;
signal \N__37252\ : std_logic;
signal \N__37251\ : std_logic;
signal \N__37248\ : std_logic;
signal \N__37245\ : std_logic;
signal \N__37240\ : std_logic;
signal \N__37237\ : std_logic;
signal \N__37236\ : std_logic;
signal \N__37233\ : std_logic;
signal \N__37230\ : std_logic;
signal \N__37225\ : std_logic;
signal \N__37222\ : std_logic;
signal \N__37219\ : std_logic;
signal \N__37218\ : std_logic;
signal \N__37215\ : std_logic;
signal \N__37212\ : std_logic;
signal \N__37207\ : std_logic;
signal \N__37204\ : std_logic;
signal \N__37203\ : std_logic;
signal \N__37200\ : std_logic;
signal \N__37197\ : std_logic;
signal \N__37192\ : std_logic;
signal \N__37189\ : std_logic;
signal \N__37186\ : std_logic;
signal \N__37185\ : std_logic;
signal \N__37182\ : std_logic;
signal \N__37179\ : std_logic;
signal \N__37174\ : std_logic;
signal \N__37171\ : std_logic;
signal \N__37170\ : std_logic;
signal \N__37167\ : std_logic;
signal \N__37164\ : std_logic;
signal \N__37159\ : std_logic;
signal \N__37156\ : std_logic;
signal \N__37153\ : std_logic;
signal \N__37150\ : std_logic;
signal \N__37147\ : std_logic;
signal \N__37144\ : std_logic;
signal \N__37141\ : std_logic;
signal \N__37138\ : std_logic;
signal \N__37135\ : std_logic;
signal \N__37132\ : std_logic;
signal \N__37129\ : std_logic;
signal \N__37126\ : std_logic;
signal \N__37125\ : std_logic;
signal \N__37122\ : std_logic;
signal \N__37119\ : std_logic;
signal \N__37114\ : std_logic;
signal \N__37111\ : std_logic;
signal \N__37110\ : std_logic;
signal \N__37107\ : std_logic;
signal \N__37104\ : std_logic;
signal \N__37099\ : std_logic;
signal \N__37096\ : std_logic;
signal \N__37093\ : std_logic;
signal \N__37092\ : std_logic;
signal \N__37089\ : std_logic;
signal \N__37086\ : std_logic;
signal \N__37081\ : std_logic;
signal \N__37078\ : std_logic;
signal \N__37077\ : std_logic;
signal \N__37074\ : std_logic;
signal \N__37071\ : std_logic;
signal \N__37066\ : std_logic;
signal \N__37063\ : std_logic;
signal \N__37062\ : std_logic;
signal \N__37059\ : std_logic;
signal \N__37056\ : std_logic;
signal \N__37053\ : std_logic;
signal \N__37050\ : std_logic;
signal \N__37047\ : std_logic;
signal \N__37042\ : std_logic;
signal \N__37039\ : std_logic;
signal \N__37038\ : std_logic;
signal \N__37035\ : std_logic;
signal \N__37032\ : std_logic;
signal \N__37029\ : std_logic;
signal \N__37024\ : std_logic;
signal \N__37021\ : std_logic;
signal \N__37018\ : std_logic;
signal \N__37017\ : std_logic;
signal \N__37014\ : std_logic;
signal \N__37011\ : std_logic;
signal \N__37006\ : std_logic;
signal \N__37003\ : std_logic;
signal \N__37000\ : std_logic;
signal \N__36997\ : std_logic;
signal \N__36994\ : std_logic;
signal \N__36991\ : std_logic;
signal \N__36988\ : std_logic;
signal \N__36985\ : std_logic;
signal \N__36982\ : std_logic;
signal \N__36979\ : std_logic;
signal \N__36978\ : std_logic;
signal \N__36977\ : std_logic;
signal \N__36974\ : std_logic;
signal \N__36969\ : std_logic;
signal \N__36964\ : std_logic;
signal \N__36961\ : std_logic;
signal \N__36958\ : std_logic;
signal \N__36955\ : std_logic;
signal \N__36952\ : std_logic;
signal \N__36949\ : std_logic;
signal \N__36948\ : std_logic;
signal \N__36947\ : std_logic;
signal \N__36944\ : std_logic;
signal \N__36941\ : std_logic;
signal \N__36938\ : std_logic;
signal \N__36935\ : std_logic;
signal \N__36932\ : std_logic;
signal \N__36925\ : std_logic;
signal \N__36922\ : std_logic;
signal \N__36921\ : std_logic;
signal \N__36920\ : std_logic;
signal \N__36917\ : std_logic;
signal \N__36914\ : std_logic;
signal \N__36911\ : std_logic;
signal \N__36908\ : std_logic;
signal \N__36905\ : std_logic;
signal \N__36898\ : std_logic;
signal \N__36897\ : std_logic;
signal \N__36896\ : std_logic;
signal \N__36895\ : std_logic;
signal \N__36894\ : std_logic;
signal \N__36891\ : std_logic;
signal \N__36888\ : std_logic;
signal \N__36885\ : std_logic;
signal \N__36882\ : std_logic;
signal \N__36881\ : std_logic;
signal \N__36880\ : std_logic;
signal \N__36877\ : std_logic;
signal \N__36874\ : std_logic;
signal \N__36871\ : std_logic;
signal \N__36868\ : std_logic;
signal \N__36865\ : std_logic;
signal \N__36862\ : std_logic;
signal \N__36859\ : std_logic;
signal \N__36858\ : std_logic;
signal \N__36855\ : std_logic;
signal \N__36850\ : std_logic;
signal \N__36843\ : std_logic;
signal \N__36840\ : std_logic;
signal \N__36837\ : std_logic;
signal \N__36834\ : std_logic;
signal \N__36831\ : std_logic;
signal \N__36826\ : std_logic;
signal \N__36823\ : std_logic;
signal \N__36814\ : std_logic;
signal \N__36811\ : std_logic;
signal \N__36808\ : std_logic;
signal \N__36807\ : std_logic;
signal \N__36804\ : std_logic;
signal \N__36803\ : std_logic;
signal \N__36800\ : std_logic;
signal \N__36797\ : std_logic;
signal \N__36796\ : std_logic;
signal \N__36795\ : std_logic;
signal \N__36792\ : std_logic;
signal \N__36791\ : std_logic;
signal \N__36790\ : std_logic;
signal \N__36787\ : std_logic;
signal \N__36784\ : std_logic;
signal \N__36781\ : std_logic;
signal \N__36780\ : std_logic;
signal \N__36777\ : std_logic;
signal \N__36774\ : std_logic;
signal \N__36771\ : std_logic;
signal \N__36768\ : std_logic;
signal \N__36761\ : std_logic;
signal \N__36758\ : std_logic;
signal \N__36755\ : std_logic;
signal \N__36752\ : std_logic;
signal \N__36749\ : std_logic;
signal \N__36742\ : std_logic;
signal \N__36737\ : std_logic;
signal \N__36734\ : std_logic;
signal \N__36731\ : std_logic;
signal \N__36724\ : std_logic;
signal \N__36721\ : std_logic;
signal \N__36718\ : std_logic;
signal \N__36717\ : std_logic;
signal \N__36714\ : std_logic;
signal \N__36713\ : std_logic;
signal \N__36710\ : std_logic;
signal \N__36707\ : std_logic;
signal \N__36704\ : std_logic;
signal \N__36697\ : std_logic;
signal \N__36694\ : std_logic;
signal \N__36691\ : std_logic;
signal \N__36688\ : std_logic;
signal \N__36685\ : std_logic;
signal \N__36682\ : std_logic;
signal \N__36679\ : std_logic;
signal \N__36678\ : std_logic;
signal \N__36675\ : std_logic;
signal \N__36672\ : std_logic;
signal \N__36669\ : std_logic;
signal \N__36664\ : std_logic;
signal \N__36661\ : std_logic;
signal \N__36658\ : std_logic;
signal \N__36657\ : std_logic;
signal \N__36654\ : std_logic;
signal \N__36653\ : std_logic;
signal \N__36650\ : std_logic;
signal \N__36647\ : std_logic;
signal \N__36644\ : std_logic;
signal \N__36637\ : std_logic;
signal \N__36636\ : std_logic;
signal \N__36631\ : std_logic;
signal \N__36628\ : std_logic;
signal \N__36627\ : std_logic;
signal \N__36624\ : std_logic;
signal \N__36621\ : std_logic;
signal \N__36618\ : std_logic;
signal \N__36613\ : std_logic;
signal \N__36612\ : std_logic;
signal \N__36609\ : std_logic;
signal \N__36606\ : std_logic;
signal \N__36603\ : std_logic;
signal \N__36598\ : std_logic;
signal \N__36595\ : std_logic;
signal \N__36592\ : std_logic;
signal \N__36589\ : std_logic;
signal \N__36588\ : std_logic;
signal \N__36587\ : std_logic;
signal \N__36584\ : std_logic;
signal \N__36579\ : std_logic;
signal \N__36574\ : std_logic;
signal \N__36571\ : std_logic;
signal \N__36568\ : std_logic;
signal \N__36565\ : std_logic;
signal \N__36564\ : std_logic;
signal \N__36563\ : std_logic;
signal \N__36560\ : std_logic;
signal \N__36557\ : std_logic;
signal \N__36554\ : std_logic;
signal \N__36551\ : std_logic;
signal \N__36548\ : std_logic;
signal \N__36545\ : std_logic;
signal \N__36538\ : std_logic;
signal \N__36535\ : std_logic;
signal \N__36532\ : std_logic;
signal \N__36529\ : std_logic;
signal \N__36526\ : std_logic;
signal \N__36523\ : std_logic;
signal \N__36520\ : std_logic;
signal \N__36517\ : std_logic;
signal \N__36514\ : std_logic;
signal \N__36511\ : std_logic;
signal \N__36508\ : std_logic;
signal \N__36505\ : std_logic;
signal \N__36502\ : std_logic;
signal \N__36499\ : std_logic;
signal \N__36496\ : std_logic;
signal \N__36493\ : std_logic;
signal \N__36490\ : std_logic;
signal \N__36487\ : std_logic;
signal \N__36484\ : std_logic;
signal \N__36481\ : std_logic;
signal \N__36478\ : std_logic;
signal \N__36477\ : std_logic;
signal \N__36474\ : std_logic;
signal \N__36471\ : std_logic;
signal \N__36468\ : std_logic;
signal \N__36465\ : std_logic;
signal \N__36462\ : std_logic;
signal \N__36459\ : std_logic;
signal \N__36456\ : std_logic;
signal \N__36453\ : std_logic;
signal \N__36450\ : std_logic;
signal \N__36447\ : std_logic;
signal \N__36444\ : std_logic;
signal \N__36441\ : std_logic;
signal \N__36438\ : std_logic;
signal \N__36433\ : std_logic;
signal \N__36430\ : std_logic;
signal \N__36427\ : std_logic;
signal \N__36426\ : std_logic;
signal \N__36423\ : std_logic;
signal \N__36420\ : std_logic;
signal \N__36417\ : std_logic;
signal \N__36412\ : std_logic;
signal \N__36411\ : std_logic;
signal \N__36408\ : std_logic;
signal \N__36405\ : std_logic;
signal \N__36402\ : std_logic;
signal \N__36397\ : std_logic;
signal \N__36396\ : std_logic;
signal \N__36395\ : std_logic;
signal \N__36394\ : std_logic;
signal \N__36391\ : std_logic;
signal \N__36388\ : std_logic;
signal \N__36385\ : std_logic;
signal \N__36382\ : std_logic;
signal \N__36379\ : std_logic;
signal \N__36378\ : std_logic;
signal \N__36375\ : std_logic;
signal \N__36370\ : std_logic;
signal \N__36367\ : std_logic;
signal \N__36364\ : std_logic;
signal \N__36361\ : std_logic;
signal \N__36358\ : std_logic;
signal \N__36353\ : std_logic;
signal \N__36346\ : std_logic;
signal \N__36345\ : std_logic;
signal \N__36340\ : std_logic;
signal \N__36337\ : std_logic;
signal \N__36334\ : std_logic;
signal \N__36333\ : std_logic;
signal \N__36330\ : std_logic;
signal \N__36327\ : std_logic;
signal \N__36324\ : std_logic;
signal \N__36319\ : std_logic;
signal \N__36318\ : std_logic;
signal \N__36315\ : std_logic;
signal \N__36312\ : std_logic;
signal \N__36309\ : std_logic;
signal \N__36304\ : std_logic;
signal \N__36303\ : std_logic;
signal \N__36302\ : std_logic;
signal \N__36299\ : std_logic;
signal \N__36296\ : std_logic;
signal \N__36293\ : std_logic;
signal \N__36290\ : std_logic;
signal \N__36287\ : std_logic;
signal \N__36280\ : std_logic;
signal \N__36277\ : std_logic;
signal \N__36274\ : std_logic;
signal \N__36271\ : std_logic;
signal \N__36268\ : std_logic;
signal \N__36265\ : std_logic;
signal \N__36262\ : std_logic;
signal \N__36259\ : std_logic;
signal \N__36256\ : std_logic;
signal \N__36255\ : std_logic;
signal \N__36254\ : std_logic;
signal \N__36253\ : std_logic;
signal \N__36252\ : std_logic;
signal \N__36249\ : std_logic;
signal \N__36246\ : std_logic;
signal \N__36243\ : std_logic;
signal \N__36242\ : std_logic;
signal \N__36241\ : std_logic;
signal \N__36238\ : std_logic;
signal \N__36237\ : std_logic;
signal \N__36234\ : std_logic;
signal \N__36233\ : std_logic;
signal \N__36228\ : std_logic;
signal \N__36225\ : std_logic;
signal \N__36222\ : std_logic;
signal \N__36219\ : std_logic;
signal \N__36216\ : std_logic;
signal \N__36213\ : std_logic;
signal \N__36210\ : std_logic;
signal \N__36207\ : std_logic;
signal \N__36204\ : std_logic;
signal \N__36199\ : std_logic;
signal \N__36188\ : std_logic;
signal \N__36185\ : std_logic;
signal \N__36182\ : std_logic;
signal \N__36179\ : std_logic;
signal \N__36176\ : std_logic;
signal \N__36171\ : std_logic;
signal \N__36166\ : std_logic;
signal \N__36165\ : std_logic;
signal \N__36164\ : std_logic;
signal \N__36161\ : std_logic;
signal \N__36154\ : std_logic;
signal \N__36151\ : std_logic;
signal \N__36148\ : std_logic;
signal \N__36145\ : std_logic;
signal \N__36144\ : std_logic;
signal \N__36143\ : std_logic;
signal \N__36140\ : std_logic;
signal \N__36137\ : std_logic;
signal \N__36134\ : std_logic;
signal \N__36131\ : std_logic;
signal \N__36124\ : std_logic;
signal \N__36121\ : std_logic;
signal \N__36118\ : std_logic;
signal \N__36115\ : std_logic;
signal \N__36112\ : std_logic;
signal \N__36109\ : std_logic;
signal \N__36108\ : std_logic;
signal \N__36105\ : std_logic;
signal \N__36104\ : std_logic;
signal \N__36101\ : std_logic;
signal \N__36098\ : std_logic;
signal \N__36095\ : std_logic;
signal \N__36088\ : std_logic;
signal \N__36085\ : std_logic;
signal \N__36082\ : std_logic;
signal \N__36079\ : std_logic;
signal \N__36076\ : std_logic;
signal \N__36073\ : std_logic;
signal \N__36070\ : std_logic;
signal \N__36067\ : std_logic;
signal \N__36064\ : std_logic;
signal \N__36061\ : std_logic;
signal \N__36058\ : std_logic;
signal \N__36055\ : std_logic;
signal \N__36052\ : std_logic;
signal \N__36049\ : std_logic;
signal \N__36046\ : std_logic;
signal \N__36043\ : std_logic;
signal \N__36040\ : std_logic;
signal \N__36039\ : std_logic;
signal \N__36036\ : std_logic;
signal \N__36033\ : std_logic;
signal \N__36030\ : std_logic;
signal \N__36025\ : std_logic;
signal \N__36022\ : std_logic;
signal \N__36019\ : std_logic;
signal \N__36016\ : std_logic;
signal \N__36013\ : std_logic;
signal \N__36010\ : std_logic;
signal \N__36007\ : std_logic;
signal \N__36004\ : std_logic;
signal \N__36001\ : std_logic;
signal \N__35998\ : std_logic;
signal \N__35995\ : std_logic;
signal \N__35992\ : std_logic;
signal \N__35991\ : std_logic;
signal \N__35988\ : std_logic;
signal \N__35985\ : std_logic;
signal \N__35982\ : std_logic;
signal \N__35979\ : std_logic;
signal \N__35978\ : std_logic;
signal \N__35977\ : std_logic;
signal \N__35972\ : std_logic;
signal \N__35971\ : std_logic;
signal \N__35968\ : std_logic;
signal \N__35967\ : std_logic;
signal \N__35964\ : std_logic;
signal \N__35961\ : std_logic;
signal \N__35958\ : std_logic;
signal \N__35955\ : std_logic;
signal \N__35952\ : std_logic;
signal \N__35951\ : std_logic;
signal \N__35948\ : std_logic;
signal \N__35943\ : std_logic;
signal \N__35938\ : std_logic;
signal \N__35935\ : std_logic;
signal \N__35934\ : std_logic;
signal \N__35933\ : std_logic;
signal \N__35930\ : std_logic;
signal \N__35927\ : std_logic;
signal \N__35922\ : std_logic;
signal \N__35919\ : std_logic;
signal \N__35916\ : std_logic;
signal \N__35905\ : std_logic;
signal \N__35902\ : std_logic;
signal \N__35899\ : std_logic;
signal \N__35896\ : std_logic;
signal \N__35895\ : std_logic;
signal \N__35892\ : std_logic;
signal \N__35889\ : std_logic;
signal \N__35886\ : std_logic;
signal \N__35881\ : std_logic;
signal \N__35878\ : std_logic;
signal \N__35875\ : std_logic;
signal \N__35872\ : std_logic;
signal \N__35869\ : std_logic;
signal \N__35866\ : std_logic;
signal \N__35863\ : std_logic;
signal \N__35860\ : std_logic;
signal \N__35857\ : std_logic;
signal \N__35856\ : std_logic;
signal \N__35855\ : std_logic;
signal \N__35852\ : std_logic;
signal \N__35849\ : std_logic;
signal \N__35846\ : std_logic;
signal \N__35843\ : std_logic;
signal \N__35838\ : std_logic;
signal \N__35833\ : std_logic;
signal \N__35830\ : std_logic;
signal \N__35827\ : std_logic;
signal \N__35824\ : std_logic;
signal \N__35821\ : std_logic;
signal \N__35818\ : std_logic;
signal \N__35815\ : std_logic;
signal \N__35812\ : std_logic;
signal \N__35811\ : std_logic;
signal \N__35810\ : std_logic;
signal \N__35807\ : std_logic;
signal \N__35806\ : std_logic;
signal \N__35803\ : std_logic;
signal \N__35802\ : std_logic;
signal \N__35799\ : std_logic;
signal \N__35798\ : std_logic;
signal \N__35795\ : std_logic;
signal \N__35792\ : std_logic;
signal \N__35789\ : std_logic;
signal \N__35786\ : std_logic;
signal \N__35783\ : std_logic;
signal \N__35780\ : std_logic;
signal \N__35779\ : std_logic;
signal \N__35776\ : std_logic;
signal \N__35773\ : std_logic;
signal \N__35770\ : std_logic;
signal \N__35767\ : std_logic;
signal \N__35762\ : std_logic;
signal \N__35759\ : std_logic;
signal \N__35758\ : std_logic;
signal \N__35757\ : std_logic;
signal \N__35754\ : std_logic;
signal \N__35751\ : std_logic;
signal \N__35748\ : std_logic;
signal \N__35745\ : std_logic;
signal \N__35742\ : std_logic;
signal \N__35739\ : std_logic;
signal \N__35736\ : std_logic;
signal \N__35733\ : std_logic;
signal \N__35716\ : std_logic;
signal \N__35713\ : std_logic;
signal \N__35710\ : std_logic;
signal \N__35707\ : std_logic;
signal \N__35704\ : std_logic;
signal \N__35701\ : std_logic;
signal \N__35698\ : std_logic;
signal \N__35695\ : std_logic;
signal \N__35692\ : std_logic;
signal \N__35689\ : std_logic;
signal \N__35686\ : std_logic;
signal \N__35683\ : std_logic;
signal \N__35680\ : std_logic;
signal \N__35677\ : std_logic;
signal \N__35674\ : std_logic;
signal \N__35671\ : std_logic;
signal \N__35668\ : std_logic;
signal \N__35665\ : std_logic;
signal \N__35664\ : std_logic;
signal \N__35663\ : std_logic;
signal \N__35662\ : std_logic;
signal \N__35661\ : std_logic;
signal \N__35658\ : std_logic;
signal \N__35655\ : std_logic;
signal \N__35652\ : std_logic;
signal \N__35649\ : std_logic;
signal \N__35646\ : std_logic;
signal \N__35641\ : std_logic;
signal \N__35640\ : std_logic;
signal \N__35637\ : std_logic;
signal \N__35636\ : std_logic;
signal \N__35633\ : std_logic;
signal \N__35628\ : std_logic;
signal \N__35625\ : std_logic;
signal \N__35622\ : std_logic;
signal \N__35619\ : std_logic;
signal \N__35618\ : std_logic;
signal \N__35617\ : std_logic;
signal \N__35614\ : std_logic;
signal \N__35611\ : std_logic;
signal \N__35608\ : std_logic;
signal \N__35603\ : std_logic;
signal \N__35600\ : std_logic;
signal \N__35597\ : std_logic;
signal \N__35584\ : std_logic;
signal \N__35581\ : std_logic;
signal \N__35578\ : std_logic;
signal \N__35575\ : std_logic;
signal \N__35572\ : std_logic;
signal \N__35569\ : std_logic;
signal \N__35568\ : std_logic;
signal \N__35567\ : std_logic;
signal \N__35564\ : std_logic;
signal \N__35563\ : std_logic;
signal \N__35560\ : std_logic;
signal \N__35559\ : std_logic;
signal \N__35558\ : std_logic;
signal \N__35555\ : std_logic;
signal \N__35552\ : std_logic;
signal \N__35549\ : std_logic;
signal \N__35546\ : std_logic;
signal \N__35543\ : std_logic;
signal \N__35540\ : std_logic;
signal \N__35537\ : std_logic;
signal \N__35534\ : std_logic;
signal \N__35531\ : std_logic;
signal \N__35530\ : std_logic;
signal \N__35525\ : std_logic;
signal \N__35522\ : std_logic;
signal \N__35519\ : std_logic;
signal \N__35514\ : std_logic;
signal \N__35511\ : std_logic;
signal \N__35510\ : std_logic;
signal \N__35509\ : std_logic;
signal \N__35502\ : std_logic;
signal \N__35497\ : std_logic;
signal \N__35494\ : std_logic;
signal \N__35491\ : std_logic;
signal \N__35482\ : std_logic;
signal \N__35479\ : std_logic;
signal \N__35476\ : std_logic;
signal \N__35473\ : std_logic;
signal \N__35470\ : std_logic;
signal \N__35467\ : std_logic;
signal \N__35464\ : std_logic;
signal \N__35461\ : std_logic;
signal \N__35458\ : std_logic;
signal \N__35455\ : std_logic;
signal \N__35452\ : std_logic;
signal \N__35451\ : std_logic;
signal \N__35450\ : std_logic;
signal \N__35449\ : std_logic;
signal \N__35448\ : std_logic;
signal \N__35445\ : std_logic;
signal \N__35442\ : std_logic;
signal \N__35441\ : std_logic;
signal \N__35438\ : std_logic;
signal \N__35433\ : std_logic;
signal \N__35428\ : std_logic;
signal \N__35425\ : std_logic;
signal \N__35422\ : std_logic;
signal \N__35421\ : std_logic;
signal \N__35420\ : std_logic;
signal \N__35417\ : std_logic;
signal \N__35414\ : std_logic;
signal \N__35411\ : std_logic;
signal \N__35408\ : std_logic;
signal \N__35405\ : std_logic;
signal \N__35402\ : std_logic;
signal \N__35401\ : std_logic;
signal \N__35398\ : std_logic;
signal \N__35395\ : std_logic;
signal \N__35392\ : std_logic;
signal \N__35387\ : std_logic;
signal \N__35384\ : std_logic;
signal \N__35381\ : std_logic;
signal \N__35368\ : std_logic;
signal \N__35365\ : std_logic;
signal \N__35362\ : std_logic;
signal \N__35359\ : std_logic;
signal \N__35356\ : std_logic;
signal \N__35353\ : std_logic;
signal \N__35350\ : std_logic;
signal \N__35347\ : std_logic;
signal \N__35344\ : std_logic;
signal \N__35341\ : std_logic;
signal \N__35338\ : std_logic;
signal \N__35335\ : std_logic;
signal \N__35332\ : std_logic;
signal \N__35329\ : std_logic;
signal \N__35326\ : std_logic;
signal \N__35325\ : std_logic;
signal \N__35322\ : std_logic;
signal \N__35319\ : std_logic;
signal \N__35316\ : std_logic;
signal \N__35313\ : std_logic;
signal \N__35308\ : std_logic;
signal \N__35305\ : std_logic;
signal \N__35302\ : std_logic;
signal \N__35301\ : std_logic;
signal \N__35298\ : std_logic;
signal \N__35295\ : std_logic;
signal \N__35292\ : std_logic;
signal \N__35289\ : std_logic;
signal \N__35284\ : std_logic;
signal \N__35283\ : std_logic;
signal \N__35280\ : std_logic;
signal \N__35277\ : std_logic;
signal \N__35276\ : std_logic;
signal \N__35273\ : std_logic;
signal \N__35270\ : std_logic;
signal \N__35267\ : std_logic;
signal \N__35264\ : std_logic;
signal \N__35261\ : std_logic;
signal \N__35258\ : std_logic;
signal \N__35255\ : std_logic;
signal \N__35252\ : std_logic;
signal \N__35245\ : std_logic;
signal \N__35242\ : std_logic;
signal \N__35239\ : std_logic;
signal \N__35236\ : std_logic;
signal \N__35233\ : std_logic;
signal \N__35230\ : std_logic;
signal \N__35227\ : std_logic;
signal \N__35224\ : std_logic;
signal \N__35221\ : std_logic;
signal \N__35218\ : std_logic;
signal \N__35215\ : std_logic;
signal \N__35212\ : std_logic;
signal \N__35209\ : std_logic;
signal \N__35206\ : std_logic;
signal \N__35203\ : std_logic;
signal \N__35200\ : std_logic;
signal \N__35197\ : std_logic;
signal \N__35194\ : std_logic;
signal \N__35191\ : std_logic;
signal \N__35188\ : std_logic;
signal \N__35185\ : std_logic;
signal \N__35182\ : std_logic;
signal \N__35179\ : std_logic;
signal \N__35176\ : std_logic;
signal \N__35173\ : std_logic;
signal \N__35170\ : std_logic;
signal \N__35167\ : std_logic;
signal \N__35164\ : std_logic;
signal \N__35161\ : std_logic;
signal \N__35158\ : std_logic;
signal \N__35155\ : std_logic;
signal \N__35152\ : std_logic;
signal \N__35149\ : std_logic;
signal \N__35146\ : std_logic;
signal \N__35143\ : std_logic;
signal \N__35140\ : std_logic;
signal \N__35137\ : std_logic;
signal \N__35134\ : std_logic;
signal \N__35131\ : std_logic;
signal \N__35128\ : std_logic;
signal \N__35125\ : std_logic;
signal \N__35122\ : std_logic;
signal \N__35119\ : std_logic;
signal \N__35116\ : std_logic;
signal \N__35113\ : std_logic;
signal \N__35110\ : std_logic;
signal \N__35107\ : std_logic;
signal \N__35104\ : std_logic;
signal \N__35101\ : std_logic;
signal \N__35098\ : std_logic;
signal \N__35095\ : std_logic;
signal \N__35092\ : std_logic;
signal \N__35089\ : std_logic;
signal \N__35086\ : std_logic;
signal \N__35083\ : std_logic;
signal \N__35082\ : std_logic;
signal \N__35079\ : std_logic;
signal \N__35076\ : std_logic;
signal \N__35073\ : std_logic;
signal \N__35070\ : std_logic;
signal \N__35067\ : std_logic;
signal \N__35062\ : std_logic;
signal \N__35059\ : std_logic;
signal \N__35056\ : std_logic;
signal \N__35053\ : std_logic;
signal \N__35050\ : std_logic;
signal \N__35047\ : std_logic;
signal \N__35044\ : std_logic;
signal \N__35041\ : std_logic;
signal \N__35038\ : std_logic;
signal \N__35035\ : std_logic;
signal \N__35032\ : std_logic;
signal \N__35029\ : std_logic;
signal \N__35026\ : std_logic;
signal \N__35023\ : std_logic;
signal \N__35020\ : std_logic;
signal \N__35017\ : std_logic;
signal \N__35014\ : std_logic;
signal \N__35011\ : std_logic;
signal \N__35008\ : std_logic;
signal \N__35005\ : std_logic;
signal \N__35002\ : std_logic;
signal \N__34999\ : std_logic;
signal \N__34996\ : std_logic;
signal \N__34995\ : std_logic;
signal \N__34994\ : std_logic;
signal \N__34991\ : std_logic;
signal \N__34988\ : std_logic;
signal \N__34985\ : std_logic;
signal \N__34980\ : std_logic;
signal \N__34975\ : std_logic;
signal \N__34974\ : std_logic;
signal \N__34971\ : std_logic;
signal \N__34970\ : std_logic;
signal \N__34967\ : std_logic;
signal \N__34964\ : std_logic;
signal \N__34963\ : std_logic;
signal \N__34962\ : std_logic;
signal \N__34959\ : std_logic;
signal \N__34956\ : std_logic;
signal \N__34953\ : std_logic;
signal \N__34950\ : std_logic;
signal \N__34947\ : std_logic;
signal \N__34936\ : std_logic;
signal \N__34935\ : std_logic;
signal \N__34932\ : std_logic;
signal \N__34931\ : std_logic;
signal \N__34930\ : std_logic;
signal \N__34927\ : std_logic;
signal \N__34922\ : std_logic;
signal \N__34919\ : std_logic;
signal \N__34918\ : std_logic;
signal \N__34915\ : std_logic;
signal \N__34914\ : std_logic;
signal \N__34913\ : std_logic;
signal \N__34908\ : std_logic;
signal \N__34905\ : std_logic;
signal \N__34902\ : std_logic;
signal \N__34897\ : std_logic;
signal \N__34894\ : std_logic;
signal \N__34885\ : std_logic;
signal \N__34882\ : std_logic;
signal \N__34879\ : std_logic;
signal \N__34878\ : std_logic;
signal \N__34877\ : std_logic;
signal \N__34876\ : std_logic;
signal \N__34873\ : std_logic;
signal \N__34872\ : std_logic;
signal \N__34869\ : std_logic;
signal \N__34866\ : std_logic;
signal \N__34865\ : std_logic;
signal \N__34864\ : std_logic;
signal \N__34861\ : std_logic;
signal \N__34858\ : std_logic;
signal \N__34855\ : std_logic;
signal \N__34850\ : std_logic;
signal \N__34847\ : std_logic;
signal \N__34846\ : std_logic;
signal \N__34845\ : std_logic;
signal \N__34844\ : std_logic;
signal \N__34841\ : std_logic;
signal \N__34838\ : std_logic;
signal \N__34835\ : std_logic;
signal \N__34832\ : std_logic;
signal \N__34827\ : std_logic;
signal \N__34820\ : std_logic;
signal \N__34817\ : std_logic;
signal \N__34812\ : std_logic;
signal \N__34805\ : std_logic;
signal \N__34802\ : std_logic;
signal \N__34799\ : std_logic;
signal \N__34796\ : std_logic;
signal \N__34793\ : std_logic;
signal \N__34790\ : std_logic;
signal \N__34787\ : std_logic;
signal \N__34784\ : std_logic;
signal \N__34779\ : std_logic;
signal \N__34774\ : std_logic;
signal \N__34773\ : std_logic;
signal \N__34772\ : std_logic;
signal \N__34771\ : std_logic;
signal \N__34770\ : std_logic;
signal \N__34769\ : std_logic;
signal \N__34768\ : std_logic;
signal \N__34765\ : std_logic;
signal \N__34762\ : std_logic;
signal \N__34755\ : std_logic;
signal \N__34752\ : std_logic;
signal \N__34751\ : std_logic;
signal \N__34748\ : std_logic;
signal \N__34747\ : std_logic;
signal \N__34746\ : std_logic;
signal \N__34745\ : std_logic;
signal \N__34744\ : std_logic;
signal \N__34743\ : std_logic;
signal \N__34742\ : std_logic;
signal \N__34741\ : std_logic;
signal \N__34740\ : std_logic;
signal \N__34739\ : std_logic;
signal \N__34736\ : std_logic;
signal \N__34731\ : std_logic;
signal \N__34728\ : std_logic;
signal \N__34725\ : std_logic;
signal \N__34724\ : std_logic;
signal \N__34723\ : std_logic;
signal \N__34720\ : std_logic;
signal \N__34717\ : std_logic;
signal \N__34716\ : std_logic;
signal \N__34713\ : std_logic;
signal \N__34712\ : std_logic;
signal \N__34709\ : std_logic;
signal \N__34704\ : std_logic;
signal \N__34701\ : std_logic;
signal \N__34698\ : std_logic;
signal \N__34693\ : std_logic;
signal \N__34686\ : std_logic;
signal \N__34679\ : std_logic;
signal \N__34674\ : std_logic;
signal \N__34667\ : std_logic;
signal \N__34648\ : std_logic;
signal \N__34645\ : std_logic;
signal \N__34642\ : std_logic;
signal \N__34641\ : std_logic;
signal \N__34640\ : std_logic;
signal \N__34639\ : std_logic;
signal \N__34638\ : std_logic;
signal \N__34637\ : std_logic;
signal \N__34636\ : std_logic;
signal \N__34635\ : std_logic;
signal \N__34634\ : std_logic;
signal \N__34633\ : std_logic;
signal \N__34632\ : std_logic;
signal \N__34631\ : std_logic;
signal \N__34630\ : std_logic;
signal \N__34629\ : std_logic;
signal \N__34628\ : std_logic;
signal \N__34627\ : std_logic;
signal \N__34626\ : std_logic;
signal \N__34625\ : std_logic;
signal \N__34624\ : std_logic;
signal \N__34621\ : std_logic;
signal \N__34620\ : std_logic;
signal \N__34617\ : std_logic;
signal \N__34602\ : std_logic;
signal \N__34595\ : std_logic;
signal \N__34594\ : std_logic;
signal \N__34593\ : std_logic;
signal \N__34590\ : std_logic;
signal \N__34589\ : std_logic;
signal \N__34588\ : std_logic;
signal \N__34585\ : std_logic;
signal \N__34584\ : std_logic;
signal \N__34575\ : std_logic;
signal \N__34574\ : std_logic;
signal \N__34573\ : std_logic;
signal \N__34572\ : std_logic;
signal \N__34571\ : std_logic;
signal \N__34570\ : std_logic;
signal \N__34569\ : std_logic;
signal \N__34568\ : std_logic;
signal \N__34567\ : std_logic;
signal \N__34566\ : std_logic;
signal \N__34565\ : std_logic;
signal \N__34564\ : std_logic;
signal \N__34563\ : std_logic;
signal \N__34562\ : std_logic;
signal \N__34561\ : std_logic;
signal \N__34556\ : std_logic;
signal \N__34553\ : std_logic;
signal \N__34546\ : std_logic;
signal \N__34541\ : std_logic;
signal \N__34536\ : std_logic;
signal \N__34533\ : std_logic;
signal \N__34530\ : std_logic;
signal \N__34527\ : std_logic;
signal \N__34524\ : std_logic;
signal \N__34507\ : std_logic;
signal \N__34504\ : std_logic;
signal \N__34503\ : std_logic;
signal \N__34500\ : std_logic;
signal \N__34497\ : std_logic;
signal \N__34494\ : std_logic;
signal \N__34491\ : std_logic;
signal \N__34490\ : std_logic;
signal \N__34489\ : std_logic;
signal \N__34488\ : std_logic;
signal \N__34487\ : std_logic;
signal \N__34486\ : std_logic;
signal \N__34485\ : std_logic;
signal \N__34482\ : std_logic;
signal \N__34479\ : std_logic;
signal \N__34476\ : std_logic;
signal \N__34467\ : std_logic;
signal \N__34466\ : std_logic;
signal \N__34465\ : std_logic;
signal \N__34456\ : std_logic;
signal \N__34453\ : std_logic;
signal \N__34446\ : std_logic;
signal \N__34443\ : std_logic;
signal \N__34436\ : std_logic;
signal \N__34425\ : std_logic;
signal \N__34418\ : std_logic;
signal \N__34413\ : std_logic;
signal \N__34406\ : std_logic;
signal \N__34393\ : std_logic;
signal \N__34390\ : std_logic;
signal \N__34387\ : std_logic;
signal \N__34386\ : std_logic;
signal \N__34385\ : std_logic;
signal \N__34384\ : std_logic;
signal \N__34381\ : std_logic;
signal \N__34376\ : std_logic;
signal \N__34375\ : std_logic;
signal \N__34374\ : std_logic;
signal \N__34373\ : std_logic;
signal \N__34372\ : std_logic;
signal \N__34371\ : std_logic;
signal \N__34370\ : std_logic;
signal \N__34369\ : std_logic;
signal \N__34368\ : std_logic;
signal \N__34367\ : std_logic;
signal \N__34366\ : std_logic;
signal \N__34365\ : std_logic;
signal \N__34364\ : std_logic;
signal \N__34363\ : std_logic;
signal \N__34362\ : std_logic;
signal \N__34361\ : std_logic;
signal \N__34360\ : std_logic;
signal \N__34357\ : std_logic;
signal \N__34356\ : std_logic;
signal \N__34355\ : std_logic;
signal \N__34350\ : std_logic;
signal \N__34347\ : std_logic;
signal \N__34336\ : std_logic;
signal \N__34333\ : std_logic;
signal \N__34330\ : std_logic;
signal \N__34317\ : std_logic;
signal \N__34314\ : std_logic;
signal \N__34311\ : std_logic;
signal \N__34308\ : std_logic;
signal \N__34307\ : std_logic;
signal \N__34306\ : std_logic;
signal \N__34305\ : std_logic;
signal \N__34304\ : std_logic;
signal \N__34303\ : std_logic;
signal \N__34302\ : std_logic;
signal \N__34301\ : std_logic;
signal \N__34300\ : std_logic;
signal \N__34299\ : std_logic;
signal \N__34296\ : std_logic;
signal \N__34295\ : std_logic;
signal \N__34294\ : std_logic;
signal \N__34293\ : std_logic;
signal \N__34292\ : std_logic;
signal \N__34291\ : std_logic;
signal \N__34290\ : std_logic;
signal \N__34289\ : std_logic;
signal \N__34286\ : std_logic;
signal \N__34281\ : std_logic;
signal \N__34276\ : std_logic;
signal \N__34273\ : std_logic;
signal \N__34268\ : std_logic;
signal \N__34263\ : std_logic;
signal \N__34262\ : std_logic;
signal \N__34261\ : std_logic;
signal \N__34260\ : std_logic;
signal \N__34259\ : std_logic;
signal \N__34258\ : std_logic;
signal \N__34257\ : std_logic;
signal \N__34256\ : std_logic;
signal \N__34255\ : std_logic;
signal \N__34252\ : std_logic;
signal \N__34239\ : std_logic;
signal \N__34236\ : std_logic;
signal \N__34233\ : std_logic;
signal \N__34224\ : std_logic;
signal \N__34215\ : std_logic;
signal \N__34210\ : std_logic;
signal \N__34201\ : std_logic;
signal \N__34184\ : std_logic;
signal \N__34181\ : std_logic;
signal \N__34162\ : std_logic;
signal \N__34159\ : std_logic;
signal \N__34158\ : std_logic;
signal \N__34157\ : std_logic;
signal \N__34156\ : std_logic;
signal \N__34155\ : std_logic;
signal \N__34154\ : std_logic;
signal \N__34153\ : std_logic;
signal \N__34152\ : std_logic;
signal \N__34151\ : std_logic;
signal \N__34150\ : std_logic;
signal \N__34149\ : std_logic;
signal \N__34148\ : std_logic;
signal \N__34147\ : std_logic;
signal \N__34142\ : std_logic;
signal \N__34141\ : std_logic;
signal \N__34136\ : std_logic;
signal \N__34133\ : std_logic;
signal \N__34128\ : std_logic;
signal \N__34123\ : std_logic;
signal \N__34122\ : std_logic;
signal \N__34121\ : std_logic;
signal \N__34120\ : std_logic;
signal \N__34115\ : std_logic;
signal \N__34114\ : std_logic;
signal \N__34113\ : std_logic;
signal \N__34112\ : std_logic;
signal \N__34109\ : std_logic;
signal \N__34106\ : std_logic;
signal \N__34103\ : std_logic;
signal \N__34100\ : std_logic;
signal \N__34097\ : std_logic;
signal \N__34096\ : std_logic;
signal \N__34095\ : std_logic;
signal \N__34094\ : std_logic;
signal \N__34089\ : std_logic;
signal \N__34086\ : std_logic;
signal \N__34083\ : std_logic;
signal \N__34080\ : std_logic;
signal \N__34077\ : std_logic;
signal \N__34074\ : std_logic;
signal \N__34071\ : std_logic;
signal \N__34066\ : std_logic;
signal \N__34063\ : std_logic;
signal \N__34060\ : std_logic;
signal \N__34057\ : std_logic;
signal \N__34052\ : std_logic;
signal \N__34045\ : std_logic;
signal \N__34042\ : std_logic;
signal \N__34037\ : std_logic;
signal \N__34012\ : std_logic;
signal \N__34009\ : std_logic;
signal \N__34006\ : std_logic;
signal \N__34003\ : std_logic;
signal \N__34000\ : std_logic;
signal \N__33997\ : std_logic;
signal \N__33994\ : std_logic;
signal \N__33991\ : std_logic;
signal \N__33988\ : std_logic;
signal \N__33985\ : std_logic;
signal \N__33982\ : std_logic;
signal \N__33979\ : std_logic;
signal \N__33976\ : std_logic;
signal \N__33973\ : std_logic;
signal \N__33970\ : std_logic;
signal \N__33967\ : std_logic;
signal \N__33964\ : std_logic;
signal \N__33961\ : std_logic;
signal \N__33960\ : std_logic;
signal \N__33957\ : std_logic;
signal \N__33954\ : std_logic;
signal \N__33951\ : std_logic;
signal \N__33948\ : std_logic;
signal \N__33945\ : std_logic;
signal \N__33940\ : std_logic;
signal \N__33937\ : std_logic;
signal \N__33936\ : std_logic;
signal \N__33933\ : std_logic;
signal \N__33930\ : std_logic;
signal \N__33927\ : std_logic;
signal \N__33924\ : std_logic;
signal \N__33923\ : std_logic;
signal \N__33918\ : std_logic;
signal \N__33915\ : std_logic;
signal \N__33914\ : std_logic;
signal \N__33911\ : std_logic;
signal \N__33908\ : std_logic;
signal \N__33905\ : std_logic;
signal \N__33898\ : std_logic;
signal \N__33895\ : std_logic;
signal \N__33894\ : std_logic;
signal \N__33891\ : std_logic;
signal \N__33888\ : std_logic;
signal \N__33885\ : std_logic;
signal \N__33882\ : std_logic;
signal \N__33877\ : std_logic;
signal \N__33874\ : std_logic;
signal \N__33871\ : std_logic;
signal \N__33868\ : std_logic;
signal \N__33865\ : std_logic;
signal \N__33864\ : std_logic;
signal \N__33861\ : std_logic;
signal \N__33858\ : std_logic;
signal \N__33857\ : std_logic;
signal \N__33854\ : std_logic;
signal \N__33851\ : std_logic;
signal \N__33848\ : std_logic;
signal \N__33843\ : std_logic;
signal \N__33838\ : std_logic;
signal \N__33835\ : std_logic;
signal \N__33832\ : std_logic;
signal \N__33829\ : std_logic;
signal \N__33826\ : std_logic;
signal \N__33823\ : std_logic;
signal \N__33820\ : std_logic;
signal \N__33819\ : std_logic;
signal \N__33818\ : std_logic;
signal \N__33815\ : std_logic;
signal \N__33812\ : std_logic;
signal \N__33809\ : std_logic;
signal \N__33802\ : std_logic;
signal \N__33799\ : std_logic;
signal \N__33796\ : std_logic;
signal \N__33793\ : std_logic;
signal \N__33790\ : std_logic;
signal \N__33787\ : std_logic;
signal \N__33784\ : std_logic;
signal \N__33781\ : std_logic;
signal \N__33780\ : std_logic;
signal \N__33777\ : std_logic;
signal \N__33774\ : std_logic;
signal \N__33769\ : std_logic;
signal \N__33766\ : std_logic;
signal \N__33763\ : std_logic;
signal \N__33760\ : std_logic;
signal \N__33757\ : std_logic;
signal \N__33754\ : std_logic;
signal \N__33753\ : std_logic;
signal \N__33750\ : std_logic;
signal \N__33747\ : std_logic;
signal \N__33744\ : std_logic;
signal \N__33739\ : std_logic;
signal \N__33736\ : std_logic;
signal \N__33733\ : std_logic;
signal \N__33730\ : std_logic;
signal \N__33729\ : std_logic;
signal \N__33726\ : std_logic;
signal \N__33723\ : std_logic;
signal \N__33720\ : std_logic;
signal \N__33715\ : std_logic;
signal \N__33712\ : std_logic;
signal \N__33709\ : std_logic;
signal \N__33706\ : std_logic;
signal \N__33703\ : std_logic;
signal \N__33700\ : std_logic;
signal \N__33697\ : std_logic;
signal \N__33696\ : std_logic;
signal \N__33693\ : std_logic;
signal \N__33690\ : std_logic;
signal \N__33687\ : std_logic;
signal \N__33682\ : std_logic;
signal \N__33679\ : std_logic;
signal \N__33676\ : std_logic;
signal \N__33675\ : std_logic;
signal \N__33672\ : std_logic;
signal \N__33669\ : std_logic;
signal \N__33666\ : std_logic;
signal \N__33661\ : std_logic;
signal \N__33658\ : std_logic;
signal \N__33655\ : std_logic;
signal \N__33654\ : std_logic;
signal \N__33651\ : std_logic;
signal \N__33648\ : std_logic;
signal \N__33645\ : std_logic;
signal \N__33640\ : std_logic;
signal \N__33637\ : std_logic;
signal \N__33634\ : std_logic;
signal \N__33631\ : std_logic;
signal \N__33630\ : std_logic;
signal \N__33627\ : std_logic;
signal \N__33624\ : std_logic;
signal \N__33621\ : std_logic;
signal \N__33616\ : std_logic;
signal \N__33613\ : std_logic;
signal \N__33610\ : std_logic;
signal \N__33607\ : std_logic;
signal \N__33606\ : std_logic;
signal \N__33603\ : std_logic;
signal \N__33600\ : std_logic;
signal \N__33597\ : std_logic;
signal \N__33592\ : std_logic;
signal \N__33589\ : std_logic;
signal \N__33586\ : std_logic;
signal \N__33583\ : std_logic;
signal \N__33580\ : std_logic;
signal \N__33577\ : std_logic;
signal \N__33574\ : std_logic;
signal \N__33571\ : std_logic;
signal \N__33568\ : std_logic;
signal \N__33565\ : std_logic;
signal \N__33562\ : std_logic;
signal \N__33559\ : std_logic;
signal \N__33558\ : std_logic;
signal \N__33555\ : std_logic;
signal \N__33552\ : std_logic;
signal \N__33549\ : std_logic;
signal \N__33546\ : std_logic;
signal \N__33541\ : std_logic;
signal \N__33538\ : std_logic;
signal \N__33535\ : std_logic;
signal \N__33534\ : std_logic;
signal \N__33533\ : std_logic;
signal \N__33530\ : std_logic;
signal \N__33527\ : std_logic;
signal \N__33524\ : std_logic;
signal \N__33521\ : std_logic;
signal \N__33514\ : std_logic;
signal \N__33511\ : std_logic;
signal \N__33508\ : std_logic;
signal \N__33505\ : std_logic;
signal \N__33502\ : std_logic;
signal \N__33499\ : std_logic;
signal \N__33496\ : std_logic;
signal \N__33493\ : std_logic;
signal \N__33492\ : std_logic;
signal \N__33489\ : std_logic;
signal \N__33486\ : std_logic;
signal \N__33481\ : std_logic;
signal \N__33478\ : std_logic;
signal \N__33475\ : std_logic;
signal \N__33472\ : std_logic;
signal \N__33469\ : std_logic;
signal \N__33466\ : std_logic;
signal \N__33463\ : std_logic;
signal \N__33462\ : std_logic;
signal \N__33461\ : std_logic;
signal \N__33458\ : std_logic;
signal \N__33455\ : std_logic;
signal \N__33452\ : std_logic;
signal \N__33449\ : std_logic;
signal \N__33442\ : std_logic;
signal \N__33439\ : std_logic;
signal \N__33438\ : std_logic;
signal \N__33435\ : std_logic;
signal \N__33432\ : std_logic;
signal \N__33429\ : std_logic;
signal \N__33426\ : std_logic;
signal \N__33421\ : std_logic;
signal \N__33418\ : std_logic;
signal \N__33415\ : std_logic;
signal \N__33412\ : std_logic;
signal \N__33409\ : std_logic;
signal \N__33406\ : std_logic;
signal \N__33403\ : std_logic;
signal \N__33400\ : std_logic;
signal \N__33397\ : std_logic;
signal \N__33394\ : std_logic;
signal \N__33391\ : std_logic;
signal \N__33390\ : std_logic;
signal \N__33387\ : std_logic;
signal \N__33384\ : std_logic;
signal \N__33381\ : std_logic;
signal \N__33376\ : std_logic;
signal \N__33373\ : std_logic;
signal \N__33370\ : std_logic;
signal \N__33367\ : std_logic;
signal \N__33364\ : std_logic;
signal \N__33361\ : std_logic;
signal \N__33358\ : std_logic;
signal \N__33355\ : std_logic;
signal \N__33354\ : std_logic;
signal \N__33353\ : std_logic;
signal \N__33350\ : std_logic;
signal \N__33345\ : std_logic;
signal \N__33340\ : std_logic;
signal \N__33337\ : std_logic;
signal \N__33336\ : std_logic;
signal \N__33333\ : std_logic;
signal \N__33330\ : std_logic;
signal \N__33325\ : std_logic;
signal \N__33322\ : std_logic;
signal \N__33319\ : std_logic;
signal \N__33316\ : std_logic;
signal \N__33313\ : std_logic;
signal \N__33310\ : std_logic;
signal \N__33307\ : std_logic;
signal \N__33304\ : std_logic;
signal \N__33301\ : std_logic;
signal \N__33298\ : std_logic;
signal \N__33295\ : std_logic;
signal \N__33292\ : std_logic;
signal \N__33289\ : std_logic;
signal \N__33286\ : std_logic;
signal \N__33283\ : std_logic;
signal \N__33280\ : std_logic;
signal \N__33277\ : std_logic;
signal \N__33274\ : std_logic;
signal \N__33271\ : std_logic;
signal \N__33268\ : std_logic;
signal \N__33265\ : std_logic;
signal \N__33262\ : std_logic;
signal \N__33261\ : std_logic;
signal \N__33258\ : std_logic;
signal \N__33255\ : std_logic;
signal \N__33252\ : std_logic;
signal \N__33249\ : std_logic;
signal \N__33244\ : std_logic;
signal \N__33241\ : std_logic;
signal \N__33238\ : std_logic;
signal \N__33235\ : std_logic;
signal \N__33232\ : std_logic;
signal \N__33229\ : std_logic;
signal \N__33226\ : std_logic;
signal \N__33223\ : std_logic;
signal \N__33220\ : std_logic;
signal \N__33217\ : std_logic;
signal \N__33214\ : std_logic;
signal \N__33211\ : std_logic;
signal \N__33208\ : std_logic;
signal \N__33207\ : std_logic;
signal \N__33204\ : std_logic;
signal \N__33201\ : std_logic;
signal \N__33198\ : std_logic;
signal \N__33195\ : std_logic;
signal \N__33190\ : std_logic;
signal \N__33187\ : std_logic;
signal \N__33184\ : std_logic;
signal \N__33181\ : std_logic;
signal \N__33178\ : std_logic;
signal \N__33175\ : std_logic;
signal \N__33172\ : std_logic;
signal \N__33169\ : std_logic;
signal \N__33166\ : std_logic;
signal \N__33163\ : std_logic;
signal \N__33162\ : std_logic;
signal \N__33159\ : std_logic;
signal \N__33156\ : std_logic;
signal \N__33151\ : std_logic;
signal \N__33148\ : std_logic;
signal \N__33145\ : std_logic;
signal \N__33142\ : std_logic;
signal \N__33139\ : std_logic;
signal \N__33136\ : std_logic;
signal \N__33133\ : std_logic;
signal \N__33130\ : std_logic;
signal \N__33127\ : std_logic;
signal \N__33124\ : std_logic;
signal \N__33121\ : std_logic;
signal \N__33118\ : std_logic;
signal \N__33115\ : std_logic;
signal \N__33112\ : std_logic;
signal \N__33109\ : std_logic;
signal \N__33106\ : std_logic;
signal \N__33103\ : std_logic;
signal \N__33100\ : std_logic;
signal \N__33097\ : std_logic;
signal \N__33094\ : std_logic;
signal \N__33091\ : std_logic;
signal \N__33088\ : std_logic;
signal \N__33085\ : std_logic;
signal \N__33082\ : std_logic;
signal \N__33079\ : std_logic;
signal \N__33076\ : std_logic;
signal \N__33075\ : std_logic;
signal \N__33072\ : std_logic;
signal \N__33069\ : std_logic;
signal \N__33066\ : std_logic;
signal \N__33061\ : std_logic;
signal \N__33058\ : std_logic;
signal \N__33055\ : std_logic;
signal \N__33052\ : std_logic;
signal \N__33049\ : std_logic;
signal \N__33046\ : std_logic;
signal \N__33043\ : std_logic;
signal \N__33040\ : std_logic;
signal \N__33037\ : std_logic;
signal \N__33034\ : std_logic;
signal \N__33033\ : std_logic;
signal \N__33032\ : std_logic;
signal \N__33031\ : std_logic;
signal \N__33024\ : std_logic;
signal \N__33021\ : std_logic;
signal \N__33016\ : std_logic;
signal \N__33015\ : std_logic;
signal \N__33012\ : std_logic;
signal \N__33011\ : std_logic;
signal \N__33010\ : std_logic;
signal \N__33009\ : std_logic;
signal \N__33006\ : std_logic;
signal \N__32997\ : std_logic;
signal \N__32994\ : std_logic;
signal \N__32989\ : std_logic;
signal \N__32988\ : std_logic;
signal \N__32987\ : std_logic;
signal \N__32984\ : std_logic;
signal \N__32979\ : std_logic;
signal \N__32976\ : std_logic;
signal \N__32971\ : std_logic;
signal \N__32968\ : std_logic;
signal \N__32965\ : std_logic;
signal \N__32962\ : std_logic;
signal \N__32959\ : std_logic;
signal \N__32956\ : std_logic;
signal \N__32953\ : std_logic;
signal \N__32952\ : std_logic;
signal \N__32951\ : std_logic;
signal \N__32948\ : std_logic;
signal \N__32943\ : std_logic;
signal \N__32938\ : std_logic;
signal \N__32935\ : std_logic;
signal \N__32932\ : std_logic;
signal \N__32931\ : std_logic;
signal \N__32930\ : std_logic;
signal \N__32927\ : std_logic;
signal \N__32924\ : std_logic;
signal \N__32921\ : std_logic;
signal \N__32914\ : std_logic;
signal \N__32913\ : std_logic;
signal \N__32912\ : std_logic;
signal \N__32909\ : std_logic;
signal \N__32908\ : std_logic;
signal \N__32905\ : std_logic;
signal \N__32904\ : std_logic;
signal \N__32903\ : std_logic;
signal \N__32900\ : std_logic;
signal \N__32897\ : std_logic;
signal \N__32896\ : std_logic;
signal \N__32895\ : std_logic;
signal \N__32894\ : std_logic;
signal \N__32893\ : std_logic;
signal \N__32890\ : std_logic;
signal \N__32887\ : std_logic;
signal \N__32886\ : std_logic;
signal \N__32885\ : std_logic;
signal \N__32884\ : std_logic;
signal \N__32881\ : std_logic;
signal \N__32880\ : std_logic;
signal \N__32877\ : std_logic;
signal \N__32874\ : std_logic;
signal \N__32873\ : std_logic;
signal \N__32872\ : std_logic;
signal \N__32871\ : std_logic;
signal \N__32868\ : std_logic;
signal \N__32865\ : std_logic;
signal \N__32862\ : std_logic;
signal \N__32861\ : std_logic;
signal \N__32858\ : std_logic;
signal \N__32855\ : std_logic;
signal \N__32850\ : std_logic;
signal \N__32847\ : std_logic;
signal \N__32846\ : std_logic;
signal \N__32843\ : std_logic;
signal \N__32842\ : std_logic;
signal \N__32839\ : std_logic;
signal \N__32836\ : std_logic;
signal \N__32833\ : std_logic;
signal \N__32830\ : std_logic;
signal \N__32827\ : std_logic;
signal \N__32824\ : std_logic;
signal \N__32821\ : std_logic;
signal \N__32818\ : std_logic;
signal \N__32815\ : std_logic;
signal \N__32810\ : std_logic;
signal \N__32807\ : std_logic;
signal \N__32806\ : std_logic;
signal \N__32801\ : std_logic;
signal \N__32796\ : std_logic;
signal \N__32793\ : std_logic;
signal \N__32790\ : std_logic;
signal \N__32787\ : std_logic;
signal \N__32784\ : std_logic;
signal \N__32779\ : std_logic;
signal \N__32778\ : std_logic;
signal \N__32775\ : std_logic;
signal \N__32770\ : std_logic;
signal \N__32765\ : std_logic;
signal \N__32762\ : std_logic;
signal \N__32757\ : std_logic;
signal \N__32754\ : std_logic;
signal \N__32751\ : std_logic;
signal \N__32746\ : std_logic;
signal \N__32741\ : std_logic;
signal \N__32736\ : std_logic;
signal \N__32733\ : std_logic;
signal \N__32728\ : std_logic;
signal \N__32727\ : std_logic;
signal \N__32724\ : std_logic;
signal \N__32719\ : std_logic;
signal \N__32716\ : std_logic;
signal \N__32711\ : std_logic;
signal \N__32704\ : std_logic;
signal \N__32701\ : std_logic;
signal \N__32698\ : std_logic;
signal \N__32693\ : std_logic;
signal \N__32688\ : std_logic;
signal \N__32685\ : std_logic;
signal \N__32680\ : std_logic;
signal \N__32671\ : std_logic;
signal \N__32668\ : std_logic;
signal \N__32665\ : std_logic;
signal \N__32662\ : std_logic;
signal \N__32659\ : std_logic;
signal \N__32656\ : std_logic;
signal \N__32653\ : std_logic;
signal \N__32650\ : std_logic;
signal \N__32647\ : std_logic;
signal \N__32644\ : std_logic;
signal \N__32641\ : std_logic;
signal \N__32640\ : std_logic;
signal \N__32637\ : std_logic;
signal \N__32634\ : std_logic;
signal \N__32633\ : std_logic;
signal \N__32632\ : std_logic;
signal \N__32629\ : std_logic;
signal \N__32626\ : std_logic;
signal \N__32625\ : std_logic;
signal \N__32622\ : std_logic;
signal \N__32619\ : std_logic;
signal \N__32616\ : std_logic;
signal \N__32613\ : std_logic;
signal \N__32610\ : std_logic;
signal \N__32599\ : std_logic;
signal \N__32596\ : std_logic;
signal \N__32595\ : std_logic;
signal \N__32592\ : std_logic;
signal \N__32591\ : std_logic;
signal \N__32590\ : std_logic;
signal \N__32589\ : std_logic;
signal \N__32586\ : std_logic;
signal \N__32583\ : std_logic;
signal \N__32580\ : std_logic;
signal \N__32575\ : std_logic;
signal \N__32566\ : std_logic;
signal \N__32563\ : std_logic;
signal \N__32560\ : std_logic;
signal \N__32557\ : std_logic;
signal \N__32554\ : std_logic;
signal \N__32551\ : std_logic;
signal \N__32548\ : std_logic;
signal \N__32547\ : std_logic;
signal \N__32546\ : std_logic;
signal \N__32543\ : std_logic;
signal \N__32542\ : std_logic;
signal \N__32541\ : std_logic;
signal \N__32538\ : std_logic;
signal \N__32535\ : std_logic;
signal \N__32532\ : std_logic;
signal \N__32527\ : std_logic;
signal \N__32518\ : std_logic;
signal \N__32515\ : std_logic;
signal \N__32512\ : std_logic;
signal \N__32511\ : std_logic;
signal \N__32510\ : std_logic;
signal \N__32509\ : std_logic;
signal \N__32506\ : std_logic;
signal \N__32505\ : std_logic;
signal \N__32502\ : std_logic;
signal \N__32499\ : std_logic;
signal \N__32496\ : std_logic;
signal \N__32493\ : std_logic;
signal \N__32488\ : std_logic;
signal \N__32479\ : std_logic;
signal \N__32476\ : std_logic;
signal \N__32473\ : std_logic;
signal \N__32470\ : std_logic;
signal \N__32467\ : std_logic;
signal \N__32466\ : std_logic;
signal \N__32465\ : std_logic;
signal \N__32464\ : std_logic;
signal \N__32463\ : std_logic;
signal \N__32460\ : std_logic;
signal \N__32457\ : std_logic;
signal \N__32450\ : std_logic;
signal \N__32447\ : std_logic;
signal \N__32440\ : std_logic;
signal \N__32437\ : std_logic;
signal \N__32436\ : std_logic;
signal \N__32435\ : std_logic;
signal \N__32432\ : std_logic;
signal \N__32429\ : std_logic;
signal \N__32426\ : std_logic;
signal \N__32419\ : std_logic;
signal \N__32416\ : std_logic;
signal \N__32413\ : std_logic;
signal \N__32410\ : std_logic;
signal \N__32409\ : std_logic;
signal \N__32404\ : std_logic;
signal \N__32401\ : std_logic;
signal \N__32398\ : std_logic;
signal \N__32395\ : std_logic;
signal \N__32392\ : std_logic;
signal \N__32389\ : std_logic;
signal \N__32386\ : std_logic;
signal \N__32383\ : std_logic;
signal \N__32382\ : std_logic;
signal \N__32379\ : std_logic;
signal \N__32376\ : std_logic;
signal \N__32371\ : std_logic;
signal \N__32370\ : std_logic;
signal \N__32367\ : std_logic;
signal \N__32366\ : std_logic;
signal \N__32363\ : std_logic;
signal \N__32360\ : std_logic;
signal \N__32355\ : std_logic;
signal \N__32350\ : std_logic;
signal \N__32347\ : std_logic;
signal \N__32344\ : std_logic;
signal \N__32341\ : std_logic;
signal \N__32338\ : std_logic;
signal \N__32337\ : std_logic;
signal \N__32336\ : std_logic;
signal \N__32333\ : std_logic;
signal \N__32330\ : std_logic;
signal \N__32327\ : std_logic;
signal \N__32320\ : std_logic;
signal \N__32317\ : std_logic;
signal \N__32314\ : std_logic;
signal \N__32311\ : std_logic;
signal \N__32310\ : std_logic;
signal \N__32307\ : std_logic;
signal \N__32304\ : std_logic;
signal \N__32301\ : std_logic;
signal \N__32300\ : std_logic;
signal \N__32297\ : std_logic;
signal \N__32294\ : std_logic;
signal \N__32291\ : std_logic;
signal \N__32288\ : std_logic;
signal \N__32281\ : std_logic;
signal \N__32278\ : std_logic;
signal \N__32275\ : std_logic;
signal \N__32272\ : std_logic;
signal \N__32271\ : std_logic;
signal \N__32268\ : std_logic;
signal \N__32265\ : std_logic;
signal \N__32262\ : std_logic;
signal \N__32259\ : std_logic;
signal \N__32258\ : std_logic;
signal \N__32255\ : std_logic;
signal \N__32252\ : std_logic;
signal \N__32249\ : std_logic;
signal \N__32246\ : std_logic;
signal \N__32239\ : std_logic;
signal \N__32238\ : std_logic;
signal \N__32235\ : std_logic;
signal \N__32232\ : std_logic;
signal \N__32231\ : std_logic;
signal \N__32228\ : std_logic;
signal \N__32225\ : std_logic;
signal \N__32222\ : std_logic;
signal \N__32219\ : std_logic;
signal \N__32212\ : std_logic;
signal \N__32209\ : std_logic;
signal \N__32206\ : std_logic;
signal \N__32203\ : std_logic;
signal \N__32200\ : std_logic;
signal \N__32197\ : std_logic;
signal \N__32194\ : std_logic;
signal \N__32191\ : std_logic;
signal \N__32188\ : std_logic;
signal \N__32185\ : std_logic;
signal \N__32182\ : std_logic;
signal \N__32181\ : std_logic;
signal \N__32180\ : std_logic;
signal \N__32179\ : std_logic;
signal \N__32178\ : std_logic;
signal \N__32173\ : std_logic;
signal \N__32170\ : std_logic;
signal \N__32165\ : std_logic;
signal \N__32164\ : std_logic;
signal \N__32163\ : std_logic;
signal \N__32162\ : std_logic;
signal \N__32161\ : std_logic;
signal \N__32160\ : std_logic;
signal \N__32159\ : std_logic;
signal \N__32158\ : std_logic;
signal \N__32157\ : std_logic;
signal \N__32156\ : std_logic;
signal \N__32155\ : std_logic;
signal \N__32152\ : std_logic;
signal \N__32147\ : std_logic;
signal \N__32138\ : std_logic;
signal \N__32131\ : std_logic;
signal \N__32128\ : std_logic;
signal \N__32125\ : std_logic;
signal \N__32122\ : std_logic;
signal \N__32117\ : std_logic;
signal \N__32108\ : std_logic;
signal \N__32101\ : std_logic;
signal \N__32100\ : std_logic;
signal \N__32099\ : std_logic;
signal \N__32096\ : std_logic;
signal \N__32095\ : std_logic;
signal \N__32094\ : std_logic;
signal \N__32091\ : std_logic;
signal \N__32088\ : std_logic;
signal \N__32087\ : std_logic;
signal \N__32084\ : std_logic;
signal \N__32079\ : std_logic;
signal \N__32074\ : std_logic;
signal \N__32071\ : std_logic;
signal \N__32070\ : std_logic;
signal \N__32069\ : std_logic;
signal \N__32068\ : std_logic;
signal \N__32067\ : std_logic;
signal \N__32064\ : std_logic;
signal \N__32061\ : std_logic;
signal \N__32058\ : std_logic;
signal \N__32055\ : std_logic;
signal \N__32052\ : std_logic;
signal \N__32045\ : std_logic;
signal \N__32032\ : std_logic;
signal \N__32029\ : std_logic;
signal \N__32026\ : std_logic;
signal \N__32023\ : std_logic;
signal \N__32020\ : std_logic;
signal \N__32017\ : std_logic;
signal \N__32016\ : std_logic;
signal \N__32013\ : std_logic;
signal \N__32012\ : std_logic;
signal \N__32009\ : std_logic;
signal \N__32006\ : std_logic;
signal \N__32003\ : std_logic;
signal \N__31998\ : std_logic;
signal \N__31995\ : std_logic;
signal \N__31990\ : std_logic;
signal \N__31987\ : std_logic;
signal \N__31986\ : std_logic;
signal \N__31983\ : std_logic;
signal \N__31980\ : std_logic;
signal \N__31979\ : std_logic;
signal \N__31976\ : std_logic;
signal \N__31973\ : std_logic;
signal \N__31970\ : std_logic;
signal \N__31965\ : std_logic;
signal \N__31960\ : std_logic;
signal \N__31957\ : std_logic;
signal \N__31954\ : std_logic;
signal \N__31951\ : std_logic;
signal \N__31948\ : std_logic;
signal \N__31945\ : std_logic;
signal \N__31942\ : std_logic;
signal \N__31939\ : std_logic;
signal \N__31936\ : std_logic;
signal \N__31933\ : std_logic;
signal \N__31932\ : std_logic;
signal \N__31931\ : std_logic;
signal \N__31928\ : std_logic;
signal \N__31925\ : std_logic;
signal \N__31922\ : std_logic;
signal \N__31917\ : std_logic;
signal \N__31914\ : std_logic;
signal \N__31911\ : std_logic;
signal \N__31906\ : std_logic;
signal \N__31905\ : std_logic;
signal \N__31904\ : std_logic;
signal \N__31899\ : std_logic;
signal \N__31896\ : std_logic;
signal \N__31891\ : std_logic;
signal \N__31888\ : std_logic;
signal \N__31885\ : std_logic;
signal \N__31884\ : std_logic;
signal \N__31883\ : std_logic;
signal \N__31882\ : std_logic;
signal \N__31879\ : std_logic;
signal \N__31876\ : std_logic;
signal \N__31873\ : std_logic;
signal \N__31870\ : std_logic;
signal \N__31861\ : std_logic;
signal \N__31860\ : std_logic;
signal \N__31859\ : std_logic;
signal \N__31858\ : std_logic;
signal \N__31855\ : std_logic;
signal \N__31852\ : std_logic;
signal \N__31847\ : std_logic;
signal \N__31840\ : std_logic;
signal \N__31837\ : std_logic;
signal \N__31834\ : std_logic;
signal \N__31831\ : std_logic;
signal \N__31828\ : std_logic;
signal \N__31827\ : std_logic;
signal \N__31824\ : std_logic;
signal \N__31821\ : std_logic;
signal \N__31820\ : std_logic;
signal \N__31815\ : std_logic;
signal \N__31812\ : std_logic;
signal \N__31809\ : std_logic;
signal \N__31804\ : std_logic;
signal \N__31801\ : std_logic;
signal \N__31798\ : std_logic;
signal \N__31795\ : std_logic;
signal \N__31792\ : std_logic;
signal \N__31789\ : std_logic;
signal \N__31786\ : std_logic;
signal \N__31783\ : std_logic;
signal \N__31780\ : std_logic;
signal \N__31777\ : std_logic;
signal \N__31776\ : std_logic;
signal \N__31773\ : std_logic;
signal \N__31770\ : std_logic;
signal \N__31769\ : std_logic;
signal \N__31768\ : std_logic;
signal \N__31767\ : std_logic;
signal \N__31766\ : std_logic;
signal \N__31763\ : std_logic;
signal \N__31760\ : std_logic;
signal \N__31757\ : std_logic;
signal \N__31754\ : std_logic;
signal \N__31753\ : std_logic;
signal \N__31752\ : std_logic;
signal \N__31751\ : std_logic;
signal \N__31750\ : std_logic;
signal \N__31747\ : std_logic;
signal \N__31744\ : std_logic;
signal \N__31741\ : std_logic;
signal \N__31736\ : std_logic;
signal \N__31733\ : std_logic;
signal \N__31730\ : std_logic;
signal \N__31727\ : std_logic;
signal \N__31726\ : std_logic;
signal \N__31723\ : std_logic;
signal \N__31720\ : std_logic;
signal \N__31719\ : std_logic;
signal \N__31716\ : std_logic;
signal \N__31713\ : std_logic;
signal \N__31708\ : std_logic;
signal \N__31703\ : std_logic;
signal \N__31700\ : std_logic;
signal \N__31697\ : std_logic;
signal \N__31694\ : std_logic;
signal \N__31691\ : std_logic;
signal \N__31688\ : std_logic;
signal \N__31685\ : std_logic;
signal \N__31682\ : std_logic;
signal \N__31677\ : std_logic;
signal \N__31672\ : std_logic;
signal \N__31665\ : std_logic;
signal \N__31662\ : std_logic;
signal \N__31659\ : std_logic;
signal \N__31654\ : std_logic;
signal \N__31651\ : std_logic;
signal \N__31648\ : std_logic;
signal \N__31641\ : std_logic;
signal \N__31636\ : std_logic;
signal \N__31633\ : std_logic;
signal \N__31630\ : std_logic;
signal \N__31627\ : std_logic;
signal \N__31624\ : std_logic;
signal \N__31621\ : std_logic;
signal \N__31618\ : std_logic;
signal \N__31615\ : std_logic;
signal \N__31612\ : std_logic;
signal \N__31609\ : std_logic;
signal \N__31606\ : std_logic;
signal \N__31603\ : std_logic;
signal \N__31600\ : std_logic;
signal \N__31597\ : std_logic;
signal \N__31594\ : std_logic;
signal \N__31591\ : std_logic;
signal \N__31588\ : std_logic;
signal \N__31587\ : std_logic;
signal \N__31584\ : std_logic;
signal \N__31581\ : std_logic;
signal \N__31578\ : std_logic;
signal \N__31575\ : std_logic;
signal \N__31572\ : std_logic;
signal \N__31569\ : std_logic;
signal \N__31566\ : std_logic;
signal \N__31563\ : std_logic;
signal \N__31560\ : std_logic;
signal \N__31557\ : std_logic;
signal \N__31554\ : std_logic;
signal \N__31551\ : std_logic;
signal \N__31548\ : std_logic;
signal \N__31545\ : std_logic;
signal \N__31542\ : std_logic;
signal \N__31537\ : std_logic;
signal \N__31534\ : std_logic;
signal \N__31533\ : std_logic;
signal \N__31530\ : std_logic;
signal \N__31529\ : std_logic;
signal \N__31526\ : std_logic;
signal \N__31523\ : std_logic;
signal \N__31520\ : std_logic;
signal \N__31513\ : std_logic;
signal \N__31510\ : std_logic;
signal \N__31507\ : std_logic;
signal \N__31504\ : std_logic;
signal \N__31501\ : std_logic;
signal \N__31498\ : std_logic;
signal \N__31495\ : std_logic;
signal \N__31492\ : std_logic;
signal \N__31489\ : std_logic;
signal \N__31488\ : std_logic;
signal \N__31483\ : std_logic;
signal \N__31480\ : std_logic;
signal \N__31477\ : std_logic;
signal \N__31474\ : std_logic;
signal \N__31471\ : std_logic;
signal \N__31468\ : std_logic;
signal \N__31465\ : std_logic;
signal \N__31462\ : std_logic;
signal \N__31459\ : std_logic;
signal \N__31456\ : std_logic;
signal \N__31453\ : std_logic;
signal \N__31450\ : std_logic;
signal \N__31447\ : std_logic;
signal \N__31444\ : std_logic;
signal \N__31441\ : std_logic;
signal \N__31438\ : std_logic;
signal \N__31435\ : std_logic;
signal \N__31434\ : std_logic;
signal \N__31431\ : std_logic;
signal \N__31428\ : std_logic;
signal \N__31425\ : std_logic;
signal \N__31422\ : std_logic;
signal \N__31419\ : std_logic;
signal \N__31416\ : std_logic;
signal \N__31413\ : std_logic;
signal \N__31410\ : std_logic;
signal \N__31407\ : std_logic;
signal \N__31404\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31398\ : std_logic;
signal \N__31395\ : std_logic;
signal \N__31392\ : std_logic;
signal \N__31389\ : std_logic;
signal \N__31384\ : std_logic;
signal \N__31381\ : std_logic;
signal \N__31378\ : std_logic;
signal \N__31377\ : std_logic;
signal \N__31376\ : std_logic;
signal \N__31373\ : std_logic;
signal \N__31370\ : std_logic;
signal \N__31367\ : std_logic;
signal \N__31364\ : std_logic;
signal \N__31357\ : std_logic;
signal \N__31356\ : std_logic;
signal \N__31353\ : std_logic;
signal \N__31350\ : std_logic;
signal \N__31347\ : std_logic;
signal \N__31342\ : std_logic;
signal \N__31339\ : std_logic;
signal \N__31336\ : std_logic;
signal \N__31333\ : std_logic;
signal \N__31332\ : std_logic;
signal \N__31329\ : std_logic;
signal \N__31326\ : std_logic;
signal \N__31323\ : std_logic;
signal \N__31320\ : std_logic;
signal \N__31317\ : std_logic;
signal \N__31312\ : std_logic;
signal \N__31309\ : std_logic;
signal \N__31306\ : std_logic;
signal \N__31303\ : std_logic;
signal \N__31302\ : std_logic;
signal \N__31299\ : std_logic;
signal \N__31296\ : std_logic;
signal \N__31293\ : std_logic;
signal \N__31288\ : std_logic;
signal \N__31287\ : std_logic;
signal \N__31284\ : std_logic;
signal \N__31281\ : std_logic;
signal \N__31278\ : std_logic;
signal \N__31273\ : std_logic;
signal \N__31270\ : std_logic;
signal \N__31267\ : std_logic;
signal \N__31264\ : std_logic;
signal \N__31261\ : std_logic;
signal \N__31258\ : std_logic;
signal \N__31255\ : std_logic;
signal \N__31252\ : std_logic;
signal \N__31249\ : std_logic;
signal \N__31246\ : std_logic;
signal \N__31243\ : std_logic;
signal \N__31240\ : std_logic;
signal \N__31237\ : std_logic;
signal \N__31234\ : std_logic;
signal \N__31231\ : std_logic;
signal \N__31228\ : std_logic;
signal \N__31225\ : std_logic;
signal \N__31222\ : std_logic;
signal \N__31221\ : std_logic;
signal \N__31218\ : std_logic;
signal \N__31215\ : std_logic;
signal \N__31212\ : std_logic;
signal \N__31207\ : std_logic;
signal \N__31204\ : std_logic;
signal \N__31201\ : std_logic;
signal \N__31198\ : std_logic;
signal \N__31195\ : std_logic;
signal \N__31194\ : std_logic;
signal \N__31191\ : std_logic;
signal \N__31188\ : std_logic;
signal \N__31185\ : std_logic;
signal \N__31180\ : std_logic;
signal \N__31177\ : std_logic;
signal \N__31176\ : std_logic;
signal \N__31173\ : std_logic;
signal \N__31170\ : std_logic;
signal \N__31167\ : std_logic;
signal \N__31164\ : std_logic;
signal \N__31159\ : std_logic;
signal \N__31156\ : std_logic;
signal \N__31153\ : std_logic;
signal \N__31150\ : std_logic;
signal \N__31147\ : std_logic;
signal \N__31146\ : std_logic;
signal \N__31143\ : std_logic;
signal \N__31140\ : std_logic;
signal \N__31137\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31131\ : std_logic;
signal \N__31126\ : std_logic;
signal \N__31123\ : std_logic;
signal \N__31120\ : std_logic;
signal \N__31117\ : std_logic;
signal \N__31114\ : std_logic;
signal \N__31111\ : std_logic;
signal \N__31108\ : std_logic;
signal \N__31105\ : std_logic;
signal \N__31102\ : std_logic;
signal \N__31099\ : std_logic;
signal \N__31096\ : std_logic;
signal \N__31093\ : std_logic;
signal \N__31090\ : std_logic;
signal \N__31087\ : std_logic;
signal \N__31084\ : std_logic;
signal \N__31081\ : std_logic;
signal \N__31078\ : std_logic;
signal \N__31075\ : std_logic;
signal \N__31072\ : std_logic;
signal \N__31069\ : std_logic;
signal \N__31066\ : std_logic;
signal \N__31063\ : std_logic;
signal \N__31060\ : std_logic;
signal \N__31057\ : std_logic;
signal \N__31054\ : std_logic;
signal \N__31051\ : std_logic;
signal \N__31048\ : std_logic;
signal \N__31045\ : std_logic;
signal \N__31042\ : std_logic;
signal \N__31039\ : std_logic;
signal \N__31036\ : std_logic;
signal \N__31033\ : std_logic;
signal \N__31030\ : std_logic;
signal \N__31027\ : std_logic;
signal \N__31024\ : std_logic;
signal \N__31021\ : std_logic;
signal \N__31018\ : std_logic;
signal \N__31015\ : std_logic;
signal \N__31012\ : std_logic;
signal \N__31009\ : std_logic;
signal \N__31006\ : std_logic;
signal \N__31003\ : std_logic;
signal \N__31000\ : std_logic;
signal \N__30999\ : std_logic;
signal \N__30994\ : std_logic;
signal \N__30993\ : std_logic;
signal \N__30992\ : std_logic;
signal \N__30991\ : std_logic;
signal \N__30990\ : std_logic;
signal \N__30989\ : std_logic;
signal \N__30986\ : std_logic;
signal \N__30983\ : std_logic;
signal \N__30980\ : std_logic;
signal \N__30977\ : std_logic;
signal \N__30972\ : std_logic;
signal \N__30969\ : std_logic;
signal \N__30966\ : std_logic;
signal \N__30959\ : std_logic;
signal \N__30956\ : std_logic;
signal \N__30953\ : std_logic;
signal \N__30950\ : std_logic;
signal \N__30943\ : std_logic;
signal \N__30940\ : std_logic;
signal \N__30939\ : std_logic;
signal \N__30936\ : std_logic;
signal \N__30933\ : std_logic;
signal \N__30932\ : std_logic;
signal \N__30931\ : std_logic;
signal \N__30930\ : std_logic;
signal \N__30929\ : std_logic;
signal \N__30928\ : std_logic;
signal \N__30925\ : std_logic;
signal \N__30922\ : std_logic;
signal \N__30917\ : std_logic;
signal \N__30912\ : std_logic;
signal \N__30909\ : std_logic;
signal \N__30898\ : std_logic;
signal \N__30895\ : std_logic;
signal \N__30892\ : std_logic;
signal \N__30889\ : std_logic;
signal \N__30886\ : std_logic;
signal \N__30883\ : std_logic;
signal \N__30880\ : std_logic;
signal \N__30877\ : std_logic;
signal \N__30874\ : std_logic;
signal \N__30871\ : std_logic;
signal \N__30868\ : std_logic;
signal \N__30865\ : std_logic;
signal \N__30862\ : std_logic;
signal \N__30859\ : std_logic;
signal \N__30856\ : std_logic;
signal \N__30853\ : std_logic;
signal \N__30850\ : std_logic;
signal \N__30847\ : std_logic;
signal \N__30844\ : std_logic;
signal \N__30841\ : std_logic;
signal \N__30838\ : std_logic;
signal \N__30835\ : std_logic;
signal \N__30832\ : std_logic;
signal \N__30829\ : std_logic;
signal \N__30826\ : std_logic;
signal \N__30823\ : std_logic;
signal \N__30820\ : std_logic;
signal \N__30817\ : std_logic;
signal \N__30814\ : std_logic;
signal \N__30811\ : std_logic;
signal \N__30810\ : std_logic;
signal \N__30807\ : std_logic;
signal \N__30804\ : std_logic;
signal \N__30803\ : std_logic;
signal \N__30800\ : std_logic;
signal \N__30797\ : std_logic;
signal \N__30794\ : std_logic;
signal \N__30791\ : std_logic;
signal \N__30788\ : std_logic;
signal \N__30785\ : std_logic;
signal \N__30778\ : std_logic;
signal \N__30775\ : std_logic;
signal \N__30772\ : std_logic;
signal \N__30771\ : std_logic;
signal \N__30770\ : std_logic;
signal \N__30767\ : std_logic;
signal \N__30764\ : std_logic;
signal \N__30761\ : std_logic;
signal \N__30754\ : std_logic;
signal \N__30751\ : std_logic;
signal \N__30748\ : std_logic;
signal \N__30745\ : std_logic;
signal \N__30744\ : std_logic;
signal \N__30741\ : std_logic;
signal \N__30740\ : std_logic;
signal \N__30739\ : std_logic;
signal \N__30736\ : std_logic;
signal \N__30729\ : std_logic;
signal \N__30724\ : std_logic;
signal \N__30723\ : std_logic;
signal \N__30722\ : std_logic;
signal \N__30721\ : std_logic;
signal \N__30718\ : std_logic;
signal \N__30711\ : std_logic;
signal \N__30706\ : std_logic;
signal \N__30703\ : std_logic;
signal \N__30702\ : std_logic;
signal \N__30701\ : std_logic;
signal \N__30698\ : std_logic;
signal \N__30693\ : std_logic;
signal \N__30688\ : std_logic;
signal \N__30685\ : std_logic;
signal \N__30682\ : std_logic;
signal \N__30679\ : std_logic;
signal \N__30676\ : std_logic;
signal \N__30673\ : std_logic;
signal \N__30670\ : std_logic;
signal \N__30667\ : std_logic;
signal \N__30664\ : std_logic;
signal \N__30663\ : std_logic;
signal \N__30660\ : std_logic;
signal \N__30657\ : std_logic;
signal \N__30654\ : std_logic;
signal \N__30649\ : std_logic;
signal \N__30646\ : std_logic;
signal \N__30643\ : std_logic;
signal \N__30640\ : std_logic;
signal \N__30637\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30633\ : std_logic;
signal \N__30630\ : std_logic;
signal \N__30625\ : std_logic;
signal \N__30624\ : std_logic;
signal \N__30623\ : std_logic;
signal \N__30616\ : std_logic;
signal \N__30613\ : std_logic;
signal \N__30610\ : std_logic;
signal \N__30607\ : std_logic;
signal \N__30604\ : std_logic;
signal \N__30601\ : std_logic;
signal \N__30598\ : std_logic;
signal \N__30595\ : std_logic;
signal \N__30594\ : std_logic;
signal \N__30591\ : std_logic;
signal \N__30588\ : std_logic;
signal \N__30583\ : std_logic;
signal \N__30580\ : std_logic;
signal \N__30579\ : std_logic;
signal \N__30576\ : std_logic;
signal \N__30573\ : std_logic;
signal \N__30568\ : std_logic;
signal \N__30567\ : std_logic;
signal \N__30564\ : std_logic;
signal \N__30561\ : std_logic;
signal \N__30558\ : std_logic;
signal \N__30553\ : std_logic;
signal \N__30550\ : std_logic;
signal \N__30549\ : std_logic;
signal \N__30546\ : std_logic;
signal \N__30543\ : std_logic;
signal \N__30538\ : std_logic;
signal \N__30535\ : std_logic;
signal \N__30532\ : std_logic;
signal \N__30529\ : std_logic;
signal \N__30528\ : std_logic;
signal \N__30525\ : std_logic;
signal \N__30522\ : std_logic;
signal \N__30519\ : std_logic;
signal \N__30516\ : std_logic;
signal \N__30511\ : std_logic;
signal \N__30508\ : std_logic;
signal \N__30505\ : std_logic;
signal \N__30502\ : std_logic;
signal \N__30499\ : std_logic;
signal \N__30496\ : std_logic;
signal \N__30493\ : std_logic;
signal \N__30490\ : std_logic;
signal \N__30487\ : std_logic;
signal \N__30484\ : std_logic;
signal \N__30481\ : std_logic;
signal \N__30478\ : std_logic;
signal \N__30475\ : std_logic;
signal \N__30472\ : std_logic;
signal \N__30469\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30463\ : std_logic;
signal \N__30462\ : std_logic;
signal \N__30461\ : std_logic;
signal \N__30458\ : std_logic;
signal \N__30455\ : std_logic;
signal \N__30454\ : std_logic;
signal \N__30451\ : std_logic;
signal \N__30448\ : std_logic;
signal \N__30443\ : std_logic;
signal \N__30442\ : std_logic;
signal \N__30439\ : std_logic;
signal \N__30436\ : std_logic;
signal \N__30433\ : std_logic;
signal \N__30430\ : std_logic;
signal \N__30427\ : std_logic;
signal \N__30422\ : std_logic;
signal \N__30415\ : std_logic;
signal \N__30412\ : std_logic;
signal \N__30409\ : std_logic;
signal \N__30406\ : std_logic;
signal \N__30403\ : std_logic;
signal \N__30400\ : std_logic;
signal \N__30397\ : std_logic;
signal \N__30394\ : std_logic;
signal \N__30391\ : std_logic;
signal \N__30390\ : std_logic;
signal \N__30387\ : std_logic;
signal \N__30384\ : std_logic;
signal \N__30379\ : std_logic;
signal \N__30378\ : std_logic;
signal \N__30375\ : std_logic;
signal \N__30372\ : std_logic;
signal \N__30367\ : std_logic;
signal \N__30366\ : std_logic;
signal \N__30363\ : std_logic;
signal \N__30360\ : std_logic;
signal \N__30357\ : std_logic;
signal \N__30354\ : std_logic;
signal \N__30349\ : std_logic;
signal \N__30348\ : std_logic;
signal \N__30345\ : std_logic;
signal \N__30342\ : std_logic;
signal \N__30337\ : std_logic;
signal \N__30334\ : std_logic;
signal \N__30333\ : std_logic;
signal \N__30330\ : std_logic;
signal \N__30327\ : std_logic;
signal \N__30322\ : std_logic;
signal \N__30319\ : std_logic;
signal \N__30318\ : std_logic;
signal \N__30315\ : std_logic;
signal \N__30312\ : std_logic;
signal \N__30307\ : std_logic;
signal \N__30306\ : std_logic;
signal \N__30303\ : std_logic;
signal \N__30300\ : std_logic;
signal \N__30297\ : std_logic;
signal \N__30292\ : std_logic;
signal \N__30291\ : std_logic;
signal \N__30288\ : std_logic;
signal \N__30285\ : std_logic;
signal \N__30280\ : std_logic;
signal \N__30277\ : std_logic;
signal \N__30274\ : std_logic;
signal \N__30271\ : std_logic;
signal \N__30270\ : std_logic;
signal \N__30267\ : std_logic;
signal \N__30264\ : std_logic;
signal \N__30259\ : std_logic;
signal \N__30258\ : std_logic;
signal \N__30255\ : std_logic;
signal \N__30252\ : std_logic;
signal \N__30247\ : std_logic;
signal \N__30246\ : std_logic;
signal \N__30243\ : std_logic;
signal \N__30240\ : std_logic;
signal \N__30237\ : std_logic;
signal \N__30232\ : std_logic;
signal \N__30231\ : std_logic;
signal \N__30228\ : std_logic;
signal \N__30225\ : std_logic;
signal \N__30220\ : std_logic;
signal \N__30217\ : std_logic;
signal \N__30214\ : std_logic;
signal \N__30211\ : std_logic;
signal \N__30208\ : std_logic;
signal \N__30205\ : std_logic;
signal \N__30204\ : std_logic;
signal \N__30203\ : std_logic;
signal \N__30200\ : std_logic;
signal \N__30197\ : std_logic;
signal \N__30194\ : std_logic;
signal \N__30187\ : std_logic;
signal \N__30186\ : std_logic;
signal \N__30185\ : std_logic;
signal \N__30182\ : std_logic;
signal \N__30179\ : std_logic;
signal \N__30176\ : std_logic;
signal \N__30173\ : std_logic;
signal \N__30170\ : std_logic;
signal \N__30163\ : std_logic;
signal \N__30160\ : std_logic;
signal \N__30157\ : std_logic;
signal \N__30154\ : std_logic;
signal \N__30151\ : std_logic;
signal \N__30148\ : std_logic;
signal \N__30145\ : std_logic;
signal \N__30142\ : std_logic;
signal \N__30141\ : std_logic;
signal \N__30140\ : std_logic;
signal \N__30139\ : std_logic;
signal \N__30134\ : std_logic;
signal \N__30133\ : std_logic;
signal \N__30128\ : std_logic;
signal \N__30125\ : std_logic;
signal \N__30122\ : std_logic;
signal \N__30119\ : std_logic;
signal \N__30116\ : std_logic;
signal \N__30111\ : std_logic;
signal \N__30106\ : std_logic;
signal \N__30103\ : std_logic;
signal \N__30100\ : std_logic;
signal \N__30099\ : std_logic;
signal \N__30096\ : std_logic;
signal \N__30093\ : std_logic;
signal \N__30090\ : std_logic;
signal \N__30087\ : std_logic;
signal \N__30084\ : std_logic;
signal \N__30079\ : std_logic;
signal \N__30078\ : std_logic;
signal \N__30075\ : std_logic;
signal \N__30072\ : std_logic;
signal \N__30069\ : std_logic;
signal \N__30064\ : std_logic;
signal \N__30061\ : std_logic;
signal \N__30058\ : std_logic;
signal \N__30055\ : std_logic;
signal \N__30052\ : std_logic;
signal \N__30049\ : std_logic;
signal \N__30046\ : std_logic;
signal \N__30045\ : std_logic;
signal \N__30042\ : std_logic;
signal \N__30041\ : std_logic;
signal \N__30038\ : std_logic;
signal \N__30035\ : std_logic;
signal \N__30032\ : std_logic;
signal \N__30029\ : std_logic;
signal \N__30022\ : std_logic;
signal \N__30021\ : std_logic;
signal \N__30018\ : std_logic;
signal \N__30015\ : std_logic;
signal \N__30014\ : std_logic;
signal \N__30013\ : std_logic;
signal \N__30012\ : std_logic;
signal \N__30009\ : std_logic;
signal \N__30006\ : std_logic;
signal \N__30005\ : std_logic;
signal \N__30004\ : std_logic;
signal \N__30003\ : std_logic;
signal \N__30000\ : std_logic;
signal \N__29999\ : std_logic;
signal \N__29996\ : std_logic;
signal \N__29995\ : std_logic;
signal \N__29994\ : std_logic;
signal \N__29991\ : std_logic;
signal \N__29990\ : std_logic;
signal \N__29987\ : std_logic;
signal \N__29984\ : std_logic;
signal \N__29981\ : std_logic;
signal \N__29974\ : std_logic;
signal \N__29961\ : std_logic;
signal \N__29950\ : std_logic;
signal \N__29949\ : std_logic;
signal \N__29946\ : std_logic;
signal \N__29943\ : std_logic;
signal \N__29940\ : std_logic;
signal \N__29937\ : std_logic;
signal \N__29936\ : std_logic;
signal \N__29935\ : std_logic;
signal \N__29934\ : std_logic;
signal \N__29933\ : std_logic;
signal \N__29932\ : std_logic;
signal \N__29931\ : std_logic;
signal \N__29930\ : std_logic;
signal \N__29929\ : std_logic;
signal \N__29928\ : std_logic;
signal \N__29927\ : std_logic;
signal \N__29924\ : std_logic;
signal \N__29921\ : std_logic;
signal \N__29918\ : std_logic;
signal \N__29909\ : std_logic;
signal \N__29898\ : std_logic;
signal \N__29887\ : std_logic;
signal \N__29886\ : std_logic;
signal \N__29883\ : std_logic;
signal \N__29880\ : std_logic;
signal \N__29879\ : std_logic;
signal \N__29876\ : std_logic;
signal \N__29873\ : std_logic;
signal \N__29870\ : std_logic;
signal \N__29863\ : std_logic;
signal \N__29862\ : std_logic;
signal \N__29859\ : std_logic;
signal \N__29858\ : std_logic;
signal \N__29857\ : std_logic;
signal \N__29856\ : std_logic;
signal \N__29855\ : std_logic;
signal \N__29854\ : std_logic;
signal \N__29851\ : std_logic;
signal \N__29848\ : std_logic;
signal \N__29847\ : std_logic;
signal \N__29846\ : std_logic;
signal \N__29845\ : std_logic;
signal \N__29842\ : std_logic;
signal \N__29841\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29837\ : std_logic;
signal \N__29830\ : std_logic;
signal \N__29827\ : std_logic;
signal \N__29824\ : std_logic;
signal \N__29819\ : std_logic;
signal \N__29808\ : std_logic;
signal \N__29805\ : std_logic;
signal \N__29794\ : std_logic;
signal \N__29793\ : std_logic;
signal \N__29792\ : std_logic;
signal \N__29791\ : std_logic;
signal \N__29788\ : std_logic;
signal \N__29787\ : std_logic;
signal \N__29784\ : std_logic;
signal \N__29783\ : std_logic;
signal \N__29782\ : std_logic;
signal \N__29781\ : std_logic;
signal \N__29776\ : std_logic;
signal \N__29773\ : std_logic;
signal \N__29768\ : std_logic;
signal \N__29767\ : std_logic;
signal \N__29766\ : std_logic;
signal \N__29765\ : std_logic;
signal \N__29764\ : std_logic;
signal \N__29757\ : std_logic;
signal \N__29754\ : std_logic;
signal \N__29749\ : std_logic;
signal \N__29742\ : std_logic;
signal \N__29739\ : std_logic;
signal \N__29736\ : std_logic;
signal \N__29725\ : std_logic;
signal \N__29722\ : std_logic;
signal \N__29719\ : std_logic;
signal \N__29716\ : std_logic;
signal \N__29715\ : std_logic;
signal \N__29712\ : std_logic;
signal \N__29709\ : std_logic;
signal \N__29706\ : std_logic;
signal \N__29705\ : std_logic;
signal \N__29702\ : std_logic;
signal \N__29699\ : std_logic;
signal \N__29696\ : std_logic;
signal \N__29693\ : std_logic;
signal \N__29686\ : std_logic;
signal \N__29683\ : std_logic;
signal \N__29680\ : std_logic;
signal \N__29677\ : std_logic;
signal \N__29674\ : std_logic;
signal \N__29671\ : std_logic;
signal \N__29668\ : std_logic;
signal \N__29665\ : std_logic;
signal \N__29662\ : std_logic;
signal \N__29659\ : std_logic;
signal \N__29656\ : std_logic;
signal \N__29653\ : std_logic;
signal \N__29650\ : std_logic;
signal \N__29647\ : std_logic;
signal \N__29644\ : std_logic;
signal \N__29641\ : std_logic;
signal \N__29638\ : std_logic;
signal \N__29635\ : std_logic;
signal \N__29632\ : std_logic;
signal \N__29629\ : std_logic;
signal \N__29626\ : std_logic;
signal \N__29623\ : std_logic;
signal \N__29620\ : std_logic;
signal \N__29617\ : std_logic;
signal \N__29614\ : std_logic;
signal \N__29611\ : std_logic;
signal \N__29608\ : std_logic;
signal \N__29607\ : std_logic;
signal \N__29604\ : std_logic;
signal \N__29601\ : std_logic;
signal \N__29598\ : std_logic;
signal \N__29595\ : std_logic;
signal \N__29590\ : std_logic;
signal \N__29587\ : std_logic;
signal \N__29586\ : std_logic;
signal \N__29583\ : std_logic;
signal \N__29580\ : std_logic;
signal \N__29577\ : std_logic;
signal \N__29576\ : std_logic;
signal \N__29573\ : std_logic;
signal \N__29570\ : std_logic;
signal \N__29567\ : std_logic;
signal \N__29562\ : std_logic;
signal \N__29557\ : std_logic;
signal \N__29556\ : std_logic;
signal \N__29555\ : std_logic;
signal \N__29552\ : std_logic;
signal \N__29549\ : std_logic;
signal \N__29546\ : std_logic;
signal \N__29543\ : std_logic;
signal \N__29536\ : std_logic;
signal \N__29533\ : std_logic;
signal \N__29530\ : std_logic;
signal \N__29527\ : std_logic;
signal \N__29524\ : std_logic;
signal \N__29521\ : std_logic;
signal \N__29518\ : std_logic;
signal \N__29515\ : std_logic;
signal \N__29512\ : std_logic;
signal \N__29509\ : std_logic;
signal \N__29508\ : std_logic;
signal \N__29505\ : std_logic;
signal \N__29502\ : std_logic;
signal \N__29499\ : std_logic;
signal \N__29498\ : std_logic;
signal \N__29493\ : std_logic;
signal \N__29490\ : std_logic;
signal \N__29487\ : std_logic;
signal \N__29482\ : std_logic;
signal \N__29479\ : std_logic;
signal \N__29476\ : std_logic;
signal \N__29475\ : std_logic;
signal \N__29474\ : std_logic;
signal \N__29473\ : std_logic;
signal \N__29472\ : std_logic;
signal \N__29471\ : std_logic;
signal \N__29470\ : std_logic;
signal \N__29459\ : std_logic;
signal \N__29454\ : std_logic;
signal \N__29449\ : std_logic;
signal \N__29448\ : std_logic;
signal \N__29447\ : std_logic;
signal \N__29440\ : std_logic;
signal \N__29437\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29433\ : std_logic;
signal \N__29432\ : std_logic;
signal \N__29425\ : std_logic;
signal \N__29422\ : std_logic;
signal \N__29421\ : std_logic;
signal \N__29420\ : std_logic;
signal \N__29417\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29407\ : std_logic;
signal \N__29404\ : std_logic;
signal \N__29401\ : std_logic;
signal \N__29398\ : std_logic;
signal \N__29397\ : std_logic;
signal \N__29394\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29390\ : std_logic;
signal \N__29387\ : std_logic;
signal \N__29384\ : std_logic;
signal \N__29377\ : std_logic;
signal \N__29374\ : std_logic;
signal \N__29371\ : std_logic;
signal \N__29368\ : std_logic;
signal \N__29365\ : std_logic;
signal \N__29362\ : std_logic;
signal \N__29359\ : std_logic;
signal \N__29356\ : std_logic;
signal \N__29353\ : std_logic;
signal \N__29350\ : std_logic;
signal \N__29347\ : std_logic;
signal \N__29344\ : std_logic;
signal \N__29341\ : std_logic;
signal \N__29338\ : std_logic;
signal \N__29335\ : std_logic;
signal \N__29332\ : std_logic;
signal \N__29329\ : std_logic;
signal \N__29326\ : std_logic;
signal \N__29325\ : std_logic;
signal \N__29322\ : std_logic;
signal \N__29319\ : std_logic;
signal \N__29318\ : std_logic;
signal \N__29317\ : std_logic;
signal \N__29314\ : std_logic;
signal \N__29311\ : std_logic;
signal \N__29308\ : std_logic;
signal \N__29305\ : std_logic;
signal \N__29300\ : std_logic;
signal \N__29297\ : std_logic;
signal \N__29296\ : std_logic;
signal \N__29293\ : std_logic;
signal \N__29288\ : std_logic;
signal \N__29285\ : std_logic;
signal \N__29282\ : std_logic;
signal \N__29275\ : std_logic;
signal \N__29272\ : std_logic;
signal \N__29271\ : std_logic;
signal \N__29268\ : std_logic;
signal \N__29265\ : std_logic;
signal \N__29260\ : std_logic;
signal \N__29257\ : std_logic;
signal \N__29254\ : std_logic;
signal \N__29253\ : std_logic;
signal \N__29250\ : std_logic;
signal \N__29247\ : std_logic;
signal \N__29244\ : std_logic;
signal \N__29239\ : std_logic;
signal \N__29236\ : std_logic;
signal \N__29235\ : std_logic;
signal \N__29232\ : std_logic;
signal \N__29229\ : std_logic;
signal \N__29224\ : std_logic;
signal \N__29221\ : std_logic;
signal \N__29220\ : std_logic;
signal \N__29217\ : std_logic;
signal \N__29214\ : std_logic;
signal \N__29209\ : std_logic;
signal \N__29206\ : std_logic;
signal \N__29203\ : std_logic;
signal \N__29202\ : std_logic;
signal \N__29199\ : std_logic;
signal \N__29196\ : std_logic;
signal \N__29191\ : std_logic;
signal \N__29190\ : std_logic;
signal \N__29187\ : std_logic;
signal \N__29186\ : std_logic;
signal \N__29183\ : std_logic;
signal \N__29180\ : std_logic;
signal \N__29179\ : std_logic;
signal \N__29178\ : std_logic;
signal \N__29177\ : std_logic;
signal \N__29174\ : std_logic;
signal \N__29169\ : std_logic;
signal \N__29166\ : std_logic;
signal \N__29163\ : std_logic;
signal \N__29162\ : std_logic;
signal \N__29159\ : std_logic;
signal \N__29152\ : std_logic;
signal \N__29149\ : std_logic;
signal \N__29146\ : std_logic;
signal \N__29143\ : std_logic;
signal \N__29140\ : std_logic;
signal \N__29135\ : std_logic;
signal \N__29134\ : std_logic;
signal \N__29131\ : std_logic;
signal \N__29128\ : std_logic;
signal \N__29125\ : std_logic;
signal \N__29122\ : std_logic;
signal \N__29113\ : std_logic;
signal \N__29110\ : std_logic;
signal \N__29109\ : std_logic;
signal \N__29108\ : std_logic;
signal \N__29105\ : std_logic;
signal \N__29104\ : std_logic;
signal \N__29103\ : std_logic;
signal \N__29100\ : std_logic;
signal \N__29099\ : std_logic;
signal \N__29096\ : std_logic;
signal \N__29095\ : std_logic;
signal \N__29092\ : std_logic;
signal \N__29089\ : std_logic;
signal \N__29086\ : std_logic;
signal \N__29083\ : std_logic;
signal \N__29080\ : std_logic;
signal \N__29077\ : std_logic;
signal \N__29074\ : std_logic;
signal \N__29069\ : std_logic;
signal \N__29066\ : std_logic;
signal \N__29061\ : std_logic;
signal \N__29056\ : std_logic;
signal \N__29051\ : std_logic;
signal \N__29048\ : std_logic;
signal \N__29045\ : std_logic;
signal \N__29042\ : std_logic;
signal \N__29035\ : std_logic;
signal \N__29032\ : std_logic;
signal \N__29029\ : std_logic;
signal \N__29026\ : std_logic;
signal \N__29023\ : std_logic;
signal \N__29020\ : std_logic;
signal \N__29017\ : std_logic;
signal \N__29014\ : std_logic;
signal \N__29011\ : std_logic;
signal \N__29008\ : std_logic;
signal \N__29005\ : std_logic;
signal \N__29002\ : std_logic;
signal \N__28999\ : std_logic;
signal \N__28996\ : std_logic;
signal \N__28993\ : std_logic;
signal \N__28990\ : std_logic;
signal \N__28987\ : std_logic;
signal \N__28984\ : std_logic;
signal \N__28981\ : std_logic;
signal \N__28980\ : std_logic;
signal \N__28979\ : std_logic;
signal \N__28978\ : std_logic;
signal \N__28977\ : std_logic;
signal \N__28976\ : std_logic;
signal \N__28975\ : std_logic;
signal \N__28974\ : std_logic;
signal \N__28973\ : std_logic;
signal \N__28968\ : std_logic;
signal \N__28955\ : std_logic;
signal \N__28954\ : std_logic;
signal \N__28953\ : std_logic;
signal \N__28952\ : std_logic;
signal \N__28951\ : std_logic;
signal \N__28950\ : std_logic;
signal \N__28949\ : std_logic;
signal \N__28948\ : std_logic;
signal \N__28947\ : std_logic;
signal \N__28944\ : std_logic;
signal \N__28943\ : std_logic;
signal \N__28942\ : std_logic;
signal \N__28941\ : std_logic;
signal \N__28940\ : std_logic;
signal \N__28937\ : std_logic;
signal \N__28934\ : std_logic;
signal \N__28931\ : std_logic;
signal \N__28916\ : std_logic;
signal \N__28913\ : std_logic;
signal \N__28910\ : std_logic;
signal \N__28909\ : std_logic;
signal \N__28908\ : std_logic;
signal \N__28907\ : std_logic;
signal \N__28904\ : std_logic;
signal \N__28899\ : std_logic;
signal \N__28892\ : std_logic;
signal \N__28889\ : std_logic;
signal \N__28884\ : std_logic;
signal \N__28881\ : std_logic;
signal \N__28880\ : std_logic;
signal \N__28877\ : std_logic;
signal \N__28876\ : std_logic;
signal \N__28873\ : std_logic;
signal \N__28870\ : std_logic;
signal \N__28867\ : std_logic;
signal \N__28866\ : std_logic;
signal \N__28865\ : std_logic;
signal \N__28860\ : std_logic;
signal \N__28855\ : std_logic;
signal \N__28852\ : std_logic;
signal \N__28849\ : std_logic;
signal \N__28846\ : std_logic;
signal \N__28841\ : std_logic;
signal \N__28838\ : std_logic;
signal \N__28833\ : std_logic;
signal \N__28830\ : std_logic;
signal \N__28827\ : std_logic;
signal \N__28810\ : std_logic;
signal \N__28809\ : std_logic;
signal \N__28808\ : std_logic;
signal \N__28807\ : std_logic;
signal \N__28806\ : std_logic;
signal \N__28805\ : std_logic;
signal \N__28804\ : std_logic;
signal \N__28803\ : std_logic;
signal \N__28802\ : std_logic;
signal \N__28801\ : std_logic;
signal \N__28800\ : std_logic;
signal \N__28799\ : std_logic;
signal \N__28798\ : std_logic;
signal \N__28797\ : std_logic;
signal \N__28796\ : std_logic;
signal \N__28795\ : std_logic;
signal \N__28788\ : std_logic;
signal \N__28777\ : std_logic;
signal \N__28776\ : std_logic;
signal \N__28775\ : std_logic;
signal \N__28774\ : std_logic;
signal \N__28773\ : std_logic;
signal \N__28756\ : std_logic;
signal \N__28751\ : std_logic;
signal \N__28750\ : std_logic;
signal \N__28749\ : std_logic;
signal \N__28748\ : std_logic;
signal \N__28747\ : std_logic;
signal \N__28746\ : std_logic;
signal \N__28743\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28737\ : std_logic;
signal \N__28736\ : std_logic;
signal \N__28733\ : std_logic;
signal \N__28728\ : std_logic;
signal \N__28725\ : std_logic;
signal \N__28716\ : std_logic;
signal \N__28711\ : std_logic;
signal \N__28708\ : std_logic;
signal \N__28705\ : std_logic;
signal \N__28702\ : std_logic;
signal \N__28699\ : std_logic;
signal \N__28694\ : std_logic;
signal \N__28689\ : std_logic;
signal \N__28678\ : std_logic;
signal \N__28677\ : std_logic;
signal \N__28674\ : std_logic;
signal \N__28671\ : std_logic;
signal \N__28668\ : std_logic;
signal \N__28665\ : std_logic;
signal \N__28664\ : std_logic;
signal \N__28661\ : std_logic;
signal \N__28658\ : std_logic;
signal \N__28655\ : std_logic;
signal \N__28654\ : std_logic;
signal \N__28649\ : std_logic;
signal \N__28646\ : std_logic;
signal \N__28643\ : std_logic;
signal \N__28640\ : std_logic;
signal \N__28637\ : std_logic;
signal \N__28634\ : std_logic;
signal \N__28631\ : std_logic;
signal \N__28628\ : std_logic;
signal \N__28621\ : std_logic;
signal \N__28618\ : std_logic;
signal \N__28617\ : std_logic;
signal \N__28614\ : std_logic;
signal \N__28613\ : std_logic;
signal \N__28612\ : std_logic;
signal \N__28611\ : std_logic;
signal \N__28608\ : std_logic;
signal \N__28607\ : std_logic;
signal \N__28604\ : std_logic;
signal \N__28601\ : std_logic;
signal \N__28598\ : std_logic;
signal \N__28595\ : std_logic;
signal \N__28594\ : std_logic;
signal \N__28593\ : std_logic;
signal \N__28592\ : std_logic;
signal \N__28591\ : std_logic;
signal \N__28588\ : std_logic;
signal \N__28585\ : std_logic;
signal \N__28582\ : std_logic;
signal \N__28575\ : std_logic;
signal \N__28566\ : std_logic;
signal \N__28555\ : std_logic;
signal \N__28552\ : std_logic;
signal \N__28551\ : std_logic;
signal \N__28548\ : std_logic;
signal \N__28545\ : std_logic;
signal \N__28540\ : std_logic;
signal \N__28537\ : std_logic;
signal \N__28534\ : std_logic;
signal \N__28531\ : std_logic;
signal \N__28530\ : std_logic;
signal \N__28527\ : std_logic;
signal \N__28524\ : std_logic;
signal \N__28519\ : std_logic;
signal \N__28516\ : std_logic;
signal \N__28515\ : std_logic;
signal \N__28512\ : std_logic;
signal \N__28509\ : std_logic;
signal \N__28506\ : std_logic;
signal \N__28501\ : std_logic;
signal \N__28498\ : std_logic;
signal \N__28497\ : std_logic;
signal \N__28494\ : std_logic;
signal \N__28491\ : std_logic;
signal \N__28486\ : std_logic;
signal \N__28483\ : std_logic;
signal \N__28482\ : std_logic;
signal \N__28479\ : std_logic;
signal \N__28476\ : std_logic;
signal \N__28473\ : std_logic;
signal \N__28468\ : std_logic;
signal \N__28465\ : std_logic;
signal \N__28464\ : std_logic;
signal \N__28461\ : std_logic;
signal \N__28458\ : std_logic;
signal \N__28453\ : std_logic;
signal \N__28450\ : std_logic;
signal \N__28449\ : std_logic;
signal \N__28446\ : std_logic;
signal \N__28443\ : std_logic;
signal \N__28438\ : std_logic;
signal \N__28435\ : std_logic;
signal \N__28434\ : std_logic;
signal \N__28431\ : std_logic;
signal \N__28428\ : std_logic;
signal \N__28423\ : std_logic;
signal \N__28420\ : std_logic;
signal \N__28419\ : std_logic;
signal \N__28418\ : std_logic;
signal \N__28417\ : std_logic;
signal \N__28416\ : std_logic;
signal \N__28415\ : std_logic;
signal \N__28414\ : std_logic;
signal \N__28399\ : std_logic;
signal \N__28398\ : std_logic;
signal \N__28397\ : std_logic;
signal \N__28394\ : std_logic;
signal \N__28391\ : std_logic;
signal \N__28390\ : std_logic;
signal \N__28389\ : std_logic;
signal \N__28388\ : std_logic;
signal \N__28385\ : std_logic;
signal \N__28382\ : std_logic;
signal \N__28373\ : std_logic;
signal \N__28372\ : std_logic;
signal \N__28371\ : std_logic;
signal \N__28370\ : std_logic;
signal \N__28369\ : std_logic;
signal \N__28368\ : std_logic;
signal \N__28367\ : std_logic;
signal \N__28366\ : std_logic;
signal \N__28365\ : std_logic;
signal \N__28364\ : std_logic;
signal \N__28363\ : std_logic;
signal \N__28362\ : std_logic;
signal \N__28361\ : std_logic;
signal \N__28354\ : std_logic;
signal \N__28337\ : std_logic;
signal \N__28330\ : std_logic;
signal \N__28327\ : std_logic;
signal \N__28324\ : std_logic;
signal \N__28321\ : std_logic;
signal \N__28318\ : std_logic;
signal \N__28315\ : std_logic;
signal \N__28312\ : std_logic;
signal \N__28307\ : std_logic;
signal \N__28300\ : std_logic;
signal \N__28297\ : std_logic;
signal \N__28294\ : std_logic;
signal \N__28291\ : std_logic;
signal \N__28288\ : std_logic;
signal \N__28285\ : std_logic;
signal \N__28282\ : std_logic;
signal \N__28279\ : std_logic;
signal \N__28276\ : std_logic;
signal \N__28273\ : std_logic;
signal \N__28270\ : std_logic;
signal \N__28267\ : std_logic;
signal \N__28264\ : std_logic;
signal \N__28261\ : std_logic;
signal \N__28258\ : std_logic;
signal \N__28255\ : std_logic;
signal \N__28252\ : std_logic;
signal \N__28249\ : std_logic;
signal \N__28246\ : std_logic;
signal \N__28243\ : std_logic;
signal \N__28240\ : std_logic;
signal \N__28237\ : std_logic;
signal \N__28234\ : std_logic;
signal \N__28231\ : std_logic;
signal \N__28228\ : std_logic;
signal \N__28225\ : std_logic;
signal \N__28222\ : std_logic;
signal \N__28219\ : std_logic;
signal \N__28216\ : std_logic;
signal \N__28213\ : std_logic;
signal \N__28212\ : std_logic;
signal \N__28211\ : std_logic;
signal \N__28208\ : std_logic;
signal \N__28205\ : std_logic;
signal \N__28202\ : std_logic;
signal \N__28195\ : std_logic;
signal \N__28192\ : std_logic;
signal \N__28189\ : std_logic;
signal \N__28186\ : std_logic;
signal \N__28183\ : std_logic;
signal \N__28180\ : std_logic;
signal \N__28177\ : std_logic;
signal \N__28174\ : std_logic;
signal \N__28171\ : std_logic;
signal \N__28168\ : std_logic;
signal \N__28165\ : std_logic;
signal \N__28162\ : std_logic;
signal \N__28161\ : std_logic;
signal \N__28158\ : std_logic;
signal \N__28157\ : std_logic;
signal \N__28154\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28146\ : std_logic;
signal \N__28143\ : std_logic;
signal \N__28138\ : std_logic;
signal \N__28135\ : std_logic;
signal \N__28134\ : std_logic;
signal \N__28131\ : std_logic;
signal \N__28128\ : std_logic;
signal \N__28125\ : std_logic;
signal \N__28122\ : std_logic;
signal \N__28121\ : std_logic;
signal \N__28118\ : std_logic;
signal \N__28115\ : std_logic;
signal \N__28112\ : std_logic;
signal \N__28109\ : std_logic;
signal \N__28106\ : std_logic;
signal \N__28099\ : std_logic;
signal \N__28096\ : std_logic;
signal \N__28093\ : std_logic;
signal \N__28090\ : std_logic;
signal \N__28087\ : std_logic;
signal \N__28086\ : std_logic;
signal \N__28085\ : std_logic;
signal \N__28082\ : std_logic;
signal \N__28079\ : std_logic;
signal \N__28076\ : std_logic;
signal \N__28073\ : std_logic;
signal \N__28070\ : std_logic;
signal \N__28067\ : std_logic;
signal \N__28060\ : std_logic;
signal \N__28057\ : std_logic;
signal \N__28054\ : std_logic;
signal \N__28051\ : std_logic;
signal \N__28050\ : std_logic;
signal \N__28047\ : std_logic;
signal \N__28046\ : std_logic;
signal \N__28043\ : std_logic;
signal \N__28040\ : std_logic;
signal \N__28037\ : std_logic;
signal \N__28034\ : std_logic;
signal \N__28027\ : std_logic;
signal \N__28024\ : std_logic;
signal \N__28021\ : std_logic;
signal \N__28018\ : std_logic;
signal \N__28015\ : std_logic;
signal \N__28014\ : std_logic;
signal \N__28013\ : std_logic;
signal \N__28010\ : std_logic;
signal \N__28007\ : std_logic;
signal \N__28004\ : std_logic;
signal \N__27997\ : std_logic;
signal \N__27994\ : std_logic;
signal \N__27993\ : std_logic;
signal \N__27992\ : std_logic;
signal \N__27989\ : std_logic;
signal \N__27986\ : std_logic;
signal \N__27983\ : std_logic;
signal \N__27980\ : std_logic;
signal \N__27977\ : std_logic;
signal \N__27974\ : std_logic;
signal \N__27971\ : std_logic;
signal \N__27964\ : std_logic;
signal \N__27963\ : std_logic;
signal \N__27960\ : std_logic;
signal \N__27959\ : std_logic;
signal \N__27956\ : std_logic;
signal \N__27953\ : std_logic;
signal \N__27950\ : std_logic;
signal \N__27943\ : std_logic;
signal \N__27940\ : std_logic;
signal \N__27937\ : std_logic;
signal \N__27934\ : std_logic;
signal \N__27931\ : std_logic;
signal \N__27928\ : std_logic;
signal \N__27925\ : std_logic;
signal \N__27922\ : std_logic;
signal \N__27921\ : std_logic;
signal \N__27920\ : std_logic;
signal \N__27917\ : std_logic;
signal \N__27914\ : std_logic;
signal \N__27911\ : std_logic;
signal \N__27908\ : std_logic;
signal \N__27901\ : std_logic;
signal \N__27898\ : std_logic;
signal \N__27895\ : std_logic;
signal \N__27892\ : std_logic;
signal \N__27889\ : std_logic;
signal \N__27886\ : std_logic;
signal \N__27883\ : std_logic;
signal \N__27880\ : std_logic;
signal \N__27877\ : std_logic;
signal \N__27874\ : std_logic;
signal \N__27873\ : std_logic;
signal \N__27870\ : std_logic;
signal \N__27867\ : std_logic;
signal \N__27864\ : std_logic;
signal \N__27861\ : std_logic;
signal \N__27858\ : std_logic;
signal \N__27857\ : std_logic;
signal \N__27854\ : std_logic;
signal \N__27851\ : std_logic;
signal \N__27848\ : std_logic;
signal \N__27845\ : std_logic;
signal \N__27838\ : std_logic;
signal \N__27835\ : std_logic;
signal \N__27832\ : std_logic;
signal \N__27829\ : std_logic;
signal \N__27826\ : std_logic;
signal \N__27825\ : std_logic;
signal \N__27824\ : std_logic;
signal \N__27821\ : std_logic;
signal \N__27816\ : std_logic;
signal \N__27811\ : std_logic;
signal \N__27808\ : std_logic;
signal \N__27805\ : std_logic;
signal \N__27802\ : std_logic;
signal \N__27801\ : std_logic;
signal \N__27800\ : std_logic;
signal \N__27797\ : std_logic;
signal \N__27794\ : std_logic;
signal \N__27791\ : std_logic;
signal \N__27788\ : std_logic;
signal \N__27785\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27777\ : std_logic;
signal \N__27774\ : std_logic;
signal \N__27773\ : std_logic;
signal \N__27770\ : std_logic;
signal \N__27767\ : std_logic;
signal \N__27764\ : std_logic;
signal \N__27757\ : std_logic;
signal \N__27756\ : std_logic;
signal \N__27753\ : std_logic;
signal \N__27750\ : std_logic;
signal \N__27747\ : std_logic;
signal \N__27746\ : std_logic;
signal \N__27743\ : std_logic;
signal \N__27740\ : std_logic;
signal \N__27737\ : std_logic;
signal \N__27730\ : std_logic;
signal \N__27727\ : std_logic;
signal \N__27726\ : std_logic;
signal \N__27723\ : std_logic;
signal \N__27720\ : std_logic;
signal \N__27717\ : std_logic;
signal \N__27714\ : std_logic;
signal \N__27709\ : std_logic;
signal \N__27706\ : std_logic;
signal \N__27703\ : std_logic;
signal \N__27700\ : std_logic;
signal \N__27697\ : std_logic;
signal \N__27694\ : std_logic;
signal \N__27691\ : std_logic;
signal \N__27688\ : std_logic;
signal \N__27685\ : std_logic;
signal \N__27682\ : std_logic;
signal \N__27679\ : std_logic;
signal \N__27676\ : std_logic;
signal \N__27673\ : std_logic;
signal \N__27670\ : std_logic;
signal \N__27667\ : std_logic;
signal \N__27664\ : std_logic;
signal \N__27661\ : std_logic;
signal \N__27658\ : std_logic;
signal \N__27655\ : std_logic;
signal \N__27652\ : std_logic;
signal \N__27649\ : std_logic;
signal \N__27646\ : std_logic;
signal \N__27643\ : std_logic;
signal \N__27640\ : std_logic;
signal \N__27637\ : std_logic;
signal \N__27634\ : std_logic;
signal \N__27631\ : std_logic;
signal \N__27628\ : std_logic;
signal \N__27625\ : std_logic;
signal \N__27622\ : std_logic;
signal \N__27619\ : std_logic;
signal \N__27616\ : std_logic;
signal \N__27613\ : std_logic;
signal \N__27610\ : std_logic;
signal \N__27609\ : std_logic;
signal \N__27608\ : std_logic;
signal \N__27605\ : std_logic;
signal \N__27602\ : std_logic;
signal \N__27599\ : std_logic;
signal \N__27596\ : std_logic;
signal \N__27589\ : std_logic;
signal \N__27588\ : std_logic;
signal \N__27587\ : std_logic;
signal \N__27584\ : std_logic;
signal \N__27581\ : std_logic;
signal \N__27578\ : std_logic;
signal \N__27571\ : std_logic;
signal \N__27570\ : std_logic;
signal \N__27567\ : std_logic;
signal \N__27566\ : std_logic;
signal \N__27563\ : std_logic;
signal \N__27560\ : std_logic;
signal \N__27557\ : std_logic;
signal \N__27554\ : std_logic;
signal \N__27551\ : std_logic;
signal \N__27544\ : std_logic;
signal \N__27541\ : std_logic;
signal \N__27538\ : std_logic;
signal \N__27535\ : std_logic;
signal \N__27532\ : std_logic;
signal \N__27529\ : std_logic;
signal \N__27526\ : std_logic;
signal \N__27523\ : std_logic;
signal \N__27520\ : std_logic;
signal \N__27517\ : std_logic;
signal \N__27514\ : std_logic;
signal \N__27513\ : std_logic;
signal \N__27512\ : std_logic;
signal \N__27509\ : std_logic;
signal \N__27506\ : std_logic;
signal \N__27505\ : std_logic;
signal \N__27504\ : std_logic;
signal \N__27501\ : std_logic;
signal \N__27496\ : std_logic;
signal \N__27493\ : std_logic;
signal \N__27490\ : std_logic;
signal \N__27487\ : std_logic;
signal \N__27484\ : std_logic;
signal \N__27481\ : std_logic;
signal \N__27478\ : std_logic;
signal \N__27469\ : std_logic;
signal \N__27466\ : std_logic;
signal \N__27465\ : std_logic;
signal \N__27464\ : std_logic;
signal \N__27461\ : std_logic;
signal \N__27458\ : std_logic;
signal \N__27455\ : std_logic;
signal \N__27454\ : std_logic;
signal \N__27453\ : std_logic;
signal \N__27448\ : std_logic;
signal \N__27445\ : std_logic;
signal \N__27442\ : std_logic;
signal \N__27439\ : std_logic;
signal \N__27436\ : std_logic;
signal \N__27433\ : std_logic;
signal \N__27430\ : std_logic;
signal \N__27427\ : std_logic;
signal \N__27418\ : std_logic;
signal \N__27415\ : std_logic;
signal \N__27412\ : std_logic;
signal \N__27409\ : std_logic;
signal \N__27406\ : std_logic;
signal \N__27403\ : std_logic;
signal \N__27400\ : std_logic;
signal \N__27397\ : std_logic;
signal \N__27394\ : std_logic;
signal \N__27391\ : std_logic;
signal \N__27388\ : std_logic;
signal \N__27385\ : std_logic;
signal \N__27382\ : std_logic;
signal \N__27379\ : std_logic;
signal \N__27376\ : std_logic;
signal \N__27373\ : std_logic;
signal \N__27370\ : std_logic;
signal \N__27367\ : std_logic;
signal \N__27364\ : std_logic;
signal \N__27361\ : std_logic;
signal \N__27358\ : std_logic;
signal \N__27355\ : std_logic;
signal \N__27352\ : std_logic;
signal \N__27349\ : std_logic;
signal \N__27346\ : std_logic;
signal \N__27343\ : std_logic;
signal \N__27340\ : std_logic;
signal \N__27337\ : std_logic;
signal \N__27334\ : std_logic;
signal \N__27331\ : std_logic;
signal \N__27328\ : std_logic;
signal \N__27325\ : std_logic;
signal \N__27322\ : std_logic;
signal \N__27319\ : std_logic;
signal \N__27316\ : std_logic;
signal \N__27313\ : std_logic;
signal \N__27310\ : std_logic;
signal \N__27307\ : std_logic;
signal \N__27304\ : std_logic;
signal \N__27301\ : std_logic;
signal \N__27300\ : std_logic;
signal \N__27297\ : std_logic;
signal \N__27294\ : std_logic;
signal \N__27291\ : std_logic;
signal \N__27288\ : std_logic;
signal \N__27287\ : std_logic;
signal \N__27284\ : std_logic;
signal \N__27281\ : std_logic;
signal \N__27278\ : std_logic;
signal \N__27275\ : std_logic;
signal \N__27272\ : std_logic;
signal \N__27265\ : std_logic;
signal \N__27262\ : std_logic;
signal \N__27259\ : std_logic;
signal \N__27256\ : std_logic;
signal \N__27253\ : std_logic;
signal \N__27250\ : std_logic;
signal \N__27247\ : std_logic;
signal \N__27244\ : std_logic;
signal \N__27241\ : std_logic;
signal \N__27238\ : std_logic;
signal \N__27235\ : std_logic;
signal \N__27232\ : std_logic;
signal \N__27229\ : std_logic;
signal \N__27226\ : std_logic;
signal \N__27223\ : std_logic;
signal \N__27220\ : std_logic;
signal \N__27217\ : std_logic;
signal \N__27214\ : std_logic;
signal \N__27211\ : std_logic;
signal \N__27208\ : std_logic;
signal \N__27205\ : std_logic;
signal \N__27202\ : std_logic;
signal \N__27199\ : std_logic;
signal \N__27196\ : std_logic;
signal \N__27193\ : std_logic;
signal \N__27190\ : std_logic;
signal \N__27187\ : std_logic;
signal \N__27184\ : std_logic;
signal \N__27181\ : std_logic;
signal \N__27178\ : std_logic;
signal \N__27175\ : std_logic;
signal \N__27172\ : std_logic;
signal \N__27169\ : std_logic;
signal \N__27166\ : std_logic;
signal \N__27163\ : std_logic;
signal \N__27160\ : std_logic;
signal \N__27157\ : std_logic;
signal \N__27154\ : std_logic;
signal \N__27151\ : std_logic;
signal \N__27148\ : std_logic;
signal \N__27145\ : std_logic;
signal \N__27142\ : std_logic;
signal \N__27139\ : std_logic;
signal \N__27136\ : std_logic;
signal \N__27133\ : std_logic;
signal \N__27130\ : std_logic;
signal \N__27127\ : std_logic;
signal \N__27124\ : std_logic;
signal \N__27121\ : std_logic;
signal \N__27118\ : std_logic;
signal \N__27115\ : std_logic;
signal \N__27114\ : std_logic;
signal \N__27111\ : std_logic;
signal \N__27108\ : std_logic;
signal \N__27103\ : std_logic;
signal \N__27102\ : std_logic;
signal \N__27099\ : std_logic;
signal \N__27096\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27088\ : std_logic;
signal \N__27087\ : std_logic;
signal \N__27084\ : std_logic;
signal \N__27081\ : std_logic;
signal \N__27076\ : std_logic;
signal \N__27073\ : std_logic;
signal \N__27070\ : std_logic;
signal \N__27067\ : std_logic;
signal \N__27064\ : std_logic;
signal \N__27061\ : std_logic;
signal \N__27058\ : std_logic;
signal \N__27055\ : std_logic;
signal \N__27052\ : std_logic;
signal \N__27049\ : std_logic;
signal \N__27048\ : std_logic;
signal \N__27047\ : std_logic;
signal \N__27044\ : std_logic;
signal \N__27041\ : std_logic;
signal \N__27038\ : std_logic;
signal \N__27031\ : std_logic;
signal \N__27028\ : std_logic;
signal \N__27025\ : std_logic;
signal \N__27022\ : std_logic;
signal \N__27019\ : std_logic;
signal \N__27016\ : std_logic;
signal \N__27013\ : std_logic;
signal \N__27010\ : std_logic;
signal \N__27007\ : std_logic;
signal \N__27004\ : std_logic;
signal \N__27001\ : std_logic;
signal \N__26998\ : std_logic;
signal \N__26995\ : std_logic;
signal \N__26992\ : std_logic;
signal \N__26989\ : std_logic;
signal \N__26988\ : std_logic;
signal \N__26985\ : std_logic;
signal \N__26984\ : std_logic;
signal \N__26981\ : std_logic;
signal \N__26978\ : std_logic;
signal \N__26975\ : std_logic;
signal \N__26972\ : std_logic;
signal \N__26969\ : std_logic;
signal \N__26966\ : std_logic;
signal \N__26959\ : std_logic;
signal \N__26958\ : std_logic;
signal \N__26957\ : std_logic;
signal \N__26954\ : std_logic;
signal \N__26949\ : std_logic;
signal \N__26946\ : std_logic;
signal \N__26941\ : std_logic;
signal \N__26938\ : std_logic;
signal \N__26935\ : std_logic;
signal \N__26932\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26928\ : std_logic;
signal \N__26925\ : std_logic;
signal \N__26920\ : std_logic;
signal \N__26919\ : std_logic;
signal \N__26916\ : std_logic;
signal \N__26915\ : std_logic;
signal \N__26912\ : std_logic;
signal \N__26909\ : std_logic;
signal \N__26906\ : std_logic;
signal \N__26903\ : std_logic;
signal \N__26896\ : std_logic;
signal \N__26895\ : std_logic;
signal \N__26892\ : std_logic;
signal \N__26891\ : std_logic;
signal \N__26890\ : std_logic;
signal \N__26889\ : std_logic;
signal \N__26888\ : std_logic;
signal \N__26885\ : std_logic;
signal \N__26884\ : std_logic;
signal \N__26883\ : std_logic;
signal \N__26882\ : std_logic;
signal \N__26881\ : std_logic;
signal \N__26880\ : std_logic;
signal \N__26879\ : std_logic;
signal \N__26878\ : std_logic;
signal \N__26875\ : std_logic;
signal \N__26864\ : std_logic;
signal \N__26861\ : std_logic;
signal \N__26858\ : std_logic;
signal \N__26855\ : std_logic;
signal \N__26852\ : std_logic;
signal \N__26851\ : std_logic;
signal \N__26850\ : std_logic;
signal \N__26847\ : std_logic;
signal \N__26846\ : std_logic;
signal \N__26843\ : std_logic;
signal \N__26842\ : std_logic;
signal \N__26841\ : std_logic;
signal \N__26838\ : std_logic;
signal \N__26837\ : std_logic;
signal \N__26836\ : std_logic;
signal \N__26831\ : std_logic;
signal \N__26818\ : std_logic;
signal \N__26805\ : std_logic;
signal \N__26802\ : std_logic;
signal \N__26799\ : std_logic;
signal \N__26798\ : std_logic;
signal \N__26797\ : std_logic;
signal \N__26792\ : std_logic;
signal \N__26789\ : std_logic;
signal \N__26780\ : std_logic;
signal \N__26773\ : std_logic;
signal \N__26770\ : std_logic;
signal \N__26769\ : std_logic;
signal \N__26768\ : std_logic;
signal \N__26765\ : std_logic;
signal \N__26762\ : std_logic;
signal \N__26759\ : std_logic;
signal \N__26756\ : std_logic;
signal \N__26753\ : std_logic;
signal \N__26746\ : std_logic;
signal \N__26745\ : std_logic;
signal \N__26742\ : std_logic;
signal \N__26739\ : std_logic;
signal \N__26734\ : std_logic;
signal \N__26731\ : std_logic;
signal \N__26728\ : std_logic;
signal \N__26727\ : std_logic;
signal \N__26724\ : std_logic;
signal \N__26721\ : std_logic;
signal \N__26718\ : std_logic;
signal \N__26715\ : std_logic;
signal \N__26710\ : std_logic;
signal \N__26709\ : std_logic;
signal \N__26706\ : std_logic;
signal \N__26703\ : std_logic;
signal \N__26698\ : std_logic;
signal \N__26695\ : std_logic;
signal \N__26692\ : std_logic;
signal \N__26691\ : std_logic;
signal \N__26688\ : std_logic;
signal \N__26685\ : std_logic;
signal \N__26682\ : std_logic;
signal \N__26679\ : std_logic;
signal \N__26674\ : std_logic;
signal \N__26671\ : std_logic;
signal \N__26670\ : std_logic;
signal \N__26667\ : std_logic;
signal \N__26664\ : std_logic;
signal \N__26659\ : std_logic;
signal \N__26658\ : std_logic;
signal \N__26655\ : std_logic;
signal \N__26652\ : std_logic;
signal \N__26647\ : std_logic;
signal \N__26646\ : std_logic;
signal \N__26643\ : std_logic;
signal \N__26640\ : std_logic;
signal \N__26635\ : std_logic;
signal \N__26632\ : std_logic;
signal \N__26629\ : std_logic;
signal \N__26628\ : std_logic;
signal \N__26625\ : std_logic;
signal \N__26622\ : std_logic;
signal \N__26619\ : std_logic;
signal \N__26616\ : std_logic;
signal \N__26611\ : std_logic;
signal \N__26610\ : std_logic;
signal \N__26609\ : std_logic;
signal \N__26606\ : std_logic;
signal \N__26603\ : std_logic;
signal \N__26600\ : std_logic;
signal \N__26597\ : std_logic;
signal \N__26590\ : std_logic;
signal \N__26587\ : std_logic;
signal \N__26586\ : std_logic;
signal \N__26585\ : std_logic;
signal \N__26582\ : std_logic;
signal \N__26577\ : std_logic;
signal \N__26574\ : std_logic;
signal \N__26569\ : std_logic;
signal \N__26568\ : std_logic;
signal \N__26565\ : std_logic;
signal \N__26564\ : std_logic;
signal \N__26561\ : std_logic;
signal \N__26558\ : std_logic;
signal \N__26555\ : std_logic;
signal \N__26552\ : std_logic;
signal \N__26545\ : std_logic;
signal \N__26542\ : std_logic;
signal \N__26539\ : std_logic;
signal \N__26536\ : std_logic;
signal \N__26533\ : std_logic;
signal \N__26532\ : std_logic;
signal \N__26529\ : std_logic;
signal \N__26528\ : std_logic;
signal \N__26525\ : std_logic;
signal \N__26522\ : std_logic;
signal \N__26519\ : std_logic;
signal \N__26514\ : std_logic;
signal \N__26509\ : std_logic;
signal \N__26508\ : std_logic;
signal \N__26505\ : std_logic;
signal \N__26504\ : std_logic;
signal \N__26501\ : std_logic;
signal \N__26498\ : std_logic;
signal \N__26495\ : std_logic;
signal \N__26492\ : std_logic;
signal \N__26485\ : std_logic;
signal \N__26482\ : std_logic;
signal \N__26481\ : std_logic;
signal \N__26480\ : std_logic;
signal \N__26477\ : std_logic;
signal \N__26474\ : std_logic;
signal \N__26471\ : std_logic;
signal \N__26468\ : std_logic;
signal \N__26465\ : std_logic;
signal \N__26458\ : std_logic;
signal \N__26455\ : std_logic;
signal \N__26452\ : std_logic;
signal \N__26451\ : std_logic;
signal \N__26450\ : std_logic;
signal \N__26447\ : std_logic;
signal \N__26444\ : std_logic;
signal \N__26441\ : std_logic;
signal \N__26438\ : std_logic;
signal \N__26435\ : std_logic;
signal \N__26428\ : std_logic;
signal \N__26427\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26423\ : std_logic;
signal \N__26418\ : std_logic;
signal \N__26415\ : std_logic;
signal \N__26410\ : std_logic;
signal \N__26409\ : std_logic;
signal \N__26408\ : std_logic;
signal \N__26405\ : std_logic;
signal \N__26402\ : std_logic;
signal \N__26399\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26389\ : std_logic;
signal \N__26388\ : std_logic;
signal \N__26387\ : std_logic;
signal \N__26384\ : std_logic;
signal \N__26381\ : std_logic;
signal \N__26378\ : std_logic;
signal \N__26375\ : std_logic;
signal \N__26372\ : std_logic;
signal \N__26365\ : std_logic;
signal \N__26364\ : std_logic;
signal \N__26363\ : std_logic;
signal \N__26360\ : std_logic;
signal \N__26357\ : std_logic;
signal \N__26354\ : std_logic;
signal \N__26351\ : std_logic;
signal \N__26348\ : std_logic;
signal \N__26345\ : std_logic;
signal \N__26342\ : std_logic;
signal \N__26335\ : std_logic;
signal \N__26332\ : std_logic;
signal \N__26329\ : std_logic;
signal \N__26326\ : std_logic;
signal \N__26323\ : std_logic;
signal \N__26320\ : std_logic;
signal \N__26317\ : std_logic;
signal \N__26314\ : std_logic;
signal \N__26311\ : std_logic;
signal \N__26308\ : std_logic;
signal \N__26307\ : std_logic;
signal \N__26304\ : std_logic;
signal \N__26301\ : std_logic;
signal \N__26296\ : std_logic;
signal \N__26293\ : std_logic;
signal \N__26292\ : std_logic;
signal \N__26289\ : std_logic;
signal \N__26286\ : std_logic;
signal \N__26283\ : std_logic;
signal \N__26280\ : std_logic;
signal \N__26275\ : std_logic;
signal \N__26272\ : std_logic;
signal \N__26269\ : std_logic;
signal \N__26266\ : std_logic;
signal \N__26263\ : std_logic;
signal \N__26262\ : std_logic;
signal \N__26259\ : std_logic;
signal \N__26258\ : std_logic;
signal \N__26255\ : std_logic;
signal \N__26252\ : std_logic;
signal \N__26247\ : std_logic;
signal \N__26242\ : std_logic;
signal \N__26239\ : std_logic;
signal \N__26236\ : std_logic;
signal \N__26233\ : std_logic;
signal \N__26230\ : std_logic;
signal \N__26227\ : std_logic;
signal \N__26224\ : std_logic;
signal \N__26221\ : std_logic;
signal \N__26218\ : std_logic;
signal \N__26215\ : std_logic;
signal \N__26212\ : std_logic;
signal \N__26209\ : std_logic;
signal \N__26208\ : std_logic;
signal \N__26207\ : std_logic;
signal \N__26204\ : std_logic;
signal \N__26199\ : std_logic;
signal \N__26194\ : std_logic;
signal \N__26191\ : std_logic;
signal \N__26188\ : std_logic;
signal \N__26185\ : std_logic;
signal \N__26184\ : std_logic;
signal \N__26181\ : std_logic;
signal \N__26178\ : std_logic;
signal \N__26175\ : std_logic;
signal \N__26172\ : std_logic;
signal \N__26167\ : std_logic;
signal \N__26164\ : std_logic;
signal \N__26161\ : std_logic;
signal \N__26158\ : std_logic;
signal \N__26155\ : std_logic;
signal \N__26152\ : std_logic;
signal \N__26149\ : std_logic;
signal \N__26148\ : std_logic;
signal \N__26145\ : std_logic;
signal \N__26142\ : std_logic;
signal \N__26139\ : std_logic;
signal \N__26136\ : std_logic;
signal \N__26133\ : std_logic;
signal \N__26130\ : std_logic;
signal \N__26127\ : std_logic;
signal \N__26124\ : std_logic;
signal \N__26119\ : std_logic;
signal \N__26116\ : std_logic;
signal \N__26113\ : std_logic;
signal \N__26110\ : std_logic;
signal \N__26107\ : std_logic;
signal \N__26104\ : std_logic;
signal \N__26101\ : std_logic;
signal \N__26100\ : std_logic;
signal \N__26097\ : std_logic;
signal \N__26096\ : std_logic;
signal \N__26093\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26087\ : std_logic;
signal \N__26084\ : std_logic;
signal \N__26077\ : std_logic;
signal \N__26074\ : std_logic;
signal \N__26071\ : std_logic;
signal \N__26070\ : std_logic;
signal \N__26069\ : std_logic;
signal \N__26066\ : std_logic;
signal \N__26063\ : std_logic;
signal \N__26060\ : std_logic;
signal \N__26057\ : std_logic;
signal \N__26054\ : std_logic;
signal \N__26047\ : std_logic;
signal \N__26044\ : std_logic;
signal \N__26041\ : std_logic;
signal \N__26038\ : std_logic;
signal \N__26035\ : std_logic;
signal \N__26032\ : std_logic;
signal \N__26031\ : std_logic;
signal \N__26028\ : std_logic;
signal \N__26027\ : std_logic;
signal \N__26024\ : std_logic;
signal \N__26021\ : std_logic;
signal \N__26016\ : std_logic;
signal \N__26011\ : std_logic;
signal \N__26008\ : std_logic;
signal \N__26005\ : std_logic;
signal \N__26002\ : std_logic;
signal \N__25999\ : std_logic;
signal \N__25996\ : std_logic;
signal \N__25993\ : std_logic;
signal \N__25992\ : std_logic;
signal \N__25989\ : std_logic;
signal \N__25986\ : std_logic;
signal \N__25983\ : std_logic;
signal \N__25982\ : std_logic;
signal \N__25977\ : std_logic;
signal \N__25974\ : std_logic;
signal \N__25969\ : std_logic;
signal \N__25968\ : std_logic;
signal \N__25965\ : std_logic;
signal \N__25962\ : std_logic;
signal \N__25961\ : std_logic;
signal \N__25958\ : std_logic;
signal \N__25955\ : std_logic;
signal \N__25952\ : std_logic;
signal \N__25949\ : std_logic;
signal \N__25946\ : std_logic;
signal \N__25939\ : std_logic;
signal \N__25938\ : std_logic;
signal \N__25937\ : std_logic;
signal \N__25934\ : std_logic;
signal \N__25931\ : std_logic;
signal \N__25930\ : std_logic;
signal \N__25927\ : std_logic;
signal \N__25920\ : std_logic;
signal \N__25917\ : std_logic;
signal \N__25912\ : std_logic;
signal \N__25911\ : std_logic;
signal \N__25910\ : std_logic;
signal \N__25905\ : std_logic;
signal \N__25902\ : std_logic;
signal \N__25897\ : std_logic;
signal \N__25894\ : std_logic;
signal \N__25893\ : std_logic;
signal \N__25890\ : std_logic;
signal \N__25889\ : std_logic;
signal \N__25886\ : std_logic;
signal \N__25883\ : std_logic;
signal \N__25880\ : std_logic;
signal \N__25873\ : std_logic;
signal \N__25872\ : std_logic;
signal \N__25869\ : std_logic;
signal \N__25866\ : std_logic;
signal \N__25863\ : std_logic;
signal \N__25860\ : std_logic;
signal \N__25857\ : std_logic;
signal \N__25856\ : std_logic;
signal \N__25853\ : std_logic;
signal \N__25850\ : std_logic;
signal \N__25847\ : std_logic;
signal \N__25840\ : std_logic;
signal \N__25837\ : std_logic;
signal \N__25834\ : std_logic;
signal \N__25831\ : std_logic;
signal \N__25828\ : std_logic;
signal \N__25825\ : std_logic;
signal \N__25822\ : std_logic;
signal \N__25819\ : std_logic;
signal \N__25816\ : std_logic;
signal \N__25813\ : std_logic;
signal \N__25812\ : std_logic;
signal \N__25809\ : std_logic;
signal \N__25808\ : std_logic;
signal \N__25805\ : std_logic;
signal \N__25802\ : std_logic;
signal \N__25799\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25793\ : std_logic;
signal \N__25786\ : std_logic;
signal \N__25785\ : std_logic;
signal \N__25782\ : std_logic;
signal \N__25779\ : std_logic;
signal \N__25774\ : std_logic;
signal \N__25771\ : std_logic;
signal \N__25768\ : std_logic;
signal \N__25765\ : std_logic;
signal \N__25762\ : std_logic;
signal \N__25759\ : std_logic;
signal \N__25756\ : std_logic;
signal \N__25753\ : std_logic;
signal \N__25750\ : std_logic;
signal \N__25747\ : std_logic;
signal \N__25746\ : std_logic;
signal \N__25743\ : std_logic;
signal \N__25740\ : std_logic;
signal \N__25737\ : std_logic;
signal \N__25734\ : std_logic;
signal \N__25729\ : std_logic;
signal \N__25726\ : std_logic;
signal \N__25723\ : std_logic;
signal \N__25720\ : std_logic;
signal \N__25717\ : std_logic;
signal \N__25714\ : std_logic;
signal \N__25711\ : std_logic;
signal \N__25710\ : std_logic;
signal \N__25707\ : std_logic;
signal \N__25706\ : std_logic;
signal \N__25703\ : std_logic;
signal \N__25700\ : std_logic;
signal \N__25697\ : std_logic;
signal \N__25694\ : std_logic;
signal \N__25691\ : std_logic;
signal \N__25688\ : std_logic;
signal \N__25685\ : std_logic;
signal \N__25682\ : std_logic;
signal \N__25675\ : std_logic;
signal \N__25672\ : std_logic;
signal \N__25669\ : std_logic;
signal \N__25668\ : std_logic;
signal \N__25665\ : std_logic;
signal \N__25662\ : std_logic;
signal \N__25659\ : std_logic;
signal \N__25656\ : std_logic;
signal \N__25651\ : std_logic;
signal \N__25648\ : std_logic;
signal \N__25645\ : std_logic;
signal \N__25642\ : std_logic;
signal \N__25639\ : std_logic;
signal \N__25636\ : std_logic;
signal \N__25633\ : std_logic;
signal \N__25630\ : std_logic;
signal \N__25627\ : std_logic;
signal \N__25624\ : std_logic;
signal \N__25621\ : std_logic;
signal \N__25618\ : std_logic;
signal \N__25615\ : std_logic;
signal \N__25612\ : std_logic;
signal \N__25609\ : std_logic;
signal \N__25606\ : std_logic;
signal \N__25603\ : std_logic;
signal \N__25600\ : std_logic;
signal \N__25597\ : std_logic;
signal \N__25594\ : std_logic;
signal \N__25591\ : std_logic;
signal \N__25588\ : std_logic;
signal \N__25585\ : std_logic;
signal \N__25582\ : std_logic;
signal \N__25579\ : std_logic;
signal \N__25578\ : std_logic;
signal \N__25575\ : std_logic;
signal \N__25572\ : std_logic;
signal \N__25567\ : std_logic;
signal \N__25564\ : std_logic;
signal \N__25563\ : std_logic;
signal \N__25560\ : std_logic;
signal \N__25557\ : std_logic;
signal \N__25552\ : std_logic;
signal \N__25549\ : std_logic;
signal \N__25548\ : std_logic;
signal \N__25545\ : std_logic;
signal \N__25542\ : std_logic;
signal \N__25537\ : std_logic;
signal \N__25534\ : std_logic;
signal \N__25533\ : std_logic;
signal \N__25530\ : std_logic;
signal \N__25527\ : std_logic;
signal \N__25522\ : std_logic;
signal \N__25519\ : std_logic;
signal \N__25518\ : std_logic;
signal \N__25515\ : std_logic;
signal \N__25512\ : std_logic;
signal \N__25507\ : std_logic;
signal \N__25504\ : std_logic;
signal \N__25503\ : std_logic;
signal \N__25500\ : std_logic;
signal \N__25497\ : std_logic;
signal \N__25492\ : std_logic;
signal \N__25489\ : std_logic;
signal \N__25486\ : std_logic;
signal \N__25483\ : std_logic;
signal \N__25480\ : std_logic;
signal \N__25477\ : std_logic;
signal \N__25474\ : std_logic;
signal \N__25471\ : std_logic;
signal \N__25468\ : std_logic;
signal \N__25465\ : std_logic;
signal \N__25464\ : std_logic;
signal \N__25463\ : std_logic;
signal \N__25460\ : std_logic;
signal \N__25457\ : std_logic;
signal \N__25454\ : std_logic;
signal \N__25451\ : std_logic;
signal \N__25444\ : std_logic;
signal \N__25443\ : std_logic;
signal \N__25440\ : std_logic;
signal \N__25437\ : std_logic;
signal \N__25432\ : std_logic;
signal \N__25429\ : std_logic;
signal \N__25428\ : std_logic;
signal \N__25425\ : std_logic;
signal \N__25424\ : std_logic;
signal \N__25421\ : std_logic;
signal \N__25418\ : std_logic;
signal \N__25415\ : std_logic;
signal \N__25412\ : std_logic;
signal \N__25405\ : std_logic;
signal \N__25402\ : std_logic;
signal \N__25401\ : std_logic;
signal \N__25398\ : std_logic;
signal \N__25395\ : std_logic;
signal \N__25392\ : std_logic;
signal \N__25389\ : std_logic;
signal \N__25386\ : std_logic;
signal \N__25381\ : std_logic;
signal \N__25378\ : std_logic;
signal \N__25377\ : std_logic;
signal \N__25374\ : std_logic;
signal \N__25371\ : std_logic;
signal \N__25366\ : std_logic;
signal \N__25363\ : std_logic;
signal \N__25362\ : std_logic;
signal \N__25359\ : std_logic;
signal \N__25356\ : std_logic;
signal \N__25351\ : std_logic;
signal \N__25348\ : std_logic;
signal \N__25347\ : std_logic;
signal \N__25344\ : std_logic;
signal \N__25341\ : std_logic;
signal \N__25336\ : std_logic;
signal \N__25333\ : std_logic;
signal \N__25332\ : std_logic;
signal \N__25329\ : std_logic;
signal \N__25326\ : std_logic;
signal \N__25321\ : std_logic;
signal \N__25318\ : std_logic;
signal \N__25317\ : std_logic;
signal \N__25314\ : std_logic;
signal \N__25311\ : std_logic;
signal \N__25306\ : std_logic;
signal \N__25303\ : std_logic;
signal \N__25302\ : std_logic;
signal \N__25299\ : std_logic;
signal \N__25296\ : std_logic;
signal \N__25291\ : std_logic;
signal \N__25288\ : std_logic;
signal \N__25287\ : std_logic;
signal \N__25286\ : std_logic;
signal \N__25283\ : std_logic;
signal \N__25278\ : std_logic;
signal \N__25275\ : std_logic;
signal \N__25270\ : std_logic;
signal \N__25267\ : std_logic;
signal \N__25266\ : std_logic;
signal \N__25263\ : std_logic;
signal \N__25260\ : std_logic;
signal \N__25255\ : std_logic;
signal \N__25252\ : std_logic;
signal \N__25249\ : std_logic;
signal \N__25248\ : std_logic;
signal \N__25247\ : std_logic;
signal \N__25244\ : std_logic;
signal \N__25241\ : std_logic;
signal \N__25238\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25232\ : std_logic;
signal \N__25229\ : std_logic;
signal \N__25222\ : std_logic;
signal \N__25221\ : std_logic;
signal \N__25218\ : std_logic;
signal \N__25215\ : std_logic;
signal \N__25210\ : std_logic;
signal \N__25207\ : std_logic;
signal \N__25204\ : std_logic;
signal \N__25201\ : std_logic;
signal \N__25198\ : std_logic;
signal \N__25197\ : std_logic;
signal \N__25194\ : std_logic;
signal \N__25193\ : std_logic;
signal \N__25190\ : std_logic;
signal \N__25187\ : std_logic;
signal \N__25184\ : std_logic;
signal \N__25181\ : std_logic;
signal \N__25174\ : std_logic;
signal \N__25171\ : std_logic;
signal \N__25168\ : std_logic;
signal \N__25165\ : std_logic;
signal \N__25162\ : std_logic;
signal \N__25159\ : std_logic;
signal \N__25156\ : std_logic;
signal \N__25153\ : std_logic;
signal \N__25150\ : std_logic;
signal \N__25149\ : std_logic;
signal \N__25148\ : std_logic;
signal \N__25145\ : std_logic;
signal \N__25140\ : std_logic;
signal \N__25137\ : std_logic;
signal \N__25132\ : std_logic;
signal \N__25129\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25123\ : std_logic;
signal \N__25122\ : std_logic;
signal \N__25121\ : std_logic;
signal \N__25118\ : std_logic;
signal \N__25113\ : std_logic;
signal \N__25110\ : std_logic;
signal \N__25105\ : std_logic;
signal \N__25102\ : std_logic;
signal \N__25099\ : std_logic;
signal \N__25096\ : std_logic;
signal \N__25093\ : std_logic;
signal \N__25090\ : std_logic;
signal \N__25087\ : std_logic;
signal \N__25084\ : std_logic;
signal \N__25081\ : std_logic;
signal \N__25078\ : std_logic;
signal \N__25077\ : std_logic;
signal \N__25076\ : std_logic;
signal \N__25071\ : std_logic;
signal \N__25068\ : std_logic;
signal \N__25063\ : std_logic;
signal \N__25060\ : std_logic;
signal \N__25057\ : std_logic;
signal \N__25054\ : std_logic;
signal \N__25051\ : std_logic;
signal \N__25048\ : std_logic;
signal \N__25045\ : std_logic;
signal \N__25042\ : std_logic;
signal \N__25041\ : std_logic;
signal \N__25038\ : std_logic;
signal \N__25035\ : std_logic;
signal \N__25032\ : std_logic;
signal \N__25027\ : std_logic;
signal \N__25024\ : std_logic;
signal \N__25021\ : std_logic;
signal \N__25018\ : std_logic;
signal \N__25015\ : std_logic;
signal \N__25012\ : std_logic;
signal \N__25009\ : std_logic;
signal \N__25008\ : std_logic;
signal \N__25007\ : std_logic;
signal \N__25004\ : std_logic;
signal \N__25001\ : std_logic;
signal \N__24998\ : std_logic;
signal \N__24997\ : std_logic;
signal \N__24990\ : std_logic;
signal \N__24989\ : std_logic;
signal \N__24986\ : std_logic;
signal \N__24983\ : std_logic;
signal \N__24978\ : std_logic;
signal \N__24975\ : std_logic;
signal \N__24972\ : std_logic;
signal \N__24969\ : std_logic;
signal \N__24966\ : std_logic;
signal \N__24963\ : std_logic;
signal \N__24958\ : std_logic;
signal \N__24955\ : std_logic;
signal \N__24952\ : std_logic;
signal \N__24949\ : std_logic;
signal \N__24946\ : std_logic;
signal \N__24943\ : std_logic;
signal \N__24940\ : std_logic;
signal \N__24937\ : std_logic;
signal \N__24934\ : std_logic;
signal \N__24931\ : std_logic;
signal \N__24928\ : std_logic;
signal \N__24925\ : std_logic;
signal \N__24922\ : std_logic;
signal \N__24919\ : std_logic;
signal \N__24916\ : std_logic;
signal \N__24913\ : std_logic;
signal \N__24910\ : std_logic;
signal \N__24907\ : std_logic;
signal \N__24904\ : std_logic;
signal \N__24903\ : std_logic;
signal \N__24900\ : std_logic;
signal \N__24899\ : std_logic;
signal \N__24896\ : std_logic;
signal \N__24891\ : std_logic;
signal \N__24886\ : std_logic;
signal \N__24885\ : std_logic;
signal \N__24882\ : std_logic;
signal \N__24879\ : std_logic;
signal \N__24874\ : std_logic;
signal \N__24871\ : std_logic;
signal \N__24870\ : std_logic;
signal \N__24867\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24859\ : std_logic;
signal \N__24856\ : std_logic;
signal \N__24855\ : std_logic;
signal \N__24850\ : std_logic;
signal \N__24847\ : std_logic;
signal \N__24844\ : std_logic;
signal \N__24841\ : std_logic;
signal \N__24838\ : std_logic;
signal \N__24837\ : std_logic;
signal \N__24834\ : std_logic;
signal \N__24831\ : std_logic;
signal \N__24828\ : std_logic;
signal \N__24825\ : std_logic;
signal \N__24820\ : std_logic;
signal \N__24817\ : std_logic;
signal \N__24814\ : std_logic;
signal \N__24811\ : std_logic;
signal \N__24808\ : std_logic;
signal \N__24807\ : std_logic;
signal \N__24804\ : std_logic;
signal \N__24801\ : std_logic;
signal \N__24796\ : std_logic;
signal \N__24795\ : std_logic;
signal \N__24792\ : std_logic;
signal \N__24789\ : std_logic;
signal \N__24784\ : std_logic;
signal \N__24783\ : std_logic;
signal \N__24780\ : std_logic;
signal \N__24777\ : std_logic;
signal \N__24774\ : std_logic;
signal \N__24769\ : std_logic;
signal \N__24768\ : std_logic;
signal \N__24765\ : std_logic;
signal \N__24762\ : std_logic;
signal \N__24757\ : std_logic;
signal \N__24756\ : std_logic;
signal \N__24753\ : std_logic;
signal \N__24750\ : std_logic;
signal \N__24745\ : std_logic;
signal \N__24744\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24738\ : std_logic;
signal \N__24733\ : std_logic;
signal \N__24730\ : std_logic;
signal \N__24729\ : std_logic;
signal \N__24726\ : std_logic;
signal \N__24723\ : std_logic;
signal \N__24718\ : std_logic;
signal \N__24715\ : std_logic;
signal \N__24712\ : std_logic;
signal \N__24711\ : std_logic;
signal \N__24708\ : std_logic;
signal \N__24705\ : std_logic;
signal \N__24700\ : std_logic;
signal \N__24697\ : std_logic;
signal \N__24694\ : std_logic;
signal \N__24691\ : std_logic;
signal \N__24690\ : std_logic;
signal \N__24687\ : std_logic;
signal \N__24684\ : std_logic;
signal \N__24683\ : std_logic;
signal \N__24678\ : std_logic;
signal \N__24675\ : std_logic;
signal \N__24672\ : std_logic;
signal \N__24667\ : std_logic;
signal \N__24666\ : std_logic;
signal \N__24661\ : std_logic;
signal \N__24658\ : std_logic;
signal \N__24657\ : std_logic;
signal \N__24654\ : std_logic;
signal \N__24651\ : std_logic;
signal \N__24646\ : std_logic;
signal \N__24645\ : std_logic;
signal \N__24644\ : std_logic;
signal \N__24641\ : std_logic;
signal \N__24638\ : std_logic;
signal \N__24635\ : std_logic;
signal \N__24632\ : std_logic;
signal \N__24629\ : std_logic;
signal \N__24626\ : std_logic;
signal \N__24623\ : std_logic;
signal \N__24616\ : std_logic;
signal \N__24613\ : std_logic;
signal \N__24612\ : std_logic;
signal \N__24611\ : std_logic;
signal \N__24608\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24602\ : std_logic;
signal \N__24595\ : std_logic;
signal \N__24592\ : std_logic;
signal \N__24589\ : std_logic;
signal \N__24586\ : std_logic;
signal \N__24583\ : std_logic;
signal \N__24580\ : std_logic;
signal \N__24577\ : std_logic;
signal \N__24574\ : std_logic;
signal \N__24573\ : std_logic;
signal \N__24570\ : std_logic;
signal \N__24567\ : std_logic;
signal \N__24562\ : std_logic;
signal \N__24559\ : std_logic;
signal \N__24558\ : std_logic;
signal \N__24553\ : std_logic;
signal \N__24550\ : std_logic;
signal \N__24547\ : std_logic;
signal \N__24544\ : std_logic;
signal \N__24541\ : std_logic;
signal \N__24538\ : std_logic;
signal \N__24535\ : std_logic;
signal \N__24532\ : std_logic;
signal \N__24529\ : std_logic;
signal \N__24526\ : std_logic;
signal \N__24523\ : std_logic;
signal \N__24520\ : std_logic;
signal \N__24517\ : std_logic;
signal \N__24514\ : std_logic;
signal \N__24513\ : std_logic;
signal \N__24510\ : std_logic;
signal \N__24507\ : std_logic;
signal \N__24504\ : std_logic;
signal \N__24501\ : std_logic;
signal \N__24498\ : std_logic;
signal \N__24495\ : std_logic;
signal \N__24492\ : std_logic;
signal \N__24489\ : std_logic;
signal \N__24486\ : std_logic;
signal \N__24483\ : std_logic;
signal \N__24480\ : std_logic;
signal \N__24477\ : std_logic;
signal \N__24474\ : std_logic;
signal \N__24471\ : std_logic;
signal \N__24468\ : std_logic;
signal \N__24465\ : std_logic;
signal \N__24462\ : std_logic;
signal \N__24457\ : std_logic;
signal \N__24454\ : std_logic;
signal \N__24453\ : std_logic;
signal \N__24450\ : std_logic;
signal \N__24447\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24443\ : std_logic;
signal \N__24438\ : std_logic;
signal \N__24433\ : std_logic;
signal \N__24432\ : std_logic;
signal \N__24427\ : std_logic;
signal \N__24424\ : std_logic;
signal \N__24421\ : std_logic;
signal \N__24420\ : std_logic;
signal \N__24417\ : std_logic;
signal \N__24414\ : std_logic;
signal \N__24413\ : std_logic;
signal \N__24410\ : std_logic;
signal \N__24407\ : std_logic;
signal \N__24404\ : std_logic;
signal \N__24399\ : std_logic;
signal \N__24394\ : std_logic;
signal \N__24391\ : std_logic;
signal \N__24388\ : std_logic;
signal \N__24385\ : std_logic;
signal \N__24382\ : std_logic;
signal \N__24379\ : std_logic;
signal \N__24376\ : std_logic;
signal \N__24373\ : std_logic;
signal \N__24370\ : std_logic;
signal \N__24367\ : std_logic;
signal \N__24364\ : std_logic;
signal \N__24361\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24355\ : std_logic;
signal \N__24352\ : std_logic;
signal \N__24349\ : std_logic;
signal \N__24346\ : std_logic;
signal \N__24343\ : std_logic;
signal \N__24342\ : std_logic;
signal \N__24339\ : std_logic;
signal \N__24338\ : std_logic;
signal \N__24335\ : std_logic;
signal \N__24332\ : std_logic;
signal \N__24329\ : std_logic;
signal \N__24326\ : std_logic;
signal \N__24323\ : std_logic;
signal \N__24320\ : std_logic;
signal \N__24315\ : std_logic;
signal \N__24310\ : std_logic;
signal \N__24309\ : std_logic;
signal \N__24306\ : std_logic;
signal \N__24303\ : std_logic;
signal \N__24300\ : std_logic;
signal \N__24297\ : std_logic;
signal \N__24292\ : std_logic;
signal \N__24289\ : std_logic;
signal \N__24286\ : std_logic;
signal \N__24283\ : std_logic;
signal \N__24280\ : std_logic;
signal \N__24279\ : std_logic;
signal \N__24276\ : std_logic;
signal \N__24273\ : std_logic;
signal \N__24268\ : std_logic;
signal \N__24265\ : std_logic;
signal \N__24262\ : std_logic;
signal \N__24259\ : std_logic;
signal \N__24256\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24252\ : std_logic;
signal \N__24251\ : std_logic;
signal \N__24248\ : std_logic;
signal \N__24245\ : std_logic;
signal \N__24242\ : std_logic;
signal \N__24235\ : std_logic;
signal \N__24234\ : std_logic;
signal \N__24231\ : std_logic;
signal \N__24230\ : std_logic;
signal \N__24227\ : std_logic;
signal \N__24224\ : std_logic;
signal \N__24221\ : std_logic;
signal \N__24214\ : std_logic;
signal \N__24211\ : std_logic;
signal \N__24208\ : std_logic;
signal \N__24205\ : std_logic;
signal \N__24202\ : std_logic;
signal \N__24199\ : std_logic;
signal \N__24196\ : std_logic;
signal \N__24195\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24191\ : std_logic;
signal \N__24188\ : std_logic;
signal \N__24185\ : std_logic;
signal \N__24182\ : std_logic;
signal \N__24179\ : std_logic;
signal \N__24176\ : std_logic;
signal \N__24175\ : std_logic;
signal \N__24172\ : std_logic;
signal \N__24167\ : std_logic;
signal \N__24166\ : std_logic;
signal \N__24163\ : std_logic;
signal \N__24160\ : std_logic;
signal \N__24157\ : std_logic;
signal \N__24154\ : std_logic;
signal \N__24151\ : std_logic;
signal \N__24142\ : std_logic;
signal \N__24139\ : std_logic;
signal \N__24138\ : std_logic;
signal \N__24135\ : std_logic;
signal \N__24132\ : std_logic;
signal \N__24129\ : std_logic;
signal \N__24128\ : std_logic;
signal \N__24125\ : std_logic;
signal \N__24122\ : std_logic;
signal \N__24119\ : std_logic;
signal \N__24112\ : std_logic;
signal \N__24111\ : std_logic;
signal \N__24110\ : std_logic;
signal \N__24107\ : std_logic;
signal \N__24102\ : std_logic;
signal \N__24097\ : std_logic;
signal \N__24094\ : std_logic;
signal \N__24091\ : std_logic;
signal \N__24090\ : std_logic;
signal \N__24089\ : std_logic;
signal \N__24086\ : std_logic;
signal \N__24081\ : std_logic;
signal \N__24076\ : std_logic;
signal \N__24073\ : std_logic;
signal \N__24072\ : std_logic;
signal \N__24069\ : std_logic;
signal \N__24066\ : std_logic;
signal \N__24063\ : std_logic;
signal \N__24060\ : std_logic;
signal \N__24055\ : std_logic;
signal \N__24052\ : std_logic;
signal \N__24049\ : std_logic;
signal \N__24046\ : std_logic;
signal \N__24045\ : std_logic;
signal \N__24044\ : std_logic;
signal \N__24041\ : std_logic;
signal \N__24036\ : std_logic;
signal \N__24031\ : std_logic;
signal \N__24030\ : std_logic;
signal \N__24027\ : std_logic;
signal \N__24024\ : std_logic;
signal \N__24021\ : std_logic;
signal \N__24020\ : std_logic;
signal \N__24017\ : std_logic;
signal \N__24014\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24004\ : std_logic;
signal \N__24001\ : std_logic;
signal \N__23998\ : std_logic;
signal \N__23995\ : std_logic;
signal \N__23992\ : std_logic;
signal \N__23989\ : std_logic;
signal \N__23986\ : std_logic;
signal \N__23985\ : std_logic;
signal \N__23982\ : std_logic;
signal \N__23979\ : std_logic;
signal \N__23976\ : std_logic;
signal \N__23973\ : std_logic;
signal \N__23968\ : std_logic;
signal \N__23965\ : std_logic;
signal \N__23962\ : std_logic;
signal \N__23961\ : std_logic;
signal \N__23960\ : std_logic;
signal \N__23957\ : std_logic;
signal \N__23954\ : std_logic;
signal \N__23951\ : std_logic;
signal \N__23946\ : std_logic;
signal \N__23941\ : std_logic;
signal \N__23938\ : std_logic;
signal \N__23935\ : std_logic;
signal \N__23932\ : std_logic;
signal \N__23929\ : std_logic;
signal \N__23926\ : std_logic;
signal \N__23923\ : std_logic;
signal \N__23920\ : std_logic;
signal \N__23917\ : std_logic;
signal \N__23914\ : std_logic;
signal \N__23911\ : std_logic;
signal \N__23908\ : std_logic;
signal \N__23905\ : std_logic;
signal \N__23902\ : std_logic;
signal \N__23899\ : std_logic;
signal \N__23896\ : std_logic;
signal \N__23893\ : std_logic;
signal \N__23890\ : std_logic;
signal \N__23887\ : std_logic;
signal \N__23884\ : std_logic;
signal \N__23881\ : std_logic;
signal \N__23878\ : std_logic;
signal \N__23875\ : std_logic;
signal \N__23874\ : std_logic;
signal \N__23871\ : std_logic;
signal \N__23868\ : std_logic;
signal \N__23865\ : std_logic;
signal \N__23862\ : std_logic;
signal \N__23857\ : std_logic;
signal \N__23856\ : std_logic;
signal \N__23853\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23849\ : std_logic;
signal \N__23846\ : std_logic;
signal \N__23843\ : std_logic;
signal \N__23840\ : std_logic;
signal \N__23837\ : std_logic;
signal \N__23830\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23824\ : std_logic;
signal \N__23823\ : std_logic;
signal \N__23820\ : std_logic;
signal \N__23819\ : std_logic;
signal \N__23816\ : std_logic;
signal \N__23813\ : std_logic;
signal \N__23810\ : std_logic;
signal \N__23807\ : std_logic;
signal \N__23806\ : std_logic;
signal \N__23805\ : std_logic;
signal \N__23800\ : std_logic;
signal \N__23797\ : std_logic;
signal \N__23792\ : std_logic;
signal \N__23785\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23779\ : std_logic;
signal \N__23778\ : std_logic;
signal \N__23777\ : std_logic;
signal \N__23774\ : std_logic;
signal \N__23771\ : std_logic;
signal \N__23768\ : std_logic;
signal \N__23767\ : std_logic;
signal \N__23764\ : std_logic;
signal \N__23763\ : std_logic;
signal \N__23760\ : std_logic;
signal \N__23755\ : std_logic;
signal \N__23752\ : std_logic;
signal \N__23749\ : std_logic;
signal \N__23744\ : std_logic;
signal \N__23737\ : std_logic;
signal \N__23734\ : std_logic;
signal \N__23733\ : std_logic;
signal \N__23732\ : std_logic;
signal \N__23729\ : std_logic;
signal \N__23724\ : std_logic;
signal \N__23719\ : std_logic;
signal \N__23718\ : std_logic;
signal \N__23717\ : std_logic;
signal \N__23714\ : std_logic;
signal \N__23711\ : std_logic;
signal \N__23708\ : std_logic;
signal \N__23701\ : std_logic;
signal \N__23698\ : std_logic;
signal \N__23697\ : std_logic;
signal \N__23694\ : std_logic;
signal \N__23691\ : std_logic;
signal \N__23688\ : std_logic;
signal \N__23683\ : std_logic;
signal \N__23682\ : std_logic;
signal \N__23681\ : std_logic;
signal \N__23680\ : std_logic;
signal \N__23677\ : std_logic;
signal \N__23674\ : std_logic;
signal \N__23671\ : std_logic;
signal \N__23668\ : std_logic;
signal \N__23659\ : std_logic;
signal \N__23656\ : std_logic;
signal \N__23653\ : std_logic;
signal \N__23650\ : std_logic;
signal \N__23647\ : std_logic;
signal \N__23646\ : std_logic;
signal \N__23643\ : std_logic;
signal \N__23640\ : std_logic;
signal \N__23635\ : std_logic;
signal \N__23632\ : std_logic;
signal \N__23629\ : std_logic;
signal \N__23628\ : std_logic;
signal \N__23627\ : std_logic;
signal \N__23624\ : std_logic;
signal \N__23621\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23612\ : std_logic;
signal \N__23609\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23596\ : std_logic;
signal \N__23593\ : std_logic;
signal \N__23590\ : std_logic;
signal \N__23587\ : std_logic;
signal \N__23584\ : std_logic;
signal \N__23581\ : std_logic;
signal \N__23578\ : std_logic;
signal \N__23577\ : std_logic;
signal \N__23574\ : std_logic;
signal \N__23571\ : std_logic;
signal \N__23568\ : std_logic;
signal \N__23565\ : std_logic;
signal \N__23560\ : std_logic;
signal \N__23557\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23553\ : std_logic;
signal \N__23550\ : std_logic;
signal \N__23547\ : std_logic;
signal \N__23542\ : std_logic;
signal \N__23541\ : std_logic;
signal \N__23538\ : std_logic;
signal \N__23535\ : std_logic;
signal \N__23532\ : std_logic;
signal \N__23529\ : std_logic;
signal \N__23524\ : std_logic;
signal \N__23523\ : std_logic;
signal \N__23520\ : std_logic;
signal \N__23517\ : std_logic;
signal \N__23514\ : std_logic;
signal \N__23511\ : std_logic;
signal \N__23508\ : std_logic;
signal \N__23505\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23499\ : std_logic;
signal \N__23496\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23490\ : std_logic;
signal \N__23487\ : std_logic;
signal \N__23482\ : std_logic;
signal \N__23479\ : std_logic;
signal \N__23478\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23474\ : std_logic;
signal \N__23471\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23463\ : std_logic;
signal \N__23458\ : std_logic;
signal \N__23457\ : std_logic;
signal \N__23454\ : std_logic;
signal \N__23451\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23444\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23436\ : std_logic;
signal \N__23431\ : std_logic;
signal \N__23428\ : std_logic;
signal \N__23425\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23419\ : std_logic;
signal \N__23416\ : std_logic;
signal \N__23415\ : std_logic;
signal \N__23412\ : std_logic;
signal \N__23409\ : std_logic;
signal \N__23404\ : std_logic;
signal \N__23401\ : std_logic;
signal \N__23398\ : std_logic;
signal \N__23395\ : std_logic;
signal \N__23392\ : std_logic;
signal \N__23391\ : std_logic;
signal \N__23388\ : std_logic;
signal \N__23385\ : std_logic;
signal \N__23382\ : std_logic;
signal \N__23379\ : std_logic;
signal \N__23374\ : std_logic;
signal \N__23371\ : std_logic;
signal \N__23368\ : std_logic;
signal \N__23367\ : std_logic;
signal \N__23364\ : std_logic;
signal \N__23361\ : std_logic;
signal \N__23358\ : std_logic;
signal \N__23355\ : std_logic;
signal \N__23350\ : std_logic;
signal \N__23347\ : std_logic;
signal \N__23344\ : std_logic;
signal \N__23343\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23337\ : std_logic;
signal \N__23334\ : std_logic;
signal \N__23331\ : std_logic;
signal \N__23326\ : std_logic;
signal \N__23325\ : std_logic;
signal \N__23322\ : std_logic;
signal \N__23319\ : std_logic;
signal \N__23316\ : std_logic;
signal \N__23313\ : std_logic;
signal \N__23308\ : std_logic;
signal \N__23307\ : std_logic;
signal \N__23304\ : std_logic;
signal \N__23301\ : std_logic;
signal \N__23298\ : std_logic;
signal \N__23295\ : std_logic;
signal \N__23290\ : std_logic;
signal \N__23287\ : std_logic;
signal \N__23286\ : std_logic;
signal \N__23283\ : std_logic;
signal \N__23280\ : std_logic;
signal \N__23277\ : std_logic;
signal \N__23274\ : std_logic;
signal \N__23269\ : std_logic;
signal \N__23266\ : std_logic;
signal \N__23263\ : std_logic;
signal \N__23260\ : std_logic;
signal \N__23257\ : std_logic;
signal \N__23254\ : std_logic;
signal \N__23251\ : std_logic;
signal \N__23248\ : std_logic;
signal \N__23245\ : std_logic;
signal \N__23242\ : std_logic;
signal \N__23239\ : std_logic;
signal \N__23236\ : std_logic;
signal \N__23233\ : std_logic;
signal \N__23232\ : std_logic;
signal \N__23231\ : std_logic;
signal \N__23230\ : std_logic;
signal \N__23229\ : std_logic;
signal \N__23226\ : std_logic;
signal \N__23219\ : std_logic;
signal \N__23216\ : std_logic;
signal \N__23209\ : std_logic;
signal \N__23206\ : std_logic;
signal \N__23205\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23199\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23191\ : std_logic;
signal \N__23188\ : std_logic;
signal \N__23185\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23179\ : std_logic;
signal \N__23176\ : std_logic;
signal \N__23173\ : std_logic;
signal \N__23172\ : std_logic;
signal \N__23169\ : std_logic;
signal \N__23166\ : std_logic;
signal \N__23163\ : std_logic;
signal \N__23160\ : std_logic;
signal \N__23155\ : std_logic;
signal \N__23152\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23146\ : std_logic;
signal \N__23143\ : std_logic;
signal \N__23140\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23134\ : std_logic;
signal \N__23133\ : std_logic;
signal \N__23130\ : std_logic;
signal \N__23127\ : std_logic;
signal \N__23122\ : std_logic;
signal \N__23119\ : std_logic;
signal \N__23118\ : std_logic;
signal \N__23115\ : std_logic;
signal \N__23112\ : std_logic;
signal \N__23107\ : std_logic;
signal \N__23104\ : std_logic;
signal \N__23103\ : std_logic;
signal \N__23100\ : std_logic;
signal \N__23097\ : std_logic;
signal \N__23094\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23086\ : std_logic;
signal \N__23085\ : std_logic;
signal \N__23082\ : std_logic;
signal \N__23079\ : std_logic;
signal \N__23074\ : std_logic;
signal \N__23071\ : std_logic;
signal \N__23070\ : std_logic;
signal \N__23067\ : std_logic;
signal \N__23064\ : std_logic;
signal \N__23059\ : std_logic;
signal \N__23056\ : std_logic;
signal \N__23053\ : std_logic;
signal \N__23052\ : std_logic;
signal \N__23049\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23041\ : std_logic;
signal \N__23038\ : std_logic;
signal \N__23035\ : std_logic;
signal \N__23032\ : std_logic;
signal \N__23029\ : std_logic;
signal \N__23026\ : std_logic;
signal \N__23023\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23017\ : std_logic;
signal \N__23014\ : std_logic;
signal \N__23011\ : std_logic;
signal \N__23008\ : std_logic;
signal \N__23005\ : std_logic;
signal \N__23002\ : std_logic;
signal \N__22999\ : std_logic;
signal \N__22998\ : std_logic;
signal \N__22995\ : std_logic;
signal \N__22994\ : std_logic;
signal \N__22993\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22983\ : std_logic;
signal \N__22982\ : std_logic;
signal \N__22977\ : std_logic;
signal \N__22974\ : std_logic;
signal \N__22971\ : std_logic;
signal \N__22968\ : std_logic;
signal \N__22965\ : std_logic;
signal \N__22962\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22951\ : std_logic;
signal \N__22948\ : std_logic;
signal \N__22945\ : std_logic;
signal \N__22942\ : std_logic;
signal \N__22941\ : std_logic;
signal \N__22938\ : std_logic;
signal \N__22935\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22926\ : std_logic;
signal \N__22923\ : std_logic;
signal \N__22920\ : std_logic;
signal \N__22917\ : std_logic;
signal \N__22912\ : std_logic;
signal \N__22909\ : std_logic;
signal \N__22906\ : std_logic;
signal \N__22905\ : std_logic;
signal \N__22900\ : std_logic;
signal \N__22897\ : std_logic;
signal \N__22896\ : std_logic;
signal \N__22891\ : std_logic;
signal \N__22888\ : std_logic;
signal \N__22887\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22879\ : std_logic;
signal \N__22876\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22872\ : std_logic;
signal \N__22869\ : std_logic;
signal \N__22864\ : std_logic;
signal \N__22861\ : std_logic;
signal \N__22858\ : std_logic;
signal \N__22855\ : std_logic;
signal \N__22852\ : std_logic;
signal \N__22849\ : std_logic;
signal \N__22846\ : std_logic;
signal \N__22845\ : std_logic;
signal \N__22842\ : std_logic;
signal \N__22839\ : std_logic;
signal \N__22838\ : std_logic;
signal \N__22835\ : std_logic;
signal \N__22830\ : std_logic;
signal \N__22825\ : std_logic;
signal \N__22822\ : std_logic;
signal \N__22819\ : std_logic;
signal \N__22818\ : std_logic;
signal \N__22815\ : std_logic;
signal \N__22812\ : std_logic;
signal \N__22807\ : std_logic;
signal \N__22804\ : std_logic;
signal \N__22803\ : std_logic;
signal \N__22800\ : std_logic;
signal \N__22797\ : std_logic;
signal \N__22796\ : std_logic;
signal \N__22793\ : std_logic;
signal \N__22788\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22782\ : std_logic;
signal \N__22779\ : std_logic;
signal \N__22776\ : std_logic;
signal \N__22775\ : std_logic;
signal \N__22768\ : std_logic;
signal \N__22765\ : std_logic;
signal \N__22762\ : std_logic;
signal \N__22759\ : std_logic;
signal \N__22756\ : std_logic;
signal \N__22753\ : std_logic;
signal \N__22750\ : std_logic;
signal \N__22747\ : std_logic;
signal \N__22744\ : std_logic;
signal \N__22741\ : std_logic;
signal \N__22740\ : std_logic;
signal \N__22739\ : std_logic;
signal \N__22734\ : std_logic;
signal \N__22731\ : std_logic;
signal \N__22726\ : std_logic;
signal \N__22725\ : std_logic;
signal \N__22724\ : std_logic;
signal \N__22721\ : std_logic;
signal \N__22716\ : std_logic;
signal \N__22711\ : std_logic;
signal \N__22708\ : std_logic;
signal \N__22705\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22703\ : std_logic;
signal \N__22700\ : std_logic;
signal \N__22697\ : std_logic;
signal \N__22694\ : std_logic;
signal \N__22691\ : std_logic;
signal \N__22688\ : std_logic;
signal \N__22681\ : std_logic;
signal \N__22678\ : std_logic;
signal \N__22677\ : std_logic;
signal \N__22674\ : std_logic;
signal \N__22673\ : std_logic;
signal \N__22670\ : std_logic;
signal \N__22667\ : std_logic;
signal \N__22664\ : std_logic;
signal \N__22657\ : std_logic;
signal \N__22656\ : std_logic;
signal \N__22653\ : std_logic;
signal \N__22652\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22643\ : std_logic;
signal \N__22640\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22634\ : std_logic;
signal \N__22627\ : std_logic;
signal \N__22626\ : std_logic;
signal \N__22623\ : std_logic;
signal \N__22620\ : std_logic;
signal \N__22619\ : std_logic;
signal \N__22614\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22606\ : std_logic;
signal \N__22605\ : std_logic;
signal \N__22600\ : std_logic;
signal \N__22597\ : std_logic;
signal \N__22596\ : std_logic;
signal \N__22595\ : std_logic;
signal \N__22592\ : std_logic;
signal \N__22589\ : std_logic;
signal \N__22586\ : std_logic;
signal \N__22583\ : std_logic;
signal \N__22580\ : std_logic;
signal \N__22577\ : std_logic;
signal \N__22570\ : std_logic;
signal \N__22567\ : std_logic;
signal \N__22566\ : std_logic;
signal \N__22563\ : std_logic;
signal \N__22560\ : std_logic;
signal \N__22559\ : std_logic;
signal \N__22556\ : std_logic;
signal \N__22553\ : std_logic;
signal \N__22550\ : std_logic;
signal \N__22543\ : std_logic;
signal \N__22540\ : std_logic;
signal \N__22537\ : std_logic;
signal \N__22534\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22522\ : std_logic;
signal \N__22519\ : std_logic;
signal \N__22518\ : std_logic;
signal \N__22515\ : std_logic;
signal \N__22512\ : std_logic;
signal \N__22509\ : std_logic;
signal \N__22506\ : std_logic;
signal \N__22501\ : std_logic;
signal \N__22498\ : std_logic;
signal \N__22495\ : std_logic;
signal \N__22492\ : std_logic;
signal \N__22491\ : std_logic;
signal \N__22490\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22484\ : std_logic;
signal \N__22481\ : std_logic;
signal \N__22478\ : std_logic;
signal \N__22475\ : std_logic;
signal \N__22468\ : std_logic;
signal \N__22465\ : std_logic;
signal \N__22462\ : std_logic;
signal \N__22459\ : std_logic;
signal \N__22456\ : std_logic;
signal \N__22453\ : std_logic;
signal \N__22452\ : std_logic;
signal \N__22449\ : std_logic;
signal \N__22446\ : std_logic;
signal \N__22443\ : std_logic;
signal \N__22440\ : std_logic;
signal \N__22435\ : std_logic;
signal \N__22432\ : std_logic;
signal \N__22429\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22425\ : std_logic;
signal \N__22424\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22416\ : std_logic;
signal \N__22411\ : std_logic;
signal \N__22410\ : std_logic;
signal \N__22409\ : std_logic;
signal \N__22408\ : std_logic;
signal \N__22405\ : std_logic;
signal \N__22404\ : std_logic;
signal \N__22403\ : std_logic;
signal \N__22402\ : std_logic;
signal \N__22399\ : std_logic;
signal \N__22396\ : std_logic;
signal \N__22395\ : std_logic;
signal \N__22394\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22390\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22388\ : std_logic;
signal \N__22387\ : std_logic;
signal \N__22384\ : std_logic;
signal \N__22381\ : std_logic;
signal \N__22378\ : std_logic;
signal \N__22375\ : std_logic;
signal \N__22362\ : std_logic;
signal \N__22361\ : std_logic;
signal \N__22360\ : std_logic;
signal \N__22359\ : std_logic;
signal \N__22356\ : std_logic;
signal \N__22355\ : std_logic;
signal \N__22354\ : std_logic;
signal \N__22353\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22351\ : std_logic;
signal \N__22350\ : std_logic;
signal \N__22345\ : std_logic;
signal \N__22342\ : std_logic;
signal \N__22337\ : std_logic;
signal \N__22334\ : std_logic;
signal \N__22333\ : std_logic;
signal \N__22330\ : std_logic;
signal \N__22325\ : std_logic;
signal \N__22324\ : std_logic;
signal \N__22323\ : std_logic;
signal \N__22316\ : std_logic;
signal \N__22313\ : std_logic;
signal \N__22310\ : std_logic;
signal \N__22303\ : std_logic;
signal \N__22294\ : std_logic;
signal \N__22291\ : std_logic;
signal \N__22286\ : std_logic;
signal \N__22281\ : std_logic;
signal \N__22278\ : std_logic;
signal \N__22261\ : std_logic;
signal \N__22260\ : std_logic;
signal \N__22259\ : std_logic;
signal \N__22258\ : std_logic;
signal \N__22257\ : std_logic;
signal \N__22256\ : std_logic;
signal \N__22255\ : std_logic;
signal \N__22254\ : std_logic;
signal \N__22253\ : std_logic;
signal \N__22252\ : std_logic;
signal \N__22249\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22246\ : std_logic;
signal \N__22243\ : std_logic;
signal \N__22240\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22224\ : std_logic;
signal \N__22223\ : std_logic;
signal \N__22222\ : std_logic;
signal \N__22221\ : std_logic;
signal \N__22220\ : std_logic;
signal \N__22219\ : std_logic;
signal \N__22212\ : std_logic;
signal \N__22209\ : std_logic;
signal \N__22204\ : std_logic;
signal \N__22199\ : std_logic;
signal \N__22196\ : std_logic;
signal \N__22195\ : std_logic;
signal \N__22194\ : std_logic;
signal \N__22193\ : std_logic;
signal \N__22192\ : std_logic;
signal \N__22191\ : std_logic;
signal \N__22190\ : std_logic;
signal \N__22187\ : std_logic;
signal \N__22182\ : std_logic;
signal \N__22179\ : std_logic;
signal \N__22176\ : std_logic;
signal \N__22169\ : std_logic;
signal \N__22166\ : std_logic;
signal \N__22163\ : std_logic;
signal \N__22158\ : std_logic;
signal \N__22151\ : std_logic;
signal \N__22132\ : std_logic;
signal \N__22131\ : std_logic;
signal \N__22130\ : std_logic;
signal \N__22129\ : std_logic;
signal \N__22128\ : std_logic;
signal \N__22127\ : std_logic;
signal \N__22126\ : std_logic;
signal \N__22125\ : std_logic;
signal \N__22124\ : std_logic;
signal \N__22123\ : std_logic;
signal \N__22122\ : std_logic;
signal \N__22121\ : std_logic;
signal \N__22120\ : std_logic;
signal \N__22119\ : std_logic;
signal \N__22118\ : std_logic;
signal \N__22117\ : std_logic;
signal \N__22116\ : std_logic;
signal \N__22115\ : std_logic;
signal \N__22114\ : std_logic;
signal \N__22113\ : std_logic;
signal \N__22110\ : std_logic;
signal \N__22109\ : std_logic;
signal \N__22106\ : std_logic;
signal \N__22105\ : std_logic;
signal \N__22104\ : std_logic;
signal \N__22103\ : std_logic;
signal \N__22102\ : std_logic;
signal \N__22101\ : std_logic;
signal \N__22100\ : std_logic;
signal \N__22099\ : std_logic;
signal \N__22096\ : std_logic;
signal \N__22095\ : std_logic;
signal \N__22094\ : std_logic;
signal \N__22093\ : std_logic;
signal \N__22088\ : std_logic;
signal \N__22085\ : std_logic;
signal \N__22076\ : std_logic;
signal \N__22069\ : std_logic;
signal \N__22064\ : std_logic;
signal \N__22057\ : std_logic;
signal \N__22044\ : std_logic;
signal \N__22041\ : std_logic;
signal \N__22038\ : std_logic;
signal \N__22037\ : std_logic;
signal \N__22036\ : std_logic;
signal \N__22035\ : std_logic;
signal \N__22034\ : std_logic;
signal \N__22033\ : std_logic;
signal \N__22032\ : std_logic;
signal \N__22031\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22027\ : std_logic;
signal \N__22026\ : std_logic;
signal \N__22025\ : std_logic;
signal \N__22018\ : std_logic;
signal \N__22015\ : std_logic;
signal \N__22008\ : std_logic;
signal \N__21999\ : std_logic;
signal \N__21992\ : std_logic;
signal \N__21991\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21989\ : std_logic;
signal \N__21984\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21968\ : std_logic;
signal \N__21965\ : std_logic;
signal \N__21962\ : std_logic;
signal \N__21959\ : std_logic;
signal \N__21956\ : std_logic;
signal \N__21953\ : std_logic;
signal \N__21944\ : std_logic;
signal \N__21937\ : std_logic;
signal \N__21934\ : std_logic;
signal \N__21931\ : std_logic;
signal \N__21910\ : std_logic;
signal \N__21907\ : std_logic;
signal \N__21904\ : std_logic;
signal \N__21903\ : std_logic;
signal \N__21900\ : std_logic;
signal \N__21897\ : std_logic;
signal \N__21892\ : std_logic;
signal \N__21889\ : std_logic;
signal \N__21886\ : std_logic;
signal \N__21883\ : std_logic;
signal \N__21880\ : std_logic;
signal \N__21877\ : std_logic;
signal \N__21874\ : std_logic;
signal \N__21871\ : std_logic;
signal \N__21868\ : std_logic;
signal \N__21867\ : std_logic;
signal \N__21864\ : std_logic;
signal \N__21861\ : std_logic;
signal \N__21856\ : std_logic;
signal \N__21853\ : std_logic;
signal \N__21852\ : std_logic;
signal \N__21849\ : std_logic;
signal \N__21846\ : std_logic;
signal \N__21843\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21839\ : std_logic;
signal \N__21834\ : std_logic;
signal \N__21831\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21823\ : std_logic;
signal \N__21820\ : std_logic;
signal \N__21817\ : std_logic;
signal \N__21814\ : std_logic;
signal \N__21813\ : std_logic;
signal \N__21810\ : std_logic;
signal \N__21807\ : std_logic;
signal \N__21802\ : std_logic;
signal \N__21801\ : std_logic;
signal \N__21798\ : std_logic;
signal \N__21795\ : std_logic;
signal \N__21794\ : std_logic;
signal \N__21791\ : std_logic;
signal \N__21786\ : std_logic;
signal \N__21781\ : std_logic;
signal \N__21778\ : std_logic;
signal \N__21777\ : std_logic;
signal \N__21776\ : std_logic;
signal \N__21773\ : std_logic;
signal \N__21770\ : std_logic;
signal \N__21767\ : std_logic;
signal \N__21760\ : std_logic;
signal \N__21759\ : std_logic;
signal \N__21756\ : std_logic;
signal \N__21753\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21746\ : std_logic;
signal \N__21743\ : std_logic;
signal \N__21736\ : std_logic;
signal \N__21733\ : std_logic;
signal \N__21732\ : std_logic;
signal \N__21729\ : std_logic;
signal \N__21726\ : std_logic;
signal \N__21725\ : std_logic;
signal \N__21722\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21716\ : std_logic;
signal \N__21709\ : std_logic;
signal \N__21706\ : std_logic;
signal \N__21703\ : std_logic;
signal \N__21700\ : std_logic;
signal \N__21697\ : std_logic;
signal \N__21696\ : std_logic;
signal \N__21695\ : std_logic;
signal \N__21692\ : std_logic;
signal \N__21687\ : std_logic;
signal \N__21684\ : std_logic;
signal \N__21681\ : std_logic;
signal \N__21676\ : std_logic;
signal \N__21673\ : std_logic;
signal \N__21672\ : std_logic;
signal \N__21671\ : std_logic;
signal \N__21668\ : std_logic;
signal \N__21665\ : std_logic;
signal \N__21662\ : std_logic;
signal \N__21659\ : std_logic;
signal \N__21656\ : std_logic;
signal \N__21649\ : std_logic;
signal \N__21646\ : std_logic;
signal \N__21643\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21637\ : std_logic;
signal \N__21634\ : std_logic;
signal \N__21631\ : std_logic;
signal \N__21628\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21619\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21610\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21604\ : std_logic;
signal \N__21603\ : std_logic;
signal \N__21600\ : std_logic;
signal \N__21597\ : std_logic;
signal \N__21594\ : std_logic;
signal \N__21591\ : std_logic;
signal \N__21586\ : std_logic;
signal \N__21583\ : std_logic;
signal \N__21580\ : std_logic;
signal \N__21579\ : std_logic;
signal \N__21576\ : std_logic;
signal \N__21573\ : std_logic;
signal \N__21568\ : std_logic;
signal \N__21567\ : std_logic;
signal \N__21564\ : std_logic;
signal \N__21561\ : std_logic;
signal \N__21558\ : std_logic;
signal \N__21557\ : std_logic;
signal \N__21554\ : std_logic;
signal \N__21551\ : std_logic;
signal \N__21548\ : std_logic;
signal \N__21541\ : std_logic;
signal \N__21540\ : std_logic;
signal \N__21537\ : std_logic;
signal \N__21534\ : std_logic;
signal \N__21533\ : std_logic;
signal \N__21530\ : std_logic;
signal \N__21527\ : std_logic;
signal \N__21524\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21514\ : std_logic;
signal \N__21513\ : std_logic;
signal \N__21510\ : std_logic;
signal \N__21507\ : std_logic;
signal \N__21502\ : std_logic;
signal \N__21501\ : std_logic;
signal \N__21496\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21490\ : std_logic;
signal \N__21487\ : std_logic;
signal \N__21484\ : std_logic;
signal \N__21481\ : std_logic;
signal \N__21478\ : std_logic;
signal \N__21475\ : std_logic;
signal \N__21474\ : std_logic;
signal \N__21473\ : std_logic;
signal \N__21470\ : std_logic;
signal \N__21467\ : std_logic;
signal \N__21464\ : std_logic;
signal \N__21461\ : std_logic;
signal \N__21458\ : std_logic;
signal \N__21451\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21447\ : std_logic;
signal \N__21446\ : std_logic;
signal \N__21443\ : std_logic;
signal \N__21440\ : std_logic;
signal \N__21437\ : std_logic;
signal \N__21434\ : std_logic;
signal \N__21431\ : std_logic;
signal \N__21428\ : std_logic;
signal \N__21421\ : std_logic;
signal \N__21420\ : std_logic;
signal \N__21417\ : std_logic;
signal \N__21414\ : std_logic;
signal \N__21413\ : std_logic;
signal \N__21406\ : std_logic;
signal \N__21403\ : std_logic;
signal \N__21400\ : std_logic;
signal \N__21397\ : std_logic;
signal \N__21394\ : std_logic;
signal \N__21391\ : std_logic;
signal \N__21388\ : std_logic;
signal \N__21387\ : std_logic;
signal \N__21386\ : std_logic;
signal \N__21383\ : std_logic;
signal \N__21378\ : std_logic;
signal \N__21373\ : std_logic;
signal \N__21370\ : std_logic;
signal \N__21367\ : std_logic;
signal \N__21366\ : std_logic;
signal \N__21363\ : std_logic;
signal \N__21360\ : std_logic;
signal \N__21357\ : std_logic;
signal \N__21354\ : std_logic;
signal \N__21349\ : std_logic;
signal \N__21346\ : std_logic;
signal \N__21345\ : std_logic;
signal \N__21342\ : std_logic;
signal \N__21339\ : std_logic;
signal \N__21338\ : std_logic;
signal \N__21335\ : std_logic;
signal \N__21332\ : std_logic;
signal \N__21329\ : std_logic;
signal \N__21322\ : std_logic;
signal \N__21321\ : std_logic;
signal \N__21318\ : std_logic;
signal \N__21315\ : std_logic;
signal \N__21314\ : std_logic;
signal \N__21311\ : std_logic;
signal \N__21308\ : std_logic;
signal \N__21305\ : std_logic;
signal \N__21298\ : std_logic;
signal \N__21297\ : std_logic;
signal \N__21294\ : std_logic;
signal \N__21291\ : std_logic;
signal \N__21290\ : std_logic;
signal \N__21287\ : std_logic;
signal \N__21282\ : std_logic;
signal \N__21277\ : std_logic;
signal \N__21276\ : std_logic;
signal \N__21273\ : std_logic;
signal \N__21270\ : std_logic;
signal \N__21269\ : std_logic;
signal \N__21266\ : std_logic;
signal \N__21263\ : std_logic;
signal \N__21260\ : std_logic;
signal \N__21253\ : std_logic;
signal \N__21252\ : std_logic;
signal \N__21251\ : std_logic;
signal \N__21246\ : std_logic;
signal \N__21243\ : std_logic;
signal \N__21238\ : std_logic;
signal \N__21237\ : std_logic;
signal \N__21234\ : std_logic;
signal \N__21231\ : std_logic;
signal \N__21230\ : std_logic;
signal \N__21227\ : std_logic;
signal \N__21224\ : std_logic;
signal \N__21221\ : std_logic;
signal \N__21214\ : std_logic;
signal \N__21213\ : std_logic;
signal \N__21210\ : std_logic;
signal \N__21207\ : std_logic;
signal \N__21202\ : std_logic;
signal \N__21199\ : std_logic;
signal \N__21196\ : std_logic;
signal \N__21195\ : std_logic;
signal \N__21190\ : std_logic;
signal \N__21187\ : std_logic;
signal \N__21186\ : std_logic;
signal \N__21185\ : std_logic;
signal \N__21184\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21182\ : std_logic;
signal \N__21181\ : std_logic;
signal \N__21170\ : std_logic;
signal \N__21165\ : std_logic;
signal \N__21160\ : std_logic;
signal \N__21159\ : std_logic;
signal \N__21158\ : std_logic;
signal \N__21157\ : std_logic;
signal \N__21156\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21154\ : std_logic;
signal \N__21153\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21149\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21141\ : std_logic;
signal \N__21134\ : std_logic;
signal \N__21131\ : std_logic;
signal \N__21128\ : std_logic;
signal \N__21115\ : std_logic;
signal \N__21114\ : std_logic;
signal \N__21111\ : std_logic;
signal \N__21108\ : std_logic;
signal \N__21103\ : std_logic;
signal \N__21100\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21096\ : std_logic;
signal \N__21093\ : std_logic;
signal \N__21090\ : std_logic;
signal \N__21087\ : std_logic;
signal \N__21084\ : std_logic;
signal \N__21079\ : std_logic;
signal \N__21076\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21070\ : std_logic;
signal \N__21069\ : std_logic;
signal \N__21066\ : std_logic;
signal \N__21065\ : std_logic;
signal \N__21062\ : std_logic;
signal \N__21059\ : std_logic;
signal \N__21056\ : std_logic;
signal \N__21049\ : std_logic;
signal \N__21046\ : std_logic;
signal \N__21043\ : std_logic;
signal \N__21042\ : std_logic;
signal \N__21039\ : std_logic;
signal \N__21038\ : std_logic;
signal \N__21035\ : std_logic;
signal \N__21032\ : std_logic;
signal \N__21029\ : std_logic;
signal \N__21022\ : std_logic;
signal \N__21019\ : std_logic;
signal \N__21016\ : std_logic;
signal \N__21013\ : std_logic;
signal \N__21010\ : std_logic;
signal \N__21007\ : std_logic;
signal \N__21004\ : std_logic;
signal \N__21001\ : std_logic;
signal \N__20998\ : std_logic;
signal \N__20995\ : std_logic;
signal \N__20994\ : std_logic;
signal \N__20991\ : std_logic;
signal \N__20988\ : std_logic;
signal \N__20983\ : std_logic;
signal \N__20980\ : std_logic;
signal \N__20977\ : std_logic;
signal \N__20974\ : std_logic;
signal \N__20971\ : std_logic;
signal \N__20970\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20968\ : std_logic;
signal \N__20967\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20965\ : std_logic;
signal \N__20964\ : std_logic;
signal \N__20963\ : std_logic;
signal \N__20960\ : std_logic;
signal \N__20949\ : std_logic;
signal \N__20946\ : std_logic;
signal \N__20945\ : std_logic;
signal \N__20944\ : std_logic;
signal \N__20943\ : std_logic;
signal \N__20942\ : std_logic;
signal \N__20941\ : std_logic;
signal \N__20940\ : std_logic;
signal \N__20939\ : std_logic;
signal \N__20938\ : std_logic;
signal \N__20937\ : std_logic;
signal \N__20936\ : std_logic;
signal \N__20935\ : std_logic;
signal \N__20934\ : std_logic;
signal \N__20933\ : std_logic;
signal \N__20932\ : std_logic;
signal \N__20929\ : std_logic;
signal \N__20928\ : std_logic;
signal \N__20927\ : std_logic;
signal \N__20926\ : std_logic;
signal \N__20925\ : std_logic;
signal \N__20924\ : std_logic;
signal \N__20923\ : std_logic;
signal \N__20920\ : std_logic;
signal \N__20915\ : std_logic;
signal \N__20914\ : std_logic;
signal \N__20913\ : std_logic;
signal \N__20910\ : std_logic;
signal \N__20907\ : std_logic;
signal \N__20898\ : std_logic;
signal \N__20897\ : std_logic;
signal \N__20896\ : std_logic;
signal \N__20895\ : std_logic;
signal \N__20894\ : std_logic;
signal \N__20893\ : std_logic;
signal \N__20890\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20870\ : std_logic;
signal \N__20867\ : std_logic;
signal \N__20856\ : std_logic;
signal \N__20851\ : std_logic;
signal \N__20846\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20828\ : std_logic;
signal \N__20809\ : std_logic;
signal \N__20806\ : std_logic;
signal \N__20805\ : std_logic;
signal \N__20800\ : std_logic;
signal \N__20797\ : std_logic;
signal \N__20794\ : std_logic;
signal \N__20791\ : std_logic;
signal \N__20790\ : std_logic;
signal \N__20787\ : std_logic;
signal \N__20784\ : std_logic;
signal \N__20779\ : std_logic;
signal \N__20776\ : std_logic;
signal \N__20773\ : std_logic;
signal \N__20770\ : std_logic;
signal \N__20767\ : std_logic;
signal \N__20764\ : std_logic;
signal \N__20761\ : std_logic;
signal \N__20758\ : std_logic;
signal \N__20755\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20746\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20740\ : std_logic;
signal \N__20737\ : std_logic;
signal \N__20734\ : std_logic;
signal \N__20731\ : std_logic;
signal \N__20730\ : std_logic;
signal \N__20727\ : std_logic;
signal \N__20724\ : std_logic;
signal \N__20719\ : std_logic;
signal \N__20716\ : std_logic;
signal \N__20713\ : std_logic;
signal \N__20710\ : std_logic;
signal \N__20707\ : std_logic;
signal \N__20704\ : std_logic;
signal \N__20701\ : std_logic;
signal \N__20698\ : std_logic;
signal \N__20695\ : std_logic;
signal \N__20692\ : std_logic;
signal \N__20689\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20683\ : std_logic;
signal \N__20680\ : std_logic;
signal \N__20679\ : std_logic;
signal \N__20676\ : std_logic;
signal \N__20673\ : std_logic;
signal \N__20668\ : std_logic;
signal \N__20665\ : std_logic;
signal \N__20662\ : std_logic;
signal \N__20659\ : std_logic;
signal \N__20656\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20641\ : std_logic;
signal \N__20640\ : std_logic;
signal \N__20637\ : std_logic;
signal \N__20634\ : std_logic;
signal \N__20631\ : std_logic;
signal \N__20628\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20620\ : std_logic;
signal \N__20617\ : std_logic;
signal \N__20616\ : std_logic;
signal \N__20615\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20606\ : std_logic;
signal \N__20603\ : std_logic;
signal \N__20596\ : std_logic;
signal \N__20595\ : std_logic;
signal \N__20592\ : std_logic;
signal \N__20589\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20586\ : std_logic;
signal \N__20583\ : std_logic;
signal \N__20576\ : std_logic;
signal \N__20573\ : std_logic;
signal \N__20566\ : std_logic;
signal \N__20563\ : std_logic;
signal \N__20562\ : std_logic;
signal \N__20561\ : std_logic;
signal \N__20558\ : std_logic;
signal \N__20555\ : std_logic;
signal \N__20552\ : std_logic;
signal \N__20545\ : std_logic;
signal \N__20544\ : std_logic;
signal \N__20541\ : std_logic;
signal \N__20540\ : std_logic;
signal \N__20537\ : std_logic;
signal \N__20534\ : std_logic;
signal \N__20531\ : std_logic;
signal \N__20524\ : std_logic;
signal \N__20521\ : std_logic;
signal \N__20520\ : std_logic;
signal \N__20519\ : std_logic;
signal \N__20518\ : std_logic;
signal \N__20517\ : std_logic;
signal \N__20514\ : std_logic;
signal \N__20511\ : std_logic;
signal \N__20508\ : std_logic;
signal \N__20505\ : std_logic;
signal \N__20502\ : std_logic;
signal \N__20493\ : std_logic;
signal \N__20490\ : std_logic;
signal \N__20487\ : std_logic;
signal \N__20482\ : std_logic;
signal \N__20479\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20475\ : std_logic;
signal \N__20472\ : std_logic;
signal \N__20469\ : std_logic;
signal \N__20466\ : std_logic;
signal \N__20461\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20457\ : std_logic;
signal \N__20454\ : std_logic;
signal \N__20453\ : std_logic;
signal \N__20450\ : std_logic;
signal \N__20449\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20439\ : std_logic;
signal \N__20436\ : std_logic;
signal \N__20431\ : std_logic;
signal \N__20430\ : std_logic;
signal \N__20429\ : std_logic;
signal \N__20426\ : std_logic;
signal \N__20421\ : std_logic;
signal \N__20418\ : std_logic;
signal \N__20413\ : std_logic;
signal \N__20410\ : std_logic;
signal \N__20407\ : std_logic;
signal \N__20404\ : std_logic;
signal \N__20401\ : std_logic;
signal \N__20398\ : std_logic;
signal \N__20395\ : std_logic;
signal \N__20392\ : std_logic;
signal \N__20389\ : std_logic;
signal \N__20386\ : std_logic;
signal \N__20383\ : std_logic;
signal \N__20380\ : std_logic;
signal \N__20377\ : std_logic;
signal \N__20374\ : std_logic;
signal \N__20371\ : std_logic;
signal \N__20368\ : std_logic;
signal \N__20367\ : std_logic;
signal \N__20364\ : std_logic;
signal \N__20361\ : std_logic;
signal \N__20358\ : std_logic;
signal \N__20355\ : std_logic;
signal \N__20352\ : std_logic;
signal \N__20349\ : std_logic;
signal \N__20346\ : std_logic;
signal \N__20343\ : std_logic;
signal \N__20340\ : std_logic;
signal \N__20337\ : std_logic;
signal \N__20334\ : std_logic;
signal \N__20331\ : std_logic;
signal \N__20328\ : std_logic;
signal \N__20325\ : std_logic;
signal \N__20322\ : std_logic;
signal \N__20319\ : std_logic;
signal \N__20316\ : std_logic;
signal \N__20313\ : std_logic;
signal \N__20310\ : std_logic;
signal \N__20305\ : std_logic;
signal \N__20304\ : std_logic;
signal \N__20301\ : std_logic;
signal \N__20300\ : std_logic;
signal \N__20293\ : std_logic;
signal \N__20290\ : std_logic;
signal \N__20287\ : std_logic;
signal \N__20284\ : std_logic;
signal \N__20281\ : std_logic;
signal \N__20280\ : std_logic;
signal \N__20277\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20271\ : std_logic;
signal \N__20268\ : std_logic;
signal \N__20263\ : std_logic;
signal \N__20260\ : std_logic;
signal \N__20257\ : std_logic;
signal \N__20254\ : std_logic;
signal \N__20251\ : std_logic;
signal \N__20248\ : std_logic;
signal \N__20245\ : std_logic;
signal \N__20244\ : std_logic;
signal \N__20241\ : std_logic;
signal \N__20238\ : std_logic;
signal \N__20235\ : std_logic;
signal \N__20232\ : std_logic;
signal \N__20227\ : std_logic;
signal \N__20224\ : std_logic;
signal \N__20221\ : std_logic;
signal \N__20218\ : std_logic;
signal \N__20217\ : std_logic;
signal \N__20214\ : std_logic;
signal \N__20211\ : std_logic;
signal \N__20208\ : std_logic;
signal \N__20205\ : std_logic;
signal \N__20200\ : std_logic;
signal \N__20197\ : std_logic;
signal \N__20194\ : std_logic;
signal \N__20191\ : std_logic;
signal \N__20190\ : std_logic;
signal \N__20189\ : std_logic;
signal \N__20186\ : std_logic;
signal \N__20181\ : std_logic;
signal \N__20176\ : std_logic;
signal \N__20173\ : std_logic;
signal \N__20170\ : std_logic;
signal \N__20167\ : std_logic;
signal \N__20164\ : std_logic;
signal \N__20161\ : std_logic;
signal \N__20158\ : std_logic;
signal \N__20155\ : std_logic;
signal \N__20152\ : std_logic;
signal \N__20149\ : std_logic;
signal \N__20146\ : std_logic;
signal \N__20145\ : std_logic;
signal \N__20144\ : std_logic;
signal \N__20143\ : std_logic;
signal \N__20142\ : std_logic;
signal \N__20139\ : std_logic;
signal \N__20136\ : std_logic;
signal \N__20133\ : std_logic;
signal \N__20130\ : std_logic;
signal \N__20127\ : std_logic;
signal \N__20120\ : std_logic;
signal \N__20113\ : std_logic;
signal \N__20110\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20103\ : std_logic;
signal \N__20102\ : std_logic;
signal \N__20099\ : std_logic;
signal \N__20098\ : std_logic;
signal \N__20093\ : std_logic;
signal \N__20088\ : std_logic;
signal \N__20085\ : std_logic;
signal \N__20082\ : std_logic;
signal \N__20077\ : std_logic;
signal \N__20074\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20070\ : std_logic;
signal \N__20065\ : std_logic;
signal \N__20062\ : std_logic;
signal \N__20061\ : std_logic;
signal \N__20056\ : std_logic;
signal \N__20053\ : std_logic;
signal \N__20052\ : std_logic;
signal \N__20047\ : std_logic;
signal \N__20044\ : std_logic;
signal \N__20041\ : std_logic;
signal \N__20038\ : std_logic;
signal \N__20035\ : std_logic;
signal \N__20034\ : std_logic;
signal \N__20029\ : std_logic;
signal \N__20026\ : std_logic;
signal \N__20023\ : std_logic;
signal \N__20022\ : std_logic;
signal \N__20019\ : std_logic;
signal \N__20016\ : std_logic;
signal \N__20013\ : std_logic;
signal \N__20010\ : std_logic;
signal \N__20005\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__19999\ : std_logic;
signal \N__19996\ : std_logic;
signal \N__19993\ : std_logic;
signal \N__19992\ : std_logic;
signal \N__19989\ : std_logic;
signal \N__19986\ : std_logic;
signal \N__19981\ : std_logic;
signal \N__19980\ : std_logic;
signal \N__19977\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19971\ : std_logic;
signal \N__19966\ : std_logic;
signal \N__19963\ : std_logic;
signal \N__19960\ : std_logic;
signal \N__19957\ : std_logic;
signal \N__19954\ : std_logic;
signal \N__19953\ : std_logic;
signal \N__19950\ : std_logic;
signal \N__19947\ : std_logic;
signal \N__19942\ : std_logic;
signal \N__19939\ : std_logic;
signal \N__19936\ : std_logic;
signal \N__19933\ : std_logic;
signal \N__19930\ : std_logic;
signal \N__19929\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19925\ : std_logic;
signal \N__19922\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19912\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19906\ : std_logic;
signal \N__19903\ : std_logic;
signal \N__19900\ : std_logic;
signal \N__19897\ : std_logic;
signal \N__19894\ : std_logic;
signal \N__19893\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19891\ : std_logic;
signal \N__19890\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19888\ : std_logic;
signal \N__19885\ : std_logic;
signal \N__19872\ : std_logic;
signal \N__19867\ : std_logic;
signal \N__19864\ : std_logic;
signal \N__19863\ : std_logic;
signal \N__19860\ : std_logic;
signal \N__19859\ : std_logic;
signal \N__19854\ : std_logic;
signal \N__19851\ : std_logic;
signal \N__19848\ : std_logic;
signal \N__19843\ : std_logic;
signal \N__19840\ : std_logic;
signal \N__19837\ : std_logic;
signal \N__19834\ : std_logic;
signal \N__19831\ : std_logic;
signal \N__19828\ : std_logic;
signal \N__19825\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19819\ : std_logic;
signal \N__19816\ : std_logic;
signal \N__19813\ : std_logic;
signal \N__19812\ : std_logic;
signal \N__19809\ : std_logic;
signal \N__19806\ : std_logic;
signal \N__19801\ : std_logic;
signal \N__19798\ : std_logic;
signal \N__19795\ : std_logic;
signal \N__19792\ : std_logic;
signal \N__19789\ : std_logic;
signal \N__19786\ : std_logic;
signal \N__19783\ : std_logic;
signal \N__19780\ : std_logic;
signal \N__19777\ : std_logic;
signal \N__19774\ : std_logic;
signal \N__19771\ : std_logic;
signal \N__19768\ : std_logic;
signal \N__19765\ : std_logic;
signal \N__19762\ : std_logic;
signal \N__19759\ : std_logic;
signal \N__19758\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19756\ : std_logic;
signal \N__19755\ : std_logic;
signal \N__19752\ : std_logic;
signal \N__19751\ : std_logic;
signal \N__19750\ : std_logic;
signal \N__19749\ : std_logic;
signal \N__19746\ : std_logic;
signal \N__19745\ : std_logic;
signal \N__19744\ : std_logic;
signal \N__19741\ : std_logic;
signal \N__19738\ : std_logic;
signal \N__19737\ : std_logic;
signal \N__19736\ : std_logic;
signal \N__19735\ : std_logic;
signal \N__19734\ : std_logic;
signal \N__19733\ : std_logic;
signal \N__19732\ : std_logic;
signal \N__19729\ : std_logic;
signal \N__19726\ : std_logic;
signal \N__19723\ : std_logic;
signal \N__19720\ : std_logic;
signal \N__19717\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19692\ : std_logic;
signal \N__19689\ : std_logic;
signal \N__19674\ : std_logic;
signal \N__19669\ : std_logic;
signal \N__19666\ : std_logic;
signal \N__19663\ : std_logic;
signal \N__19660\ : std_logic;
signal \N__19657\ : std_logic;
signal \N__19654\ : std_logic;
signal \N__19653\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19651\ : std_logic;
signal \N__19648\ : std_logic;
signal \N__19645\ : std_logic;
signal \N__19642\ : std_logic;
signal \N__19641\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19637\ : std_logic;
signal \N__19626\ : std_logic;
signal \N__19623\ : std_logic;
signal \N__19618\ : std_logic;
signal \N__19617\ : std_logic;
signal \N__19616\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19600\ : std_logic;
signal \N__19597\ : std_logic;
signal \N__19596\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19589\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19579\ : std_logic;
signal \N__19578\ : std_logic;
signal \N__19577\ : std_logic;
signal \N__19576\ : std_logic;
signal \N__19575\ : std_logic;
signal \N__19574\ : std_logic;
signal \N__19569\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19563\ : std_logic;
signal \N__19562\ : std_logic;
signal \N__19561\ : std_logic;
signal \N__19560\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19558\ : std_logic;
signal \N__19553\ : std_logic;
signal \N__19552\ : std_logic;
signal \N__19551\ : std_logic;
signal \N__19550\ : std_logic;
signal \N__19547\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19530\ : std_logic;
signal \N__19527\ : std_logic;
signal \N__19520\ : std_logic;
signal \N__19507\ : std_logic;
signal \N__19506\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19500\ : std_logic;
signal \N__19497\ : std_logic;
signal \N__19492\ : std_logic;
signal \N__19491\ : std_logic;
signal \N__19488\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19484\ : std_logic;
signal \N__19479\ : std_logic;
signal \N__19474\ : std_logic;
signal \N__19473\ : std_logic;
signal \N__19472\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19468\ : std_logic;
signal \N__19467\ : std_logic;
signal \N__19466\ : std_logic;
signal \N__19461\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19459\ : std_logic;
signal \N__19458\ : std_logic;
signal \N__19457\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19447\ : std_logic;
signal \N__19444\ : std_logic;
signal \N__19437\ : std_logic;
signal \N__19434\ : std_logic;
signal \N__19433\ : std_logic;
signal \N__19432\ : std_logic;
signal \N__19431\ : std_logic;
signal \N__19430\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19417\ : std_logic;
signal \N__19410\ : std_logic;
signal \N__19407\ : std_logic;
signal \N__19396\ : std_logic;
signal \N__19393\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19389\ : std_logic;
signal \N__19386\ : std_logic;
signal \N__19383\ : std_logic;
signal \N__19378\ : std_logic;
signal \N__19377\ : std_logic;
signal \N__19376\ : std_logic;
signal \N__19373\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19359\ : std_logic;
signal \N__19356\ : std_logic;
signal \N__19355\ : std_logic;
signal \N__19348\ : std_logic;
signal \N__19345\ : std_logic;
signal \N__19344\ : std_logic;
signal \N__19339\ : std_logic;
signal \N__19336\ : std_logic;
signal \N__19335\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19327\ : std_logic;
signal \N__19326\ : std_logic;
signal \N__19323\ : std_logic;
signal \N__19318\ : std_logic;
signal \N__19315\ : std_logic;
signal \N__19314\ : std_logic;
signal \N__19309\ : std_logic;
signal \N__19306\ : std_logic;
signal \N__19303\ : std_logic;
signal \N__19302\ : std_logic;
signal \N__19299\ : std_logic;
signal \N__19294\ : std_logic;
signal \N__19291\ : std_logic;
signal \N__19290\ : std_logic;
signal \N__19287\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19280\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19270\ : std_logic;
signal \N__19269\ : std_logic;
signal \N__19268\ : std_logic;
signal \N__19265\ : std_logic;
signal \N__19262\ : std_logic;
signal \N__19259\ : std_logic;
signal \N__19256\ : std_logic;
signal \N__19251\ : std_logic;
signal \N__19246\ : std_logic;
signal \N__19243\ : std_logic;
signal \N__19240\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19238\ : std_logic;
signal \N__19233\ : std_logic;
signal \N__19230\ : std_logic;
signal \N__19225\ : std_logic;
signal \N__19224\ : std_logic;
signal \N__19219\ : std_logic;
signal \N__19216\ : std_logic;
signal \N__19213\ : std_logic;
signal \N__19210\ : std_logic;
signal \N__19209\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19205\ : std_logic;
signal \N__19202\ : std_logic;
signal \N__19199\ : std_logic;
signal \N__19192\ : std_logic;
signal \N__19191\ : std_logic;
signal \N__19190\ : std_logic;
signal \N__19187\ : std_logic;
signal \N__19182\ : std_logic;
signal \N__19177\ : std_logic;
signal \N__19176\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19172\ : std_logic;
signal \N__19167\ : std_logic;
signal \N__19162\ : std_logic;
signal \N__19161\ : std_logic;
signal \N__19158\ : std_logic;
signal \N__19157\ : std_logic;
signal \N__19154\ : std_logic;
signal \N__19149\ : std_logic;
signal \N__19144\ : std_logic;
signal \N__19141\ : std_logic;
signal \N__19140\ : std_logic;
signal \N__19135\ : std_logic;
signal \N__19134\ : std_logic;
signal \N__19131\ : std_logic;
signal \N__19128\ : std_logic;
signal \N__19123\ : std_logic;
signal \N__19122\ : std_logic;
signal \N__19119\ : std_logic;
signal \N__19116\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19109\ : std_logic;
signal \N__19106\ : std_logic;
signal \N__19099\ : std_logic;
signal \N__19096\ : std_logic;
signal \N__19093\ : std_logic;
signal \N__19090\ : std_logic;
signal \N__19087\ : std_logic;
signal \N__19084\ : std_logic;
signal \N__19081\ : std_logic;
signal \N__19078\ : std_logic;
signal \N__19075\ : std_logic;
signal \N__19072\ : std_logic;
signal \N__19069\ : std_logic;
signal \N__19066\ : std_logic;
signal \N__19063\ : std_logic;
signal \N__19060\ : std_logic;
signal \N__19057\ : std_logic;
signal \N__19054\ : std_logic;
signal \N__19051\ : std_logic;
signal \N__19048\ : std_logic;
signal \N__19045\ : std_logic;
signal \N__19042\ : std_logic;
signal \N__19039\ : std_logic;
signal \N__19036\ : std_logic;
signal \N__19033\ : std_logic;
signal \N__19030\ : std_logic;
signal \N__19027\ : std_logic;
signal \N__19024\ : std_logic;
signal \N__19021\ : std_logic;
signal \N__19018\ : std_logic;
signal \N__19015\ : std_logic;
signal \N__19012\ : std_logic;
signal \N__19009\ : std_logic;
signal \N__19006\ : std_logic;
signal \N__19003\ : std_logic;
signal \N__19000\ : std_logic;
signal \N__18997\ : std_logic;
signal \N__18994\ : std_logic;
signal \N__18991\ : std_logic;
signal \N__18988\ : std_logic;
signal \N__18985\ : std_logic;
signal \ICE_GPMO_2\ : std_logic;
signal \VCCG0\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged11WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged3WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged10WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged8WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged4WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged9WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged5WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged0WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged6WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged1WCLKN_net\ : std_logic;
signal \ICE_SYSCLK\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged7WCLKN_net\ : std_logic;
signal \INViac_raw_buf_vac_raw_buf_merged2WCLKN_net\ : std_logic;
signal \RTD_SCLK\ : std_logic;
signal \RTD.n8\ : std_logic;
signal \RTD_CS\ : std_logic;
signal \RTD.n11673\ : std_logic;
signal \n13279_cascade_\ : std_logic;
signal \RTD_SDO\ : std_logic;
signal read_buf_0 : std_logic;
signal read_buf_5 : std_logic;
signal read_buf_12 : std_logic;
signal read_buf_6 : std_logic;
signal read_buf_7 : std_logic;
signal read_buf_11 : std_logic;
signal \n11700_cascade_\ : std_logic;
signal read_buf_14 : std_logic;
signal read_buf_15 : std_logic;
signal read_buf_1 : std_logic;
signal read_buf_13 : std_logic;
signal read_buf_9 : std_logic;
signal adress_1 : std_logic;
signal adress_2 : std_logic;
signal adress_3 : std_logic;
signal adress_4 : std_logic;
signal adress_5 : std_logic;
signal read_buf_10 : std_logic;
signal n14465 : std_logic;
signal read_buf_8 : std_logic;
signal read_buf_4 : std_logic;
signal n13279 : std_logic;
signal read_buf_2 : std_logic;
signal read_buf_3 : std_logic;
signal n11700 : std_logic;
signal \RTD.n11726\ : std_logic;
signal \RTD.n15050\ : std_logic;
signal \RTD_SDI\ : std_logic;
signal \RTD.n11704\ : std_logic;
signal \RTD.n33_cascade_\ : std_logic;
signal n1_adj_1575 : std_logic;
signal \RTD.n16614\ : std_logic;
signal \RTD.n16614_cascade_\ : std_logic;
signal \RTD.n19482\ : std_logic;
signal \RTD.n19482_cascade_\ : std_logic;
signal \RTD.n7285_cascade_\ : std_logic;
signal \RTD.n21_cascade_\ : std_logic;
signal \RTD.n4\ : std_logic;
signal \RTD.n20969_cascade_\ : std_logic;
signal \RTD.n32\ : std_logic;
signal adress_6 : std_logic;
signal \RTD.adress_7\ : std_logic;
signal adress_0 : std_logic;
signal \RTD.n19855\ : std_logic;
signal \RTD.adress_7_N_1331_7_cascade_\ : std_logic;
signal \RTD_DRDY\ : std_logic;
signal \RTD.n11_cascade_\ : std_logic;
signal \RTD.n19_cascade_\ : std_logic;
signal n13151 : std_logic;
signal \RTD.n1_adj_1393\ : std_logic;
signal \RTD.adress_7_N_1331_7\ : std_logic;
signal \RTD.n16\ : std_logic;
signal \RTD.mode\ : std_logic;
signal \RTD.n10\ : std_logic;
signal \RTD.cfg_buf_2\ : std_logic;
signal \RTD.cfg_buf_4\ : std_logic;
signal \RTD.cfg_buf_7\ : std_logic;
signal \RTD.n12\ : std_logic;
signal cfg_buf_1 : std_logic;
signal \buf_readRTD_7\ : std_logic;
signal \n19_adj_1622_cascade_\ : std_logic;
signal buf_adcdata_vac_15 : std_logic;
signal buf_data_iac_3 : std_logic;
signal buf_data_iac_21 : std_logic;
signal cmd_rdadctmp_28_adj_1415 : std_logic;
signal \buf_readRTD_5\ : std_logic;
signal n14_adj_1577 : std_logic;
signal \n20573_cascade_\ : std_logic;
signal \VAC_CS\ : std_logic;
signal \VAC_SCLK\ : std_logic;
signal buf_data_iac_8 : std_logic;
signal \data_index_9_N_212_7\ : std_logic;
signal \CLK_DDS.n9\ : std_logic;
signal \RTD.bit_cnt_1\ : std_logic;
signal \RTD.bit_cnt_0\ : std_logic;
signal \RTD.bit_cnt_2\ : std_logic;
signal \RTD.n17638\ : std_logic;
signal \RTD.bit_cnt_3\ : std_logic;
signal \RTD.n17638_cascade_\ : std_logic;
signal \RTD.n1_adj_1392\ : std_logic;
signal \RTD.n21063_cascade_\ : std_logic;
signal bit_cnt_1 : std_logic;
signal bit_cnt_2 : std_logic;
signal n8_adj_1409 : std_logic;
signal \CLK_DDS.n16711\ : std_logic;
signal \RTD.n7285\ : std_logic;
signal \RTD.n11_adj_1394\ : std_logic;
signal \RTD.n21091\ : std_logic;
signal \RTD.n33\ : std_logic;
signal \RTD.n17676\ : std_logic;
signal \RTD.n7_adj_1395\ : std_logic;
signal \RTD.n11712\ : std_logic;
signal \RTD.cfg_tmp_1\ : std_logic;
signal \RTD.cfg_tmp_2\ : std_logic;
signal \RTD.cfg_tmp_3\ : std_logic;
signal \RTD.cfg_tmp_4\ : std_logic;
signal \RTD.cfg_tmp_5\ : std_logic;
signal \RTD.cfg_tmp_6\ : std_logic;
signal \RTD.cfg_tmp_7\ : std_logic;
signal \RTD.cfg_tmp_0\ : std_logic;
signal \RTD.adc_state_0\ : std_logic;
signal \n18586_cascade_\ : std_logic;
signal cfg_buf_0 : std_logic;
signal \RTD.n9\ : std_logic;
signal \RTD.n11\ : std_logic;
signal \RTD.n14\ : std_logic;
signal \RTD.n20722_cascade_\ : std_logic;
signal \RTD.n13198\ : std_logic;
signal \RTD.n13198_cascade_\ : std_logic;
signal \RTD.n14984\ : std_logic;
signal \RTD.cfg_buf_5\ : std_logic;
signal \RTD.n11_adj_1396\ : std_logic;
signal \RTD.cfg_buf_3\ : std_logic;
signal n18586 : std_logic;
signal n13162 : std_logic;
signal \RTD.cfg_buf_6\ : std_logic;
signal \buf_readRTD_11\ : std_logic;
signal \n22099_cascade_\ : std_logic;
signal \n22102_cascade_\ : std_logic;
signal buf_adcdata_vac_19 : std_logic;
signal \n19_adj_1610_cascade_\ : std_logic;
signal buf_adcdata_iac_3 : std_logic;
signal n22_adj_1611 : std_logic;
signal cmd_rdadctmp_29_adj_1414 : std_logic;
signal cmd_rdadctmp_10 : std_logic;
signal cmd_rdadctmp_26_adj_1417 : std_logic;
signal cmd_rdadctmp_27_adj_1416 : std_logic;
signal cmd_rdadctmp_9 : std_logic;
signal cmd_rdadctmp_23_adj_1420 : std_logic;
signal buf_adcdata_vac_3 : std_logic;
signal cmd_rdadctmp_8 : std_logic;
signal cmd_rdadctmp_22_adj_1421 : std_logic;
signal n19_adj_1487 : std_logic;
signal buf_adcdata_vac_8 : std_logic;
signal \buf_readRTD_0\ : std_logic;
signal \n19_adj_1479_cascade_\ : std_logic;
signal \n23_adj_1512_cascade_\ : std_logic;
signal cmd_rdadctmp_6_adj_1437 : std_logic;
signal cmd_rdadctmp_21_adj_1422 : std_logic;
signal buf_adcdata_vac_13 : std_logic;
signal cmd_rdadctmp_4_adj_1439 : std_logic;
signal cmd_rdadctmp_5_adj_1438 : std_logic;
signal buf_data_iac_14 : std_logic;
signal cmd_rdadctmp_20 : std_logic;
signal cmd_rdadctmp_21 : std_logic;
signal cmd_rdadctmp_19 : std_logic;
signal cmd_rdadctmp_18 : std_logic;
signal buf_data_iac_11 : std_logic;
signal cmd_rdadctmp_17 : std_logic;
signal buf_adcdata_iac_9 : std_logic;
signal \DDS_MCLK1\ : std_logic;
signal \DDS_CS1\ : std_logic;
signal \DDS_SCK1\ : std_logic;
signal \RTD.adc_state_3\ : std_logic;
signal \RTD.adc_state_1\ : std_logic;
signal adc_state_2_adj_1474 : std_logic;
signal \RTD.n20487\ : std_logic;
signal buf_data_iac_22 : std_logic;
signal \DDS_MOSI1\ : std_logic;
signal buf_adcdata_vac_21 : std_logic;
signal \buf_readRTD_8\ : std_logic;
signal \n22183_cascade_\ : std_logic;
signal buf_data_iac_2 : std_logic;
signal \buf_readRTD_13\ : std_logic;
signal n22153 : std_logic;
signal buf_adcdata_iac_2 : std_logic;
signal \n19_adj_1613_cascade_\ : std_logic;
signal n22_adj_1614 : std_logic;
signal \buf_readRTD_15\ : std_logic;
signal buf_adcdata_vac_2 : std_logic;
signal buf_adcdata_vac_22 : std_logic;
signal buf_adcdata_vac_14 : std_logic;
signal buf_adcdata_vac_17 : std_logic;
signal cmd_rdadctmp_30_adj_1413 : std_logic;
signal cmd_rdadctmp_31_adj_1412 : std_logic;
signal buf_adcdata_vac_16 : std_logic;
signal cmd_rdadctmp_10_adj_1433 : std_logic;
signal cmd_rdadctmp_11_adj_1432 : std_logic;
signal cmd_rdadctmp_7_adj_1436 : std_logic;
signal cmd_rdadctmp_8_adj_1435 : std_logic;
signal cmd_rdadctmp_9_adj_1434 : std_logic;
signal \VAC_MISO\ : std_logic;
signal n21973 : std_logic;
signal cmd_rdadctmp_17_adj_1426 : std_logic;
signal cmd_rdadctmp_16_adj_1427 : std_logic;
signal cmd_rdadctmp_0_adj_1443 : std_logic;
signal cmd_rdadctmp_1_adj_1442 : std_logic;
signal cmd_rdadctmp_2_adj_1441 : std_logic;
signal cmd_rdadctmp_3_adj_1440 : std_logic;
signal n20573 : std_logic;
signal \ADC_VAC.n12556_cascade_\ : std_logic;
signal \ADC_VAC.n20667\ : std_logic;
signal \ADC_VAC.n20747_cascade_\ : std_logic;
signal \ADC_VAC.n20763_cascade_\ : std_logic;
signal \ADC_VAC.n21031_cascade_\ : std_logic;
signal \ADC_VAC.n20668\ : std_logic;
signal \VAC_DRDY\ : std_logic;
signal \ADC_VAC.n17_cascade_\ : std_logic;
signal \ADC_VAC.n12\ : std_logic;
signal \ADC_VAC.bit_cnt_0\ : std_logic;
signal \bfn_7_17_0_\ : std_logic;
signal \ADC_VAC.bit_cnt_1\ : std_logic;
signal \ADC_VAC.n19357\ : std_logic;
signal \ADC_VAC.bit_cnt_2\ : std_logic;
signal \ADC_VAC.n19358\ : std_logic;
signal \ADC_VAC.bit_cnt_3\ : std_logic;
signal \ADC_VAC.n19359\ : std_logic;
signal \ADC_VAC.bit_cnt_4\ : std_logic;
signal \ADC_VAC.n19360\ : std_logic;
signal \ADC_VAC.bit_cnt_5\ : std_logic;
signal \ADC_VAC.n19361\ : std_logic;
signal \ADC_VAC.bit_cnt_6\ : std_logic;
signal \ADC_VAC.n19362\ : std_logic;
signal \ADC_VAC.n19363\ : std_logic;
signal \ADC_VAC.bit_cnt_7\ : std_logic;
signal \ADC_VAC.n12556\ : std_logic;
signal \ADC_VAC.n14829\ : std_logic;
signal \ADC_IAC.n12459_cascade_\ : std_logic;
signal \bfn_7_19_0_\ : std_logic;
signal \ADC_IAC.n19350\ : std_logic;
signal \ADC_IAC.n19351\ : std_logic;
signal \ADC_IAC.n19352\ : std_logic;
signal \ADC_IAC.n19353\ : std_logic;
signal \ADC_IAC.n19354\ : std_logic;
signal \ADC_IAC.n19355\ : std_logic;
signal \ADC_IAC.n19356\ : std_logic;
signal \ADC_IAC.n12459\ : std_logic;
signal \ADC_IAC.n14791\ : std_logic;
signal bit_cnt_0_adj_1449 : std_logic;
signal bit_cnt_3 : std_logic;
signal n21206 : std_logic;
signal buf_adcdata_vdc_3 : std_logic;
signal \CLK_DDS.n9_adj_1386\ : std_logic;
signal buf_adcdata_vdc_21 : std_logic;
signal buf_adcdata_vdc_13 : std_logic;
signal buf_adcdata_vdc_16 : std_logic;
signal buf_adcdata_vdc_2 : std_logic;
signal buf_adcdata_vdc_19 : std_logic;
signal buf_adcdata_vdc_15 : std_logic;
signal buf_adcdata_vdc_14 : std_logic;
signal buf_adcdata_vdc_22 : std_logic;
signal buf_adcdata_vdc_17 : std_logic;
signal buf_adcdata_vdc_0 : std_logic;
signal buf_adcdata_vac_0 : std_logic;
signal buf_adcdata_iac_0 : std_logic;
signal \n19_adj_1477_cascade_\ : std_logic;
signal \buf_readRTD_14\ : std_logic;
signal n22141 : std_logic;
signal \buf_readRTD_10\ : std_logic;
signal buf_adcdata_vdc_18 : std_logic;
signal buf_adcdata_vac_18 : std_logic;
signal \n21931_cascade_\ : std_logic;
signal \buf_cfgRTD_2\ : std_logic;
signal \buf_cfgRTD_3\ : std_logic;
signal \buf_cfgRTD_0\ : std_logic;
signal \n14490_cascade_\ : std_logic;
signal \buf_cfgRTD_1\ : std_logic;
signal \buf_readRTD_9\ : std_logic;
signal n22165 : std_logic;
signal buf_adcdata_iac_1 : std_logic;
signal buf_data_iac_1 : std_logic;
signal \n22_adj_1618_cascade_\ : std_logic;
signal buf_data_iac_16 : std_logic;
signal \n20781_cascade_\ : std_logic;
signal buf_adcdata_vdc_1 : std_logic;
signal buf_adcdata_vac_1 : std_logic;
signal n19_adj_1617 : std_logic;
signal \n22171_cascade_\ : std_logic;
signal n20775 : std_logic;
signal n20842 : std_logic;
signal n20843 : std_logic;
signal \n22051_cascade_\ : std_logic;
signal n20828 : std_logic;
signal n20814 : std_logic;
signal cmd_rdadctmp_24_adj_1419 : std_logic;
signal cmd_rdadctmp_25_adj_1418 : std_logic;
signal n22039 : std_logic;
signal n22042 : std_logic;
signal \buf_cfgRTD_7\ : std_logic;
signal cmd_rdadctmp_20_adj_1423 : std_logic;
signal cmd_rdadctmp_18_adj_1425 : std_logic;
signal buf_adcdata_vac_12 : std_logic;
signal buf_adcdata_vdc_10 : std_logic;
signal buf_adcdata_vac_10 : std_logic;
signal cmd_rdadctmp_19_adj_1424 : std_logic;
signal buf_data_iac_23 : std_logic;
signal \n26_adj_1511_cascade_\ : std_logic;
signal \n20834_cascade_\ : std_logic;
signal \n22057_cascade_\ : std_logic;
signal buf_data_iac_12 : std_logic;
signal n22135 : std_logic;
signal buf_adcdata_vac_23 : std_logic;
signal buf_adcdata_vdc_23 : std_logic;
signal n20831 : std_logic;
signal cmd_rdadctmp_7 : std_logic;
signal n16_adj_1507 : std_logic;
signal cmd_rdadctmp_6 : std_logic;
signal \data_index_9_N_212_8\ : std_logic;
signal cmd_rdadctmp_22 : std_logic;
signal n8_adj_1534 : std_logic;
signal buf_adcdata_iac_8 : std_logic;
signal cmd_rdadctmp_5 : std_logic;
signal buf_adcdata_iac_22 : std_logic;
signal cmd_rdadctmp_1 : std_logic;
signal n20553 : std_logic;
signal cmd_rdadctmp_29 : std_logic;
signal cmd_rdadctmp_27 : std_logic;
signal \IAC_MISO\ : std_logic;
signal cmd_rdadctmp_0 : std_logic;
signal cmd_rdadctmp_30 : std_logic;
signal cmd_rdadctmp_4 : std_logic;
signal cmd_rdadctmp_2 : std_logic;
signal cmd_rdadctmp_3 : std_logic;
signal \IAC_CS\ : std_logic;
signal n14_adj_1581 : std_logic;
signal \ADC_IAC.n20669\ : std_logic;
signal \ADC_IAC.bit_cnt_4\ : std_logic;
signal \ADC_IAC.bit_cnt_3\ : std_logic;
signal \ADC_IAC.bit_cnt_1\ : std_logic;
signal \ADC_IAC.bit_cnt_2\ : std_logic;
signal \ADC_IAC.bit_cnt_6\ : std_logic;
signal \ADC_IAC.bit_cnt_0\ : std_logic;
signal \ADC_IAC.n20753_cascade_\ : std_logic;
signal \ADC_IAC.bit_cnt_7\ : std_logic;
signal \ADC_IAC.bit_cnt_5\ : std_logic;
signal \ADC_IAC.n20765_cascade_\ : std_logic;
signal \ADC_IAC.n21007_cascade_\ : std_logic;
signal \ADC_IAC.n20670\ : std_logic;
signal \IAC_DRDY\ : std_logic;
signal \ADC_IAC.n17_cascade_\ : std_logic;
signal \ADC_IAC.n12\ : std_logic;
signal \ADC_VDC.n20345\ : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_0\ : std_logic;
signal \bfn_9_5_0_\ : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_1\ : std_logic;
signal \ADC_VDC.n19364\ : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_2\ : std_logic;
signal \ADC_VDC.n19365\ : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_3\ : std_logic;
signal \ADC_VDC.n19366\ : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_4\ : std_logic;
signal \ADC_VDC.n19367\ : std_logic;
signal cmd_rdadctmp_5_adj_1467 : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_5\ : std_logic;
signal \ADC_VDC.n19368\ : std_logic;
signal cmd_rdadctmp_6_adj_1466 : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_6\ : std_logic;
signal \ADC_VDC.n19369\ : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_7\ : std_logic;
signal \ADC_VDC.n19370\ : std_logic;
signal \ADC_VDC.n19371\ : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_8\ : std_logic;
signal \bfn_9_6_0_\ : std_logic;
signal cmd_rdadctmp_9_adj_1463 : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_9\ : std_logic;
signal \ADC_VDC.n19372\ : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_10\ : std_logic;
signal \ADC_VDC.n19373\ : std_logic;
signal cmd_rdadcbuf_11 : std_logic;
signal \ADC_VDC.n19374\ : std_logic;
signal cmd_rdadcbuf_12 : std_logic;
signal \ADC_VDC.n19375\ : std_logic;
signal cmd_rdadctmp_13_adj_1459 : std_logic;
signal cmd_rdadcbuf_13 : std_logic;
signal \ADC_VDC.n19376\ : std_logic;
signal cmd_rdadctmp_14_adj_1458 : std_logic;
signal cmd_rdadcbuf_14 : std_logic;
signal \ADC_VDC.n19377\ : std_logic;
signal \ADC_VDC.n19378\ : std_logic;
signal \ADC_VDC.n19379\ : std_logic;
signal \bfn_9_7_0_\ : std_logic;
signal \ADC_VDC.n19380\ : std_logic;
signal cmd_rdadctmp_18_adj_1454 : std_logic;
signal \ADC_VDC.n19381\ : std_logic;
signal \ADC_VDC.n19382\ : std_logic;
signal \ADC_VDC.n19383\ : std_logic;
signal cmd_rdadctmp_21_adj_1451 : std_logic;
signal cmd_rdadcbuf_21 : std_logic;
signal \ADC_VDC.n19384\ : std_logic;
signal cmd_rdadctmp_22_adj_1450 : std_logic;
signal \ADC_VDC.n19385\ : std_logic;
signal \ADC_VDC.cmd_rdadctmp_23\ : std_logic;
signal \ADC_VDC.n19386\ : std_logic;
signal \ADC_VDC.n19387\ : std_logic;
signal cmd_rdadcbuf_24 : std_logic;
signal \bfn_9_8_0_\ : std_logic;
signal cmd_rdadcbuf_25 : std_logic;
signal \ADC_VDC.n19388\ : std_logic;
signal cmd_rdadcbuf_26 : std_logic;
signal \ADC_VDC.n19389\ : std_logic;
signal cmd_rdadcbuf_27 : std_logic;
signal \ADC_VDC.n19390\ : std_logic;
signal cmd_rdadcbuf_28 : std_logic;
signal \ADC_VDC.n19391\ : std_logic;
signal cmd_rdadcbuf_29 : std_logic;
signal \ADC_VDC.n19392\ : std_logic;
signal cmd_rdadcbuf_30 : std_logic;
signal \ADC_VDC.n19393\ : std_logic;
signal cmd_rdadcbuf_31 : std_logic;
signal \ADC_VDC.n19394\ : std_logic;
signal \ADC_VDC.n19395\ : std_logic;
signal cmd_rdadcbuf_32 : std_logic;
signal \bfn_9_9_0_\ : std_logic;
signal cmd_rdadcbuf_33 : std_logic;
signal \ADC_VDC.n19396\ : std_logic;
signal \ADC_VDC.n19397\ : std_logic;
signal n20772 : std_logic;
signal n21943 : std_logic;
signal \n21946_cascade_\ : std_logic;
signal n22060 : std_logic;
signal n22054 : std_logic;
signal \n22015_cascade_\ : std_logic;
signal buf_data_iac_17 : std_logic;
signal \n20818_cascade_\ : std_logic;
signal n20871 : std_logic;
signal \n20820_cascade_\ : std_logic;
signal n21967 : std_logic;
signal n21970 : std_logic;
signal \n22003_cascade_\ : std_logic;
signal \n20624_cascade_\ : std_logic;
signal \SIG_DDS.n10_cascade_\ : std_logic;
signal \buf_readRTD_12\ : std_logic;
signal n22006 : std_logic;
signal \n22027_cascade_\ : std_logic;
signal n22030 : std_logic;
signal buf_adcdata_vac_20 : std_logic;
signal buf_adcdata_vdc_20 : std_logic;
signal n22207 : std_logic;
signal n20801 : std_logic;
signal buf_adcdata_iac_10 : std_logic;
signal \SIG_DDS.bit_cnt_1\ : std_logic;
signal \SIG_DDS.bit_cnt_2\ : std_logic;
signal buf_adcdata_vac_11 : std_logic;
signal cmd_rdadctmp_23 : std_logic;
signal n8 : std_logic;
signal n22117 : std_logic;
signal buf_adcdata_iac_13 : std_logic;
signal \SIG_DDS.bit_cnt_3\ : std_logic;
signal \SIG_DDS.n21292\ : std_logic;
signal \VAC_OSR0\ : std_logic;
signal buf_adcdata_iac_19 : std_logic;
signal n11417 : std_logic;
signal buf_adcdata_iac_17 : std_logic;
signal \n22201_cascade_\ : std_logic;
signal n20805 : std_logic;
signal cmd_rdadctmp_24 : std_logic;
signal cmd_rdadctmp_31 : std_logic;
signal buf_adcdata_iac_23 : std_logic;
signal \AC_ADC_SYNC\ : std_logic;
signal \VAC_FLT1\ : std_logic;
signal \IAC_SCLK\ : std_logic;
signal \ADC_VDC.n18394_cascade_\ : std_logic;
signal \EIS_SYNCCLK\ : std_logic;
signal \IAC_CLK\ : std_logic;
signal \ADC_VDC.n31_cascade_\ : std_logic;
signal \ADC_VDC.n21925_cascade_\ : std_logic;
signal \ADC_VDC.n18397\ : std_logic;
signal \ADC_VDC.n21928_cascade_\ : std_logic;
signal \ADC_VDC.n20514\ : std_logic;
signal \ADC_VDC.n6_cascade_\ : std_logic;
signal \ADC_VDC.n10519\ : std_logic;
signal \n12853_cascade_\ : std_logic;
signal cmd_rdadctmp_0_adj_1472 : std_logic;
signal cmd_rdadctmp_3_adj_1469 : std_logic;
signal cmd_rdadctmp_4_adj_1468 : std_logic;
signal \ADC_VDC.n12885\ : std_logic;
signal cmd_rdadctmp_7_adj_1465 : std_logic;
signal cmd_rdadctmp_8_adj_1464 : std_logic;
signal cmd_rdadctmp_17_adj_1455 : std_logic;
signal cmd_rdadctmp_15_adj_1457 : std_logic;
signal cmd_rdadctmp_16_adj_1456 : std_logic;
signal cmd_rdadctmp_1_adj_1471 : std_logic;
signal cmd_rdadctmp_2_adj_1470 : std_logic;
signal cmd_rdadctmp_12_adj_1460 : std_logic;
signal cmd_rdadctmp_10_adj_1462 : std_logic;
signal cmd_rdadctmp_11_adj_1461 : std_logic;
signal \ADC_VDC.n21673_cascade_\ : std_logic;
signal \VDC_SCLK\ : std_logic;
signal cmd_rdadctmp_19_adj_1453 : std_logic;
signal n12853 : std_logic;
signal cmd_rdadctmp_20_adj_1452 : std_logic;
signal cmd_rdadcbuf_23 : std_logic;
signal buf_adcdata_vdc_12 : std_logic;
signal cmd_rdadcbuf_22 : std_logic;
signal buf_adcdata_vdc_11 : std_logic;
signal cmd_rdadcbuf_15 : std_logic;
signal cmd_rdadcbuf_20 : std_logic;
signal cmd_rdadcbuf_19 : std_logic;
signal buf_adcdata_vdc_8 : std_logic;
signal cmd_rdadcbuf_18 : std_logic;
signal cmd_rdadcbuf_17 : std_logic;
signal cmd_rdadcbuf_16 : std_logic;
signal \ADC_VDC.n18394\ : std_logic;
signal \ADC_VDC.cmd_rdadcbuf_35_N_1130_34\ : std_logic;
signal \ADC_VDC.n21106_cascade_\ : std_logic;
signal cmd_rdadcbuf_34 : std_logic;
signal \ADC_VDC.n13020\ : std_logic;
signal \ADC_VDC.n21\ : std_logic;
signal \ADC_VDC.n19\ : std_logic;
signal buf_data_vac_16 : std_logic;
signal buf_data_vac_23 : std_logic;
signal buf_data_vac_22 : std_logic;
signal buf_data_vac_21 : std_logic;
signal buf_data_vac_20 : std_logic;
signal buf_data_vac_19 : std_logic;
signal buf_data_vac_18 : std_logic;
signal buf_data_vac_17 : std_logic;
signal \n21143_cascade_\ : std_logic;
signal \n12_cascade_\ : std_logic;
signal n12116 : std_logic;
signal \n12116_cascade_\ : std_logic;
signal n14756 : std_logic;
signal \n25_adj_1592_cascade_\ : std_logic;
signal \n11944_cascade_\ : std_logic;
signal \n11941_cascade_\ : std_logic;
signal \n21919_cascade_\ : std_logic;
signal buf_data_iac_18 : std_logic;
signal \n20794_cascade_\ : std_logic;
signal n21922 : std_logic;
signal \n20796_cascade_\ : std_logic;
signal n21934 : std_logic;
signal \n22213_cascade_\ : std_logic;
signal \n22216_cascade_\ : std_logic;
signal n20937 : std_logic;
signal n20936 : std_logic;
signal \n21907_cascade_\ : std_logic;
signal buf_adcdata_iac_21 : std_logic;
signal \n22033_cascade_\ : std_logic;
signal \n22036_cascade_\ : std_logic;
signal n22156 : std_logic;
signal n21910 : std_logic;
signal \n20823_cascade_\ : std_logic;
signal \n30_adj_1514_cascade_\ : std_logic;
signal n11941 : std_logic;
signal n14735 : std_logic;
signal \CLK_DDS.tmp_buf_10\ : std_logic;
signal \CLK_DDS.tmp_buf_11\ : std_logic;
signal \CLK_DDS.tmp_buf_12\ : std_logic;
signal \CLK_DDS.tmp_buf_13\ : std_logic;
signal \CLK_DDS.tmp_buf_14\ : std_logic;
signal \CLK_DDS.tmp_buf_9\ : std_logic;
signal \CLK_DDS.tmp_buf_8\ : std_logic;
signal buf_dds1_14 : std_logic;
signal buf_dds1_12 : std_logic;
signal buf_dds1_9 : std_logic;
signal tmp_buf_15_adj_1448 : std_logic;
signal \CLK_DDS.tmp_buf_0\ : std_logic;
signal \CLK_DDS.tmp_buf_1\ : std_logic;
signal \CLK_DDS.tmp_buf_2\ : std_logic;
signal \CLK_DDS.tmp_buf_3\ : std_logic;
signal \CLK_DDS.tmp_buf_4\ : std_logic;
signal \CLK_DDS.tmp_buf_5\ : std_logic;
signal \CLK_DDS.tmp_buf_6\ : std_logic;
signal \CLK_DDS.tmp_buf_7\ : std_logic;
signal buf_dds1_15 : std_logic;
signal n22045 : std_logic;
signal n22048 : std_logic;
signal \VAC_FLT0\ : std_logic;
signal n16_adj_1480 : std_logic;
signal buf_dds1_0 : std_logic;
signal buf_adcdata_iac_18 : std_logic;
signal cmd_rdadctmp_25 : std_logic;
signal cmd_rdadctmp_26 : std_logic;
signal n23_adj_1513 : std_logic;
signal cmd_rdadctmp_28 : std_logic;
signal buf_adcdata_iac_20 : std_logic;
signal \IAC_FLT1\ : std_logic;
signal \IAC_OSR1\ : std_logic;
signal \IAC_FLT0\ : std_logic;
signal buf_adcdata_iac_16 : std_logic;
signal buf_dds1_8 : std_logic;
signal \n22189_cascade_\ : std_logic;
signal n20769 : std_logic;
signal n16_adj_1489 : std_logic;
signal \IAC_OSR0\ : std_logic;
signal \bfn_11_3_0_\ : std_logic;
signal \ADC_VDC.genclk.n19410\ : std_logic;
signal \ADC_VDC.genclk.n19411\ : std_logic;
signal \ADC_VDC.genclk.n19412\ : std_logic;
signal \ADC_VDC.genclk.n19413\ : std_logic;
signal \ADC_VDC.genclk.n19414\ : std_logic;
signal \ADC_VDC.genclk.n19415\ : std_logic;
signal \ADC_VDC.genclk.n19416\ : std_logic;
signal \ADC_VDC.genclk.n19417\ : std_logic;
signal \INVADC_VDC.genclk.t0off_i0C_net\ : std_logic;
signal \bfn_11_4_0_\ : std_logic;
signal \ADC_VDC.genclk.n19418\ : std_logic;
signal \ADC_VDC.genclk.n19419\ : std_logic;
signal \ADC_VDC.genclk.n19420\ : std_logic;
signal \ADC_VDC.genclk.n19421\ : std_logic;
signal \ADC_VDC.genclk.n19422\ : std_logic;
signal \ADC_VDC.genclk.n19423\ : std_logic;
signal \ADC_VDC.genclk.n19424\ : std_logic;
signal \INVADC_VDC.genclk.t0off_i8C_net\ : std_logic;
signal n13073 : std_logic;
signal \ADC_VDC.n20618_cascade_\ : std_logic;
signal \ADC_VDC.n47\ : std_logic;
signal \ADC_VDC.n20702\ : std_logic;
signal \ADC_VDC.n20\ : std_logic;
signal dds_state_1_adj_1446 : std_logic;
signal dds_state_2_adj_1445 : std_logic;
signal trig_dds1 : std_logic;
signal dds_state_0_adj_1447 : std_logic;
signal \CLK_DDS.n12722\ : std_logic;
signal \ADC_VDC.avg_cnt_0\ : std_logic;
signal \bfn_11_7_0_\ : std_logic;
signal \ADC_VDC.avg_cnt_1\ : std_logic;
signal \ADC_VDC.n19399\ : std_logic;
signal \ADC_VDC.avg_cnt_2\ : std_logic;
signal \ADC_VDC.n19400\ : std_logic;
signal \ADC_VDC.avg_cnt_3\ : std_logic;
signal \ADC_VDC.n19401\ : std_logic;
signal \ADC_VDC.avg_cnt_4\ : std_logic;
signal \ADC_VDC.n19402\ : std_logic;
signal \ADC_VDC.avg_cnt_5\ : std_logic;
signal \ADC_VDC.n19403\ : std_logic;
signal \ADC_VDC.avg_cnt_6\ : std_logic;
signal \ADC_VDC.n19404\ : std_logic;
signal \ADC_VDC.avg_cnt_7\ : std_logic;
signal \ADC_VDC.n19405\ : std_logic;
signal \ADC_VDC.n19406\ : std_logic;
signal \ADC_VDC.avg_cnt_8\ : std_logic;
signal \bfn_11_8_0_\ : std_logic;
signal \ADC_VDC.avg_cnt_9\ : std_logic;
signal \ADC_VDC.n19407\ : std_logic;
signal \ADC_VDC.avg_cnt_10\ : std_logic;
signal \ADC_VDC.n19408\ : std_logic;
signal \ADC_VDC.n19409\ : std_logic;
signal \ADC_VDC.avg_cnt_11\ : std_logic;
signal \ADC_VDC.n13060\ : std_logic;
signal \ADC_VDC.n14900\ : std_logic;
signal \n23_adj_1510_cascade_\ : std_logic;
signal n20833 : std_logic;
signal buf_data_iac_20 : std_logic;
signal n20810 : std_logic;
signal \THERMOSTAT\ : std_logic;
signal buf_control_7 : std_logic;
signal \n21050_cascade_\ : std_logic;
signal n11905 : std_logic;
signal \buf_cfgRTD_6\ : std_logic;
signal \n11882_cascade_\ : std_logic;
signal comm_cmd_4 : std_logic;
signal comm_cmd_6 : std_logic;
signal comm_cmd_5 : std_logic;
signal \n8_adj_1522_cascade_\ : std_logic;
signal \n12214_cascade_\ : std_logic;
signal buf_dds1_13 : std_logic;
signal buf_dds1_11 : std_logic;
signal n22075 : std_logic;
signal n22078 : std_logic;
signal buf_dds1_5 : std_logic;
signal n7 : std_logic;
signal n12214 : std_logic;
signal \n16539_cascade_\ : std_logic;
signal \n17_adj_1601_cascade_\ : std_logic;
signal n16547 : std_logic;
signal \n16547_cascade_\ : std_logic;
signal \n13_cascade_\ : std_logic;
signal \INVeis_state_i0C_net\ : std_logic;
signal n19_adj_1482 : std_logic;
signal \buf_readRTD_6\ : std_logic;
signal \n21937_cascade_\ : std_logic;
signal buf_adcdata_iac_14 : std_logic;
signal \n21940_cascade_\ : std_logic;
signal \n30_adj_1490_cascade_\ : std_logic;
signal n26_adj_1495 : std_logic;
signal n21109 : std_logic;
signal \n22111_cascade_\ : std_logic;
signal n22114 : std_logic;
signal n8_adj_1536 : std_logic;
signal \AMPV_POW\ : std_logic;
signal \DTRIG_N_910\ : std_logic;
signal adc_state_1 : std_logic;
signal n10503 : std_logic;
signal \DTRIG_N_910_adj_1444\ : std_logic;
signal adc_state_1_adj_1410 : std_logic;
signal \VAC_OSR1\ : std_logic;
signal \n4_adj_1473_cascade_\ : std_logic;
signal \acadc_skipCount_13\ : std_logic;
signal buf_dds1_10 : std_logic;
signal n22147 : std_logic;
signal n22150 : std_logic;
signal \n20690_cascade_\ : std_logic;
signal acadc_trig : std_logic;
signal n20529 : std_logic;
signal eis_end : std_logic;
signal \INVacadc_trig_300C_net\ : std_logic;
signal eis_start : std_logic;
signal n17357 : std_logic;
signal \n11_adj_1620_cascade_\ : std_logic;
signal n11730 : std_logic;
signal \ADC_VDC.genclk.t0off_6\ : std_logic;
signal \ADC_VDC.genclk.t0off_1\ : std_logic;
signal \ADC_VDC.genclk.t0off_4\ : std_logic;
signal \ADC_VDC.genclk.t0off_0\ : std_logic;
signal \ADC_VDC.genclk.n21169_cascade_\ : std_logic;
signal \ADC_VDC.genclk.t0off_12\ : std_logic;
signal \ADC_VDC.genclk.t0off_2\ : std_logic;
signal \ADC_VDC.genclk.t0off_7\ : std_logic;
signal \ADC_VDC.genclk.t0off_10\ : std_logic;
signal \ADC_VDC.genclk.n27\ : std_logic;
signal \ADC_VDC.genclk.t0off_13\ : std_logic;
signal \ADC_VDC.genclk.t0off_8\ : std_logic;
signal \ADC_VDC.genclk.t0off_5\ : std_logic;
signal \ADC_VDC.genclk.t0off_3\ : std_logic;
signal \ADC_VDC.genclk.n26\ : std_logic;
signal \ADC_VDC.genclk.t0off_14\ : std_logic;
signal \ADC_VDC.genclk.t0off_9\ : std_logic;
signal \ADC_VDC.genclk.t0off_15\ : std_logic;
signal \ADC_VDC.genclk.t0off_11\ : std_logic;
signal \ADC_VDC.genclk.n28\ : std_logic;
signal \ADC_VDC.genclk.n11721\ : std_logic;
signal \ADC_VDC.n10112_cascade_\ : std_logic;
signal \ADC_VDC.n12793\ : std_logic;
signal \ADC_VDC.n17\ : std_logic;
signal \ADC_VDC.n4\ : std_logic;
signal \ADC_VDC.n12\ : std_logic;
signal \ADC_VDC.n72\ : std_logic;
signal \ADC_VDC.n20710\ : std_logic;
signal \ADC_VDC.n20490_cascade_\ : std_logic;
signal \ADC_VDC.n11251_cascade_\ : std_logic;
signal \ADC_VDC.n20523_cascade_\ : std_logic;
signal \ADC_VDC.n21178\ : std_logic;
signal \ADC_VDC.n20490\ : std_logic;
signal \ADC_VDC.n21025\ : std_logic;
signal \ADC_VDC.n7_adj_1403\ : std_logic;
signal \ADC_VDC.n20712\ : std_logic;
signal \ADC_VDC.n11662\ : std_logic;
signal \ADC_VDC.n21028\ : std_logic;
signal comm_buf_0_7 : std_logic;
signal \ADC_VDC.n10\ : std_logic;
signal \ADC_VDC.n15\ : std_logic;
signal \ADC_VDC.n19_adj_1405\ : std_logic;
signal wdtick_cnt_0 : std_logic;
signal wdtick_cnt_1 : std_logic;
signal wdtick_cnt_2 : std_logic;
signal n14490 : std_logic;
signal n11882 : std_logic;
signal buf_data_iac_0 : std_logic;
signal n22_adj_1476 : std_logic;
signal buf_data_vac_8 : std_logic;
signal buf_data_vac_15 : std_logic;
signal buf_data_vac_14 : std_logic;
signal buf_data_vac_13 : std_logic;
signal buf_data_vac_12 : std_logic;
signal buf_data_vac_11 : std_logic;
signal buf_data_vac_10 : std_logic;
signal buf_data_vac_9 : std_logic;
signal n14_adj_1516 : std_logic;
signal \bfn_12_12_0_\ : std_logic;
signal n19335 : std_logic;
signal n19336 : std_logic;
signal n19337 : std_logic;
signal n19338 : std_logic;
signal n19339 : std_logic;
signal data_idxvec_6 : std_logic;
signal n19340 : std_logic;
signal n19341 : std_logic;
signal n19342 : std_logic;
signal \bfn_12_13_0_\ : std_logic;
signal data_idxvec_9 : std_logic;
signal n19343 : std_logic;
signal data_idxvec_10 : std_logic;
signal n19344 : std_logic;
signal n19345 : std_logic;
signal data_idxvec_12 : std_logic;
signal n19346 : std_logic;
signal data_idxvec_13 : std_logic;
signal n19347 : std_logic;
signal data_idxvec_14 : std_logic;
signal n19348 : std_logic;
signal n19349 : std_logic;
signal data_idxvec_15 : std_logic;
signal data_idxvec_5 : std_logic;
signal \n26_adj_1486_cascade_\ : std_logic;
signal \n22177_cascade_\ : std_logic;
signal n22120 : std_logic;
signal \n22180_cascade_\ : std_logic;
signal \n30_adj_1485_cascade_\ : std_logic;
signal buf_data_iac_13 : std_logic;
signal n21036 : std_logic;
signal \data_index_9_N_212_0\ : std_logic;
signal \acadc_skipCount_8\ : std_logic;
signal \n20_cascade_\ : std_logic;
signal n14_adj_1498 : std_logic;
signal n18_adj_1587 : std_logic;
signal \n26_adj_1604_cascade_\ : std_logic;
signal n31 : std_logic;
signal \data_index_9_N_212_3\ : std_logic;
signal \acadc_skipCount_5\ : std_logic;
signal n16_adj_1504 : std_logic;
signal buf_dds1_1 : std_logic;
signal \acadc_skipCount_6\ : std_logic;
signal n17 : std_logic;
signal acadc_dtrig_v : std_logic;
signal acadc_dtrig_i : std_logic;
signal \iac_raw_buf_N_728_cascade_\ : std_logic;
signal n21997 : std_logic;
signal buf_dds1_3 : std_logic;
signal n20624 : std_logic;
signal \n12353_cascade_\ : std_logic;
signal n35 : std_logic;
signal \iac_raw_buf_N_726\ : std_logic;
signal \eis_end_N_716\ : std_logic;
signal acadc_rst : std_logic;
signal buf_data_iac_15 : std_logic;
signal buf_dds1_2 : std_logic;
signal buf_adcdata_iac_15 : std_logic;
signal n21961 : std_logic;
signal \n16_adj_1621_cascade_\ : std_logic;
signal buf_dds0_10 : std_logic;
signal \SIG_DDS.tmp_buf_10\ : std_logic;
signal buf_dds0_9 : std_logic;
signal \SIG_DDS.tmp_buf_9\ : std_logic;
signal buf_dds0_13 : std_logic;
signal \SIG_DDS.tmp_buf_13\ : std_logic;
signal buf_dds0_14 : std_logic;
signal buf_dds0_1 : std_logic;
signal \SIG_DDS.tmp_buf_7\ : std_logic;
signal \SIG_DDS.tmp_buf_8\ : std_logic;
signal \comm_spi.n22629\ : std_logic;
signal \comm_spi.n22629_cascade_\ : std_logic;
signal \INVADC_VDC.genclk.t_clk_24C_net\ : std_logic;
signal \comm_spi.n22632_cascade_\ : std_logic;
signal \comm_spi.imosi_cascade_\ : std_logic;
signal \comm_spi.imosi\ : std_logic;
signal \comm_spi.n14599\ : std_logic;
signal \comm_spi.DOUT_7__N_738\ : std_logic;
signal \ADC_VDC.genclk.n21167\ : std_logic;
signal \ADC_VDC.n11_cascade_\ : std_logic;
signal \ADC_VDC.n17359\ : std_logic;
signal \ADC_VDC.bit_cnt_0\ : std_logic;
signal \bfn_13_6_0_\ : std_logic;
signal \ADC_VDC.bit_cnt_1\ : std_logic;
signal \ADC_VDC.n19469\ : std_logic;
signal \ADC_VDC.n19470\ : std_logic;
signal \ADC_VDC.n19471\ : std_logic;
signal \ADC_VDC.bit_cnt_4\ : std_logic;
signal \ADC_VDC.n19472\ : std_logic;
signal \ADC_VDC.bit_cnt_5\ : std_logic;
signal \ADC_VDC.n19473\ : std_logic;
signal \ADC_VDC.bit_cnt_6\ : std_logic;
signal \ADC_VDC.n19474\ : std_logic;
signal \ADC_VDC.n19475\ : std_logic;
signal \ADC_VDC.bit_cnt_7\ : std_logic;
signal \VDC_CLK\ : std_logic;
signal \ADC_VDC.n18381\ : std_logic;
signal \INVcomm_spi.imiso_83_12193_12194_setC_net\ : std_logic;
signal buf_data_iac_6 : std_logic;
signal \ADC_VDC.bit_cnt_3\ : std_logic;
signal \ADC_VDC.bit_cnt_2\ : std_logic;
signal \ADC_VDC.n6_adj_1404\ : std_logic;
signal \comm_spi.data_tx_7__N_762\ : std_logic;
signal n11727 : std_logic;
signal \INVcomm_spi.bit_cnt_3767__i1C_net\ : std_logic;
signal \comm_spi.bit_cnt_1\ : std_logic;
signal \comm_spi.bit_cnt_0\ : std_logic;
signal \comm_spi.bit_cnt_2\ : std_logic;
signal comm_buf_3_1 : std_logic;
signal \n21991_cascade_\ : std_logic;
signal n14763 : std_logic;
signal comm_buf_3_3 : std_logic;
signal \n21979_cascade_\ : std_logic;
signal comm_buf_4_3 : std_logic;
signal comm_buf_6_3 : std_logic;
signal \n4_adj_1567_cascade_\ : std_logic;
signal \n20783_cascade_\ : std_logic;
signal n21982 : std_logic;
signal comm_buf_3_5 : std_logic;
signal \n17331_cascade_\ : std_logic;
signal \n20903_cascade_\ : std_logic;
signal \n1_adj_1561_cascade_\ : std_logic;
signal comm_buf_6_6 : std_logic;
signal comm_buf_3_6 : std_logic;
signal n2_adj_1562 : std_logic;
signal comm_buf_4_6 : std_logic;
signal n21051 : std_logic;
signal \n4_adj_1563_cascade_\ : std_logic;
signal n22093 : std_logic;
signal data_idxvec_2 : std_logic;
signal \n26_adj_1506_cascade_\ : std_logic;
signal buf_data_iac_10 : std_logic;
signal \n20816_cascade_\ : std_logic;
signal n20845 : std_logic;
signal \n22087_cascade_\ : std_logic;
signal \n22090_cascade_\ : std_logic;
signal n19_adj_1505 : std_logic;
signal \buf_readRTD_2\ : std_logic;
signal n20846 : std_logic;
signal n20815 : std_logic;
signal n19 : std_logic;
signal \buf_readRTD_4\ : std_logic;
signal buf_adcdata_iac_12 : std_logic;
signal \n22081_cascade_\ : std_logic;
signal data_idxvec_4 : std_logic;
signal n21261 : std_logic;
signal \n26_adj_1484_cascade_\ : std_logic;
signal \n22159_cascade_\ : std_logic;
signal n22084 : std_logic;
signal \n22162_cascade_\ : std_logic;
signal \n30_adj_1493_cascade_\ : std_logic;
signal data_idxvec_3 : std_logic;
signal n21285 : std_logic;
signal \n26_adj_1502_cascade_\ : std_logic;
signal \n22195_cascade_\ : std_logic;
signal \acadc_skipCount_3\ : std_logic;
signal \n22198_cascade_\ : std_logic;
signal \n30_adj_1503_cascade_\ : std_logic;
signal n19_adj_1501 : std_logic;
signal \buf_readRTD_3\ : std_logic;
signal buf_adcdata_iac_11 : std_logic;
signal \n22009_cascade_\ : std_logic;
signal n16_adj_1500 : std_logic;
signal n22012 : std_logic;
signal acadc_skipcnt_0 : std_logic;
signal \bfn_13_16_0_\ : std_logic;
signal \INVacadc_skipcnt_i0_i0C_net\ : std_logic;
signal n20757 : std_logic;
signal n19311 : std_logic;
signal \n19311_THRU_CRY_0_THRU_CO\ : std_logic;
signal \n19311_THRU_CRY_1_THRU_CO\ : std_logic;
signal \n19311_THRU_CRY_2_THRU_CO\ : std_logic;
signal \n19311_THRU_CRY_3_THRU_CO\ : std_logic;
signal \n19311_THRU_CRY_4_THRU_CO\ : std_logic;
signal \GNDG0\ : std_logic;
signal \n19311_THRU_CRY_5_THRU_CO\ : std_logic;
signal \n19311_THRU_CRY_6_THRU_CO\ : std_logic;
signal acadc_skipcnt_1 : std_logic;
signal \bfn_13_17_0_\ : std_logic;
signal n19312 : std_logic;
signal acadc_skipcnt_3 : std_logic;
signal n19313 : std_logic;
signal acadc_skipcnt_4 : std_logic;
signal n19314 : std_logic;
signal acadc_skipcnt_5 : std_logic;
signal n19315 : std_logic;
signal acadc_skipcnt_6 : std_logic;
signal n19316 : std_logic;
signal n19317 : std_logic;
signal acadc_skipcnt_8 : std_logic;
signal n19318 : std_logic;
signal n19319 : std_logic;
signal \INVacadc_skipcnt_i0_i1C_net\ : std_logic;
signal \bfn_13_18_0_\ : std_logic;
signal n19320 : std_logic;
signal n19321 : std_logic;
signal n19322 : std_logic;
signal acadc_skipcnt_13 : std_logic;
signal n19323 : std_logic;
signal n19324 : std_logic;
signal n19325 : std_logic;
signal \INVacadc_skipcnt_i0_i9C_net\ : std_logic;
signal n11538 : std_logic;
signal n14639 : std_logic;
signal \SIG_DDS.tmp_buf_11\ : std_logic;
signal buf_dds0_12 : std_logic;
signal \SIG_DDS.tmp_buf_12\ : std_logic;
signal \SIG_DDS.tmp_buf_1\ : std_logic;
signal \comm_spi.n22632\ : std_logic;
signal \comm_spi.n14600\ : std_logic;
signal \comm_spi.DOUT_7__N_739\ : std_logic;
signal \ADC_VDC.genclk.n21172_cascade_\ : std_logic;
signal \ADC_VDC.genclk.n21166\ : std_logic;
signal \ADC_VDC.genclk.n28_adj_1400\ : std_logic;
signal \ADC_VDC.genclk.n26_adj_1401\ : std_logic;
signal \ADC_VDC.genclk.n27_adj_1402\ : std_logic;
signal \comm_spi.n14586\ : std_logic;
signal \ADC_VDC.genclk.div_state_0\ : std_logic;
signal \ADC_VDC.genclk.div_state_1\ : std_logic;
signal \INVADC_VDC.genclk.div_state_i1C_net\ : std_logic;
signal \ADC_VDC.genclk.n6\ : std_logic;
signal \VDC_SDO\ : std_logic;
signal \ADC_VDC.adc_state_0\ : std_logic;
signal \ADC_VDC.n62\ : std_logic;
signal adc_state_2 : std_logic;
signal adc_state_3 : std_logic;
signal \ADC_VDC.n62_cascade_\ : std_logic;
signal \ADC_VDC.adc_state_1\ : std_logic;
signal \ADC_VDC.n11736\ : std_logic;
signal comm_buf_3_7 : std_logic;
signal n1 : std_logic;
signal \n2_adj_1559_cascade_\ : std_logic;
signal comm_buf_4_7 : std_logic;
signal comm_buf_6_7 : std_logic;
signal n4_adj_1560 : std_logic;
signal \n21276_cascade_\ : std_logic;
signal n22105 : std_logic;
signal comm_buf_3_2 : std_logic;
signal \n21985_cascade_\ : std_logic;
signal \n21988_cascade_\ : std_logic;
signal comm_buf_3_0 : std_logic;
signal \n17304_cascade_\ : std_logic;
signal \n20906_cascade_\ : std_logic;
signal comm_buf_4_2 : std_logic;
signal comm_buf_6_2 : std_logic;
signal \n4_adj_1568_cascade_\ : std_logic;
signal n20786 : std_logic;
signal n30_adj_1475 : std_logic;
signal comm_buf_2_7 : std_logic;
signal n30_adj_1595 : std_logic;
signal comm_buf_2_6 : std_logic;
signal n30_adj_1612 : std_logic;
signal comm_buf_2_3 : std_logic;
signal n30_adj_1615 : std_logic;
signal comm_buf_2_2 : std_logic;
signal n30_adj_1619 : std_logic;
signal comm_buf_2_1 : std_logic;
signal buf_data_vac_0 : std_logic;
signal comm_buf_5_0 : std_logic;
signal buf_data_vac_7 : std_logic;
signal comm_buf_5_7 : std_logic;
signal comm_rx_buf_6 : std_logic;
signal buf_data_vac_6 : std_logic;
signal comm_buf_5_6 : std_logic;
signal buf_data_vac_5 : std_logic;
signal comm_buf_5_5 : std_logic;
signal comm_rx_buf_4 : std_logic;
signal buf_data_vac_4 : std_logic;
signal comm_rx_buf_3 : std_logic;
signal buf_data_vac_3 : std_logic;
signal comm_buf_5_3 : std_logic;
signal comm_rx_buf_2 : std_logic;
signal buf_data_vac_2 : std_logic;
signal comm_buf_5_2 : std_logic;
signal buf_data_vac_1 : std_logic;
signal \buf_readRTD_1\ : std_logic;
signal buf_adcdata_vdc_9 : std_logic;
signal buf_adcdata_vac_9 : std_logic;
signal n19_adj_1508 : std_logic;
signal n20836 : std_logic;
signal \n22069_cascade_\ : std_logic;
signal n20837 : std_logic;
signal data_idxvec_1 : std_logic;
signal \n26_adj_1509_cascade_\ : std_logic;
signal buf_data_iac_9 : std_logic;
signal n20825 : std_logic;
signal comm_rx_buf_1 : std_logic;
signal n22072 : std_logic;
signal data_idxvec_0 : std_logic;
signal n21001 : std_logic;
signal \n26_cascade_\ : std_logic;
signal \acadc_skipCount_0\ : std_logic;
signal \n22021_cascade_\ : std_logic;
signal n22024 : std_logic;
signal n21976 : std_logic;
signal \n30_adj_1478_cascade_\ : std_logic;
signal comm_rx_buf_0 : std_logic;
signal cmd_rdadctmp_13_adj_1430 : std_logic;
signal buf_dds1_4 : std_logic;
signal n16 : std_logic;
signal buf_dds1_6 : std_logic;
signal n16_adj_1488 : std_logic;
signal n20824 : std_logic;
signal \data_index_9_N_212_2\ : std_logic;
signal acadc_skipcnt_14 : std_logic;
signal acadc_skipcnt_11 : std_logic;
signal comm_buf_1_3 : std_logic;
signal n8_adj_1543 : std_logic;
signal acadc_skipcnt_2 : std_logic;
signal acadc_skipcnt_7 : std_logic;
signal \acadc_skipCount_2\ : std_logic;
signal n23_adj_1586 : std_logic;
signal \n22_cascade_\ : std_logic;
signal n30_adj_1571 : std_logic;
signal data_idxvec_7 : std_logic;
signal \acadc_skipCount_14\ : std_logic;
signal n8_adj_1545 : std_logic;
signal acadc_skipcnt_9 : std_logic;
signal acadc_skipcnt_15 : std_logic;
signal \acadc_skipCount_15\ : std_logic;
signal n24 : std_logic;
signal \acadc_skipCount_1\ : std_logic;
signal n9_adj_1407 : std_logic;
signal n20949 : std_logic;
signal n26_adj_1623 : std_logic;
signal \n21949_cascade_\ : std_logic;
signal \acadc_skipCount_7\ : std_logic;
signal n21964 : std_logic;
signal \n21952_cascade_\ : std_logic;
signal \acadc_skipCount_4\ : std_logic;
signal \acadc_skipCount_9\ : std_logic;
signal comm_rx_buf_7 : std_logic;
signal n30_adj_1624 : std_logic;
signal n14742 : std_logic;
signal buf_dds0_3 : std_logic;
signal \SIG_DDS.tmp_buf_2\ : std_logic;
signal \SIG_DDS.tmp_buf_3\ : std_logic;
signal \SIG_DDS.tmp_buf_4\ : std_logic;
signal \SIG_DDS.tmp_buf_5\ : std_logic;
signal \SIG_DDS.tmp_buf_6\ : std_logic;
signal \ADC_VDC.genclk.t0on_0\ : std_logic;
signal \bfn_15_3_0_\ : std_logic;
signal \ADC_VDC.genclk.t0on_1\ : std_logic;
signal \ADC_VDC.genclk.n19425\ : std_logic;
signal \ADC_VDC.genclk.t0on_2\ : std_logic;
signal \ADC_VDC.genclk.n19426\ : std_logic;
signal \ADC_VDC.genclk.t0on_3\ : std_logic;
signal \ADC_VDC.genclk.n19427\ : std_logic;
signal \ADC_VDC.genclk.t0on_4\ : std_logic;
signal \ADC_VDC.genclk.n19428\ : std_logic;
signal \ADC_VDC.genclk.t0on_5\ : std_logic;
signal \ADC_VDC.genclk.n19429\ : std_logic;
signal \ADC_VDC.genclk.t0on_6\ : std_logic;
signal \ADC_VDC.genclk.n19430\ : std_logic;
signal \ADC_VDC.genclk.t0on_7\ : std_logic;
signal \ADC_VDC.genclk.n19431\ : std_logic;
signal \ADC_VDC.genclk.n19432\ : std_logic;
signal \INVADC_VDC.genclk.t0on_i0C_net\ : std_logic;
signal \ADC_VDC.genclk.t0on_8\ : std_logic;
signal \bfn_15_4_0_\ : std_logic;
signal \ADC_VDC.genclk.t0on_9\ : std_logic;
signal \ADC_VDC.genclk.n19433\ : std_logic;
signal \ADC_VDC.genclk.t0on_10\ : std_logic;
signal \ADC_VDC.genclk.n19434\ : std_logic;
signal \ADC_VDC.genclk.t0on_11\ : std_logic;
signal \ADC_VDC.genclk.n19435\ : std_logic;
signal \ADC_VDC.genclk.t0on_12\ : std_logic;
signal \ADC_VDC.genclk.n19436\ : std_logic;
signal \ADC_VDC.genclk.t0on_13\ : std_logic;
signal \ADC_VDC.genclk.n19437\ : std_logic;
signal \ADC_VDC.genclk.t0on_14\ : std_logic;
signal \ADC_VDC.genclk.n19438\ : std_logic;
signal \ADC_VDC.genclk.n19439\ : std_logic;
signal \ADC_VDC.genclk.t0on_15\ : std_logic;
signal \INVADC_VDC.genclk.t0on_i8C_net\ : std_logic;
signal \ADC_VDC.genclk.div_state_1__N_1266\ : std_logic;
signal \ADC_VDC.genclk.n14695\ : std_logic;
signal \comm_spi.n14585\ : std_logic;
signal \INVcomm_spi.MISO_48_12187_12188_setC_net\ : std_logic;
signal comm_tx_buf_7 : std_logic;
signal comm_tx_buf_2 : std_logic;
signal \comm_spi.imosi_N_744\ : std_logic;
signal \ICE_SPI_MOSI\ : std_logic;
signal \comm_spi.imosi_N_745\ : std_logic;
signal \comm_spi.n22644\ : std_logic;
signal \comm_spi.data_tx_7__N_778\ : std_logic;
signal \comm_spi.n14608\ : std_logic;
signal \comm_spi.data_tx_7__N_781\ : std_logic;
signal \comm_spi.n14607\ : std_logic;
signal \comm_spi.data_tx_7__N_763\ : std_logic;
signal comm_tx_buf_3 : std_logic;
signal eis_state_0 : std_logic;
signal n21067 : std_logic;
signal n10508 : std_logic;
signal \n11839_cascade_\ : std_logic;
signal n9222 : std_logic;
signal \n9222_cascade_\ : std_logic;
signal \n24_adj_1579_cascade_\ : std_logic;
signal \n21079_cascade_\ : std_logic;
signal n12643 : std_logic;
signal n16_adj_1570 : std_logic;
signal \n12080_cascade_\ : std_logic;
signal comm_buf_4_0 : std_logic;
signal n22132 : std_logic;
signal n12206 : std_logic;
signal \n12206_cascade_\ : std_logic;
signal n14770 : std_logic;
signal comm_buf_6_0 : std_logic;
signal comm_buf_2_0 : std_logic;
signal n22129 : std_logic;
signal buf_data_iac_5 : std_logic;
signal \n22_adj_1599_cascade_\ : std_logic;
signal \n30_adj_1600_cascade_\ : std_logic;
signal comm_rx_buf_5 : std_logic;
signal n12080 : std_logic;
signal n14749 : std_logic;
signal buf_adcdata_vdc_5 : std_logic;
signal buf_adcdata_vac_5 : std_logic;
signal n19_adj_1598 : std_logic;
signal comm_buf_2_5 : std_logic;
signal comm_buf_6_5 : std_logic;
signal comm_buf_4_5 : std_logic;
signal \n22123_cascade_\ : std_logic;
signal n22126 : std_logic;
signal n20602 : std_logic;
signal \SELIRNG0\ : std_logic;
signal n14_adj_1552 : std_logic;
signal \n14_adj_1552_cascade_\ : std_logic;
signal n14_adj_1550 : std_logic;
signal n12254 : std_logic;
signal n12007 : std_logic;
signal n14_adj_1527 : std_logic;
signal n14_adj_1529 : std_logic;
signal req_data_cnt_5 : std_logic;
signal req_data_cnt_4 : std_logic;
signal req_data_cnt_1 : std_logic;
signal n20_adj_1496 : std_logic;
signal \n18_adj_1553_cascade_\ : std_logic;
signal eis_stop : std_logic;
signal \n29_cascade_\ : std_logic;
signal n16_adj_1609 : std_logic;
signal n14_adj_1558 : std_logic;
signal req_data_cnt_3 : std_logic;
signal acadc_skipcnt_12 : std_logic;
signal acadc_skipcnt_10 : std_logic;
signal n21 : std_logic;
signal \n9_adj_1408_cascade_\ : std_logic;
signal cmd_rdadctmp_14_adj_1429 : std_logic;
signal comm_buf_0_2 : std_logic;
signal \acadc_skipCount_10\ : std_logic;
signal n12391 : std_logic;
signal n12367 : std_logic;
signal n11324 : std_logic;
signal \n8780_cascade_\ : std_logic;
signal eis_state_1 : std_logic;
signal buf_dds0_7 : std_logic;
signal n8_adj_1541 : std_logic;
signal \n8_adj_1541_cascade_\ : std_logic;
signal \data_index_9_N_212_4\ : std_logic;
signal data_count_0 : std_logic;
signal \bfn_15_17_0_\ : std_logic;
signal data_count_1 : std_logic;
signal n19287 : std_logic;
signal data_count_2 : std_logic;
signal n19288 : std_logic;
signal data_count_3 : std_logic;
signal n19289 : std_logic;
signal data_count_4 : std_logic;
signal n19290 : std_logic;
signal data_count_5 : std_logic;
signal n19291 : std_logic;
signal data_count_6 : std_logic;
signal n19292 : std_logic;
signal data_count_7 : std_logic;
signal n19293 : std_logic;
signal n19294 : std_logic;
signal \INVdata_count_i0_i0C_net\ : std_logic;
signal data_count_8 : std_logic;
signal \bfn_15_18_0_\ : std_logic;
signal n19295 : std_logic;
signal data_count_9 : std_logic;
signal \INVdata_count_i0_i8C_net\ : std_logic;
signal \SIG_DDS.tmp_buf_14\ : std_logic;
signal buf_dds0_0 : std_logic;
signal \SIG_DDS.tmp_buf_0\ : std_logic;
signal \SIG_DDS.n12700\ : std_logic;
signal comm_tx_buf_6 : std_logic;
signal \comm_spi.data_tx_7__N_758\ : std_logic;
signal \comm_spi.n22623\ : std_logic;
signal \comm_spi.n14592\ : std_logic;
signal \comm_spi.n14593\ : std_logic;
signal \INVcomm_spi.imiso_83_12193_12194_resetC_net\ : std_logic;
signal n17393 : std_logic;
signal n30 : std_logic;
signal \comm_state_3_N_412_3_cascade_\ : std_logic;
signal \n20700_cascade_\ : std_logic;
signal flagcntwd : std_logic;
signal n11411 : std_logic;
signal n20081 : std_logic;
signal n11333 : std_logic;
signal comm_buf_0_6 : std_logic;
signal n28 : std_logic;
signal n27 : std_logic;
signal \n26_adj_1625_cascade_\ : std_logic;
signal n25_adj_1616 : std_logic;
signal \n19553_cascade_\ : std_logic;
signal n22_adj_1594 : std_logic;
signal n10_adj_1582 : std_logic;
signal clk_cnt_1 : std_logic;
signal clk_cnt_0 : std_logic;
signal \clk_RTD\ : std_logic;
signal \TEST_LED\ : std_logic;
signal buf_adcdata_vdc_6 : std_logic;
signal buf_adcdata_vac_6 : std_logic;
signal n19_adj_1593 : std_logic;
signal n21071 : std_logic;
signal n20_adj_1607 : std_logic;
signal comm_buf_5_4 : std_logic;
signal comm_buf_4_4 : std_logic;
signal data_idxvec_8 : std_logic;
signal n20779 : std_logic;
signal \n12415_cascade_\ : std_logic;
signal \buf_cfgRTD_5\ : std_logic;
signal comm_buf_1_0 : std_logic;
signal n14_adj_1528 : std_logic;
signal n14_adj_1525 : std_logic;
signal n20850 : std_logic;
signal n30_adj_1520 : std_logic;
signal n14_adj_1524 : std_logic;
signal req_data_cnt_0 : std_logic;
signal req_data_cnt_6 : std_logic;
signal n17_adj_1554 : std_logic;
signal req_data_cnt_15 : std_logic;
signal req_data_cnt_9 : std_logic;
signal n20613 : std_logic;
signal req_data_cnt_2 : std_logic;
signal req_data_cnt_7 : std_logic;
signal n14_adj_1548 : std_logic;
signal n22_adj_1492 : std_logic;
signal \n21_adj_1494_cascade_\ : std_logic;
signal n24_adj_1530 : std_logic;
signal n30_adj_1597 : std_logic;
signal n14_adj_1549 : std_logic;
signal \buf_cfgRTD_4\ : std_logic;
signal n12415 : std_logic;
signal n14_adj_1551 : std_logic;
signal req_data_cnt_10 : std_logic;
signal req_data_cnt_8 : std_logic;
signal n19_adj_1499 : std_logic;
signal \bfn_16_15_0_\ : std_logic;
signal n19326 : std_logic;
signal data_index_2 : std_logic;
signal n7_adj_1544 : std_logic;
signal n19327 : std_logic;
signal data_index_3 : std_logic;
signal n7_adj_1542 : std_logic;
signal n19328 : std_logic;
signal data_index_4 : std_logic;
signal n7_adj_1540 : std_logic;
signal n19329 : std_logic;
signal n19330 : std_logic;
signal n19331 : std_logic;
signal data_index_7 : std_logic;
signal n7_adj_1535 : std_logic;
signal n19332 : std_logic;
signal n19333 : std_logic;
signal data_index_8 : std_logic;
signal n7_adj_1533 : std_logic;
signal \bfn_16_16_0_\ : std_logic;
signal n10579 : std_logic;
signal n19334 : std_logic;
signal \n17338_cascade_\ : std_logic;
signal \data_index_9_N_212_5\ : std_logic;
signal n7_adj_1515 : std_logic;
signal n17314 : std_logic;
signal data_index_0 : std_logic;
signal comm_buf_1_2 : std_logic;
signal buf_dds0_2 : std_logic;
signal data_index_9 : std_logic;
signal buf_dds0_4 : std_logic;
signal \n8_adj_1538_cascade_\ : std_logic;
signal data_index_6 : std_logic;
signal buf_dds0_6 : std_logic;
signal comm_buf_1_7 : std_logic;
signal buf_dds1_7 : std_logic;
signal comm_buf_0_0 : std_logic;
signal buf_dds0_8 : std_logic;
signal comm_buf_1_1 : std_logic;
signal data_index_1 : std_logic;
signal n8780 : std_logic;
signal n8_adj_1547 : std_logic;
signal \n8_adj_1547_cascade_\ : std_logic;
signal n7_adj_1546 : std_logic;
signal \data_index_9_N_212_1\ : std_logic;
signal buf_dds0_11 : std_logic;
signal buf_dds0_5 : std_logic;
signal n8_adj_1532 : std_logic;
signal n7_adj_1531 : std_logic;
signal \data_index_9_N_212_9\ : std_logic;
signal tmp_buf_15 : std_logic;
signal \DDS_MOSI\ : std_logic;
signal comm_buf_0_1 : std_logic;
signal \DDS_RNG_0\ : std_logic;
signal n8_adj_1538 : std_logic;
signal n7_adj_1537 : std_logic;
signal \data_index_9_N_212_6\ : std_logic;
signal n11901 : std_logic;
signal comm_buf_0_3 : std_logic;
signal n14869 : std_logic;
signal bit_cnt_0 : std_logic;
signal \comm_spi.n14624\ : std_logic;
signal \comm_spi.data_tx_7__N_769\ : std_logic;
signal \comm_spi.n22626\ : std_logic;
signal \comm_spi.n22626_cascade_\ : std_logic;
signal \comm_spi.n14589\ : std_logic;
signal \ICE_SPI_MISO\ : std_logic;
signal \comm_spi.n22635\ : std_logic;
signal \comm_spi.n14623\ : std_logic;
signal \comm_spi.data_tx_7__N_759\ : std_logic;
signal \comm_spi.n14596\ : std_logic;
signal \comm_spi.n14595\ : std_logic;
signal \comm_spi.n14588\ : std_logic;
signal \comm_spi.n14590\ : std_logic;
signal \INVcomm_spi.MISO_48_12187_12188_resetC_net\ : std_logic;
signal \comm_spi.data_tx_7__N_766\ : std_logic;
signal n20931 : std_logic;
signal \n21913_cascade_\ : std_logic;
signal n21916 : std_logic;
signal \n1252_cascade_\ : std_logic;
signal n2 : std_logic;
signal \n21088_cascade_\ : std_logic;
signal n14_adj_1497 : std_logic;
signal \comm_state_3_N_412_3\ : std_logic;
signal n1252 : std_logic;
signal n8_adj_1555 : std_logic;
signal \n2342_cascade_\ : std_logic;
signal \comm_state_3_N_428_2\ : std_logic;
signal \n15_adj_1602_cascade_\ : std_logic;
signal n20571 : std_logic;
signal \n20641_cascade_\ : std_logic;
signal n12_adj_1603 : std_logic;
signal n7_adj_1588 : std_logic;
signal secclk_cnt_0 : std_logic;
signal \bfn_17_9_0_\ : std_logic;
signal secclk_cnt_1 : std_logic;
signal n19447 : std_logic;
signal secclk_cnt_2 : std_logic;
signal n19448 : std_logic;
signal secclk_cnt_3 : std_logic;
signal n19449 : std_logic;
signal secclk_cnt_4 : std_logic;
signal n19450 : std_logic;
signal secclk_cnt_5 : std_logic;
signal n19451 : std_logic;
signal secclk_cnt_6 : std_logic;
signal n19452 : std_logic;
signal secclk_cnt_7 : std_logic;
signal n19453 : std_logic;
signal n19454 : std_logic;
signal secclk_cnt_8 : std_logic;
signal \bfn_17_10_0_\ : std_logic;
signal secclk_cnt_9 : std_logic;
signal n19455 : std_logic;
signal secclk_cnt_10 : std_logic;
signal n19456 : std_logic;
signal secclk_cnt_11 : std_logic;
signal n19457 : std_logic;
signal n19458 : std_logic;
signal secclk_cnt_13 : std_logic;
signal n19459 : std_logic;
signal secclk_cnt_14 : std_logic;
signal n19460 : std_logic;
signal secclk_cnt_15 : std_logic;
signal n19461 : std_logic;
signal n19462 : std_logic;
signal secclk_cnt_16 : std_logic;
signal \bfn_17_11_0_\ : std_logic;
signal secclk_cnt_17 : std_logic;
signal n19463 : std_logic;
signal secclk_cnt_18 : std_logic;
signal n19464 : std_logic;
signal n19465 : std_logic;
signal secclk_cnt_20 : std_logic;
signal n19466 : std_logic;
signal n19467 : std_logic;
signal n19468 : std_logic;
signal n14700 : std_logic;
signal comm_buf_0_5 : std_logic;
signal n14_adj_1556 : std_logic;
signal \VDC_RNG0\ : std_logic;
signal \acadc_skipCount_12\ : std_logic;
signal req_data_cnt_13 : std_logic;
signal n21022 : std_logic;
signal n21049 : std_logic;
signal comm_length_2 : std_logic;
signal \n21955_cascade_\ : std_logic;
signal n21958 : std_logic;
signal n21024 : std_logic;
signal buf_data_iac_19 : std_logic;
signal n20950 : std_logic;
signal data_idxvec_11 : std_logic;
signal n26_adj_1519 : std_logic;
signal \SELIRNG1\ : std_logic;
signal \acadc_skipCount_11\ : std_logic;
signal n23_adj_1518 : std_logic;
signal comm_length_0 : std_logic;
signal n11846 : std_logic;
signal n14652 : std_logic;
signal n10553 : std_logic;
signal n20622 : std_logic;
signal n12381 : std_logic;
signal req_data_cnt_11 : std_logic;
signal req_data_cnt_14 : std_logic;
signal n23_adj_1491 : std_logic;
signal cmd_rdadctmp_15_adj_1428 : std_logic;
signal cmd_rdadctmp_15 : std_logic;
signal cmd_rdadctmp_16 : std_logic;
signal n17338 : std_logic;
signal n17336 : std_logic;
signal data_index_5 : std_logic;
signal n16708 : std_logic;
signal n20626 : std_logic;
signal n11805 : std_logic;
signal n14_adj_1523 : std_logic;
signal n12353 : std_logic;
signal buf_dds0_15 : std_logic;
signal n9 : std_logic;
signal \SIG_DDS.n9\ : std_logic;
signal \comm_spi.n14620\ : std_logic;
signal \comm_spi.data_tx_7__N_772\ : std_logic;
signal \comm_spi.n22638\ : std_logic;
signal \comm_spi.n14619\ : std_logic;
signal \comm_spi.n14615\ : std_logic;
signal \comm_spi.data_tx_7__N_761\ : std_logic;
signal \comm_spi.n22641\ : std_logic;
signal \comm_spi.n14611\ : std_logic;
signal \comm_spi.n14612\ : std_logic;
signal \comm_spi.n14616\ : std_logic;
signal n20641 : std_logic;
signal n17656 : std_logic;
signal n21162 : std_logic;
signal \n17658_cascade_\ : std_logic;
signal n20653 : std_logic;
signal \n12220_cascade_\ : std_logic;
signal \n4_adj_1483_cascade_\ : std_logic;
signal n12205 : std_logic;
signal n4 : std_logic;
signal \n20510_cascade_\ : std_logic;
signal n3 : std_logic;
signal n20534 : std_logic;
signal n11810 : std_logic;
signal \n11810_cascade_\ : std_logic;
signal n20650 : std_logic;
signal \n20672_cascade_\ : std_logic;
signal n20510 : std_logic;
signal n20585 : std_logic;
signal n11824 : std_logic;
signal \comm_spi.bit_cnt_3\ : std_logic;
signal \comm_spi.n16858\ : std_logic;
signal \INVcomm_spi.data_valid_85C_net\ : std_logic;
signal n21087 : std_logic;
signal n4_adj_1566 : std_logic;
signal \n22063_cascade_\ : std_logic;
signal comm_buf_6_4 : std_logic;
signal n21081 : std_logic;
signal comm_buf_0_4 : std_logic;
signal comm_buf_1_4 : std_logic;
signal n1_adj_1564 : std_logic;
signal \n18824_cascade_\ : std_logic;
signal n20507 : std_logic;
signal comm_buf_2_4 : std_logic;
signal comm_buf_3_4 : std_logic;
signal n2_adj_1565 : std_logic;
signal comm_buf_5_1 : std_logic;
signal comm_buf_4_1 : std_logic;
signal \n4_adj_1569_cascade_\ : std_logic;
signal comm_buf_6_1 : std_logic;
signal \n20792_cascade_\ : std_logic;
signal n21994 : std_logic;
signal n12322 : std_logic;
signal n14784 : std_logic;
signal n21069 : std_logic;
signal \iac_raw_buf_N_728\ : std_logic;
signal data_cntvec_0 : std_logic;
signal \bfn_18_12_0_\ : std_logic;
signal data_cntvec_1 : std_logic;
signal n19296 : std_logic;
signal data_cntvec_2 : std_logic;
signal n19297 : std_logic;
signal data_cntvec_3 : std_logic;
signal n19298 : std_logic;
signal data_cntvec_4 : std_logic;
signal n19299 : std_logic;
signal data_cntvec_5 : std_logic;
signal n19300 : std_logic;
signal data_cntvec_6 : std_logic;
signal n19301 : std_logic;
signal data_cntvec_7 : std_logic;
signal n19302 : std_logic;
signal n19303 : std_logic;
signal \INVdata_cntvec_i0_i0C_net\ : std_logic;
signal data_cntvec_8 : std_logic;
signal \bfn_18_13_0_\ : std_logic;
signal data_cntvec_9 : std_logic;
signal n19304 : std_logic;
signal data_cntvec_10 : std_logic;
signal n19305 : std_logic;
signal data_cntvec_11 : std_logic;
signal n19306 : std_logic;
signal data_cntvec_12 : std_logic;
signal n19307 : std_logic;
signal data_cntvec_13 : std_logic;
signal n19308 : std_logic;
signal data_cntvec_14 : std_logic;
signal n19309 : std_logic;
signal n19310 : std_logic;
signal data_cntvec_15 : std_logic;
signal \INVdata_cntvec_i0_i8C_net\ : std_logic;
signal n13443 : std_logic;
signal n14632 : std_logic;
signal buf_adcdata_iac_6 : std_logic;
signal n20540 : std_logic;
signal adc_state_0_adj_1411 : std_logic;
signal cmd_rdadctmp_12_adj_1431 : std_logic;
signal buf_adcdata_vac_7 : std_logic;
signal buf_adcdata_vdc_7 : std_logic;
signal buf_adcdata_iac_7 : std_logic;
signal \n19_adj_1589_cascade_\ : std_logic;
signal comm_cmd_2 : std_logic;
signal buf_data_iac_7 : std_logic;
signal \n22_adj_1590_cascade_\ : std_logic;
signal n30_adj_1591 : std_logic;
signal buf_adcdata_iac_5 : std_logic;
signal cmd_rdadctmp_11 : std_logic;
signal n20543 : std_logic;
signal buf_adcdata_iac_4 : std_logic;
signal cmd_rdadctmp_14 : std_logic;
signal \comm_spi.n14581\ : std_logic;
signal \comm_spi.iclk_N_754\ : std_logic;
signal comm_tx_buf_5 : std_logic;
signal \comm_spi.data_tx_7__N_760\ : std_logic;
signal \ICE_GPMI_0\ : std_logic;
signal n11406 : std_logic;
signal n12220 : std_logic;
signal \n10_adj_1572_cascade_\ : std_logic;
signal n20643 : std_logic;
signal n4_adj_1596 : std_logic;
signal n2342 : std_logic;
signal n11836 : std_logic;
signal n14722 : std_logic;
signal \comm_spi.n22647\ : std_logic;
signal comm_buf_1_5 : std_logic;
signal n14_adj_1557 : std_logic;
signal comm_index_2 : std_logic;
signal n18824 : std_logic;
signal \n20563_cascade_\ : std_logic;
signal n20627 : std_logic;
signal \n12_adj_1539_cascade_\ : std_logic;
signal n20556 : std_logic;
signal n12164 : std_logic;
signal \ICE_SPI_CE0\ : std_logic;
signal comm_data_vld : std_logic;
signal n23_adj_1574 : std_logic;
signal \n21_adj_1573_cascade_\ : std_logic;
signal n18 : std_logic;
signal comm_index_1 : std_logic;
signal comm_length_1 : std_logic;
signal n4_adj_1576 : std_logic;
signal comm_cmd_7 : std_logic;
signal \n5_cascade_\ : std_logic;
signal n20863 : std_logic;
signal n14514 : std_logic;
signal \n21658_cascade_\ : std_logic;
signal n9273 : std_logic;
signal \n20865_cascade_\ : std_logic;
signal n20536 : std_logic;
signal n10540 : std_logic;
signal comm_index_0 : std_logic;
signal n20563 : std_logic;
signal n12_adj_1585 : std_logic;
signal comm_buf_1_6 : std_logic;
signal n14_adj_1526 : std_logic;
signal buf_adcdata_vdc_4 : std_logic;
signal buf_adcdata_vac_4 : std_logic;
signal n19_adj_1605 : std_logic;
signal comm_state_2 : std_logic;
signal n20734 : std_logic;
signal adc_state_0 : std_logic;
signal cmd_rdadctmp_12 : std_logic;
signal n12542 : std_logic;
signal cmd_rdadctmp_13 : std_logic;
signal buf_control_0 : std_logic;
signal wdtick_flag : std_logic;
signal \CONT_SD\ : std_logic;
signal trig_dds0 : std_logic;
signal \comm_spi.n14582\ : std_logic;
signal \ICE_SPI_SCLK\ : std_logic;
signal \comm_spi.iclk_N_755\ : std_logic;
signal \comm_spi.data_tx_7__N_765\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \comm_spi.data_tx_7__N_787\ : std_logic;
signal \comm_spi.n14604\ : std_logic;
signal \comm_spi.n14578\ : std_logic;
signal \comm_spi.n14577\ : std_logic;
signal \comm_spi.n14603\ : std_logic;
signal \comm_spi.iclk\ : std_logic;
signal comm_tx_buf_0 : std_logic;
signal \comm_spi.n22650\ : std_logic;
signal \comm_spi.data_tx_7__N_764\ : std_logic;
signal comm_tx_buf_1 : std_logic;
signal \comm_spi.data_tx_7__N_784\ : std_logic;
signal comm_tx_buf_4 : std_logic;
signal \comm_spi.data_tx_7__N_775\ : std_logic;
signal \n20502_cascade_\ : std_logic;
signal n12_adj_1583 : std_logic;
signal n20502 : std_logic;
signal \INVdds0_mclk_294C_net\ : std_logic;
signal secclk_cnt_19 : std_logic;
signal secclk_cnt_21 : std_logic;
signal secclk_cnt_12 : std_logic;
signal secclk_cnt_22 : std_logic;
signal n14_adj_1578 : std_logic;
signal comm_cmd_1 : std_logic;
signal comm_cmd_0 : std_logic;
signal n23_adj_1517 : std_logic;
signal req_data_cnt_12 : std_logic;
signal n20809 : std_logic;
signal n17415 : std_logic;
signal buf_data_iac_4 : std_logic;
signal comm_cmd_3 : std_logic;
signal n22_adj_1606 : std_logic;
signal n30_adj_1608 : std_logic;
signal \clk_16MHz\ : std_logic;
signal dds0_mclk : std_logic;
signal buf_control_6 : std_logic;
signal \DDS_MCLK\ : std_logic;
signal \DDS_SCK\ : std_logic;
signal dds_state_2 : std_logic;
signal dds_state_0 : std_logic;
signal dds_state_1 : std_logic;
signal \DDS_CS\ : std_logic;
signal \SIG_DDS.n9_adj_1385\ : std_logic;
signal comm_clear : std_logic;
signal \clk_32MHz\ : std_logic;
signal comm_state_3 : std_logic;
signal comm_state_1 : std_logic;
signal comm_state_0 : std_logic;
signal n11347 : std_logic;
signal dds0_mclkcnt_0 : std_logic;
signal \bfn_22_11_0_\ : std_logic;
signal dds0_mclkcnt_1 : std_logic;
signal n19440 : std_logic;
signal dds0_mclkcnt_2 : std_logic;
signal n19441 : std_logic;
signal dds0_mclkcnt_3 : std_logic;
signal n19442 : std_logic;
signal dds0_mclkcnt_4 : std_logic;
signal n19443 : std_logic;
signal dds0_mclkcnt_5 : std_logic;
signal n19444 : std_logic;
signal n10 : std_logic;
signal dds0_mclkcnt_6 : std_logic;
signal n19445 : std_logic;
signal n19446 : std_logic;
signal dds0_mclkcnt_7 : std_logic;
signal \INVdds0_mclkcnt_i7_3772__i0C_net\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \VAC_DRDY_wire\ : std_logic;
signal \IAC_FLT1_wire\ : std_logic;
signal \DDS_SCK_wire\ : std_logic;
signal \ICE_IOR_166_wire\ : std_logic;
signal \ICE_IOR_119_wire\ : std_logic;
signal \DDS_MOSI_wire\ : std_logic;
signal \VAC_MISO_wire\ : std_logic;
signal \DDS_MOSI1_wire\ : std_logic;
signal \ICE_IOR_146_wire\ : std_logic;
signal \VDC_CLK_wire\ : std_logic;
signal \ICE_IOT_222_wire\ : std_logic;
signal \IAC_CS_wire\ : std_logic;
signal \ICE_IOL_18B_wire\ : std_logic;
signal \ICE_IOL_13A_wire\ : std_logic;
signal \ICE_IOB_81_wire\ : std_logic;
signal \VAC_OSR1_wire\ : std_logic;
signal \IAC_MOSI_wire\ : std_logic;
signal \DDS_CS1_wire\ : std_logic;
signal \ICE_IOL_4B_wire\ : std_logic;
signal \ICE_IOB_94_wire\ : std_logic;
signal \VAC_CS_wire\ : std_logic;
signal \VAC_CLK_wire\ : std_logic;
signal \ICE_SPI_CE0_wire\ : std_logic;
signal \ICE_IOR_167_wire\ : std_logic;
signal \ICE_IOR_118_wire\ : std_logic;
signal \RTD_SDO_wire\ : std_logic;
signal \IAC_OSR0_wire\ : std_logic;
signal \VDC_SCLK_wire\ : std_logic;
signal \VAC_FLT1_wire\ : std_logic;
signal \ICE_SPI_MOSI_wire\ : std_logic;
signal \ICE_IOR_165_wire\ : std_logic;
signal \ICE_IOR_147_wire\ : std_logic;
signal \ICE_IOL_14A_wire\ : std_logic;
signal \ICE_IOL_13B_wire\ : std_logic;
signal \ICE_IOB_91_wire\ : std_logic;
signal \ICE_GPMO_0_wire\ : std_logic;
signal \DDS_RNG_0_wire\ : std_logic;
signal \VDC_RNG0_wire\ : std_logic;
signal \ICE_SPI_SCLK_wire\ : std_logic;
signal \ICE_IOR_152_wire\ : std_logic;
signal \ICE_IOL_12A_wire\ : std_logic;
signal \RTD_DRDY_wire\ : std_logic;
signal \ICE_SPI_MISO_wire\ : std_logic;
signal \ICE_IOT_177_wire\ : std_logic;
signal \ICE_IOR_141_wire\ : std_logic;
signal \ICE_IOB_80_wire\ : std_logic;
signal \ICE_IOB_102_wire\ : std_logic;
signal \ICE_GPMO_2_wire\ : std_logic;
signal \ICE_GPMI_0_wire\ : std_logic;
signal \IAC_MISO_wire\ : std_logic;
signal \VAC_OSR0_wire\ : std_logic;
signal \VAC_MOSI_wire\ : std_logic;
signal \TEST_LED_wire\ : std_logic;
signal \ICE_IOR_148_wire\ : std_logic;
signal \STAT_COMM_wire\ : std_logic;
signal \ICE_SYSCLK_wire\ : std_logic;
signal \ICE_IOR_161_wire\ : std_logic;
signal \ICE_IOB_95_wire\ : std_logic;
signal \ICE_IOB_82_wire\ : std_logic;
signal \ICE_IOB_104_wire\ : std_logic;
signal \IAC_CLK_wire\ : std_logic;
signal \DDS_CS_wire\ : std_logic;
signal \SELIRNG0_wire\ : std_logic;
signal \RTD_SDI_wire\ : std_logic;
signal \ICE_IOT_221_wire\ : std_logic;
signal \ICE_IOT_197_wire\ : std_logic;
signal \DDS_MCLK_wire\ : std_logic;
signal \RTD_SCLK_wire\ : std_logic;
signal \RTD_CS_wire\ : std_logic;
signal \ICE_IOR_137_wire\ : std_logic;
signal \IAC_OSR1_wire\ : std_logic;
signal \VAC_FLT0_wire\ : std_logic;
signal \ICE_IOR_144_wire\ : std_logic;
signal \ICE_IOR_128_wire\ : std_logic;
signal \ICE_GPMO_1_wire\ : std_logic;
signal \IAC_SCLK_wire\ : std_logic;
signal \EIS_SYNCCLK_wire\ : std_logic;
signal \ICE_IOR_139_wire\ : std_logic;
signal \ICE_IOL_4A_wire\ : std_logic;
signal \VAC_SCLK_wire\ : std_logic;
signal \THERMOSTAT_wire\ : std_logic;
signal \ICE_IOR_164_wire\ : std_logic;
signal \ICE_IOB_103_wire\ : std_logic;
signal \AMPV_POW_wire\ : std_logic;
signal \VDC_SDO_wire\ : std_logic;
signal \ICE_IOT_174_wire\ : std_logic;
signal \ICE_IOR_140_wire\ : std_logic;
signal \ICE_IOB_96_wire\ : std_logic;
signal \CONT_SD_wire\ : std_logic;
signal \AC_ADC_SYNC_wire\ : std_logic;
signal \SELIRNG1_wire\ : std_logic;
signal \ICE_IOL_12B_wire\ : std_logic;
signal \ICE_IOR_160_wire\ : std_logic;
signal \ICE_IOR_136_wire\ : std_logic;
signal \DDS_MCLK1_wire\ : std_logic;
signal \ICE_IOT_198_wire\ : std_logic;
signal \ICE_IOT_173_wire\ : std_logic;
signal \IAC_DRDY_wire\ : std_logic;
signal \ICE_IOT_178_wire\ : std_logic;
signal \ICE_IOR_138_wire\ : std_logic;
signal \ICE_IOR_120_wire\ : std_logic;
signal \IAC_FLT0_wire\ : std_logic;
signal \DDS_SCK1_wire\ : std_logic;
signal \pll_main.zim_pll_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged2_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged2_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged2_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged2_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged2_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged7_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged7_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged7_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged7_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged7_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged6_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged6_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged6_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged6_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged6_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged5_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged5_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged5_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged5_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged5_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged9_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged9_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged9_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged9_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged9_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged4_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged4_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged4_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged4_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged4_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged8_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged8_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged8_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged8_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged8_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged10_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged10_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged10_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged10_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged10_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged3_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged3_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged3_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged3_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged3_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged11_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged11_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged11_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged11_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \iac_raw_buf_vac_raw_buf_merged11_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    \VAC_DRDY_wire\ <= VAC_DRDY;
    IAC_FLT1 <= \IAC_FLT1_wire\;
    DDS_SCK <= \DDS_SCK_wire\;
    \ICE_IOR_166_wire\ <= ICE_IOR_166;
    \ICE_IOR_119_wire\ <= ICE_IOR_119;
    DDS_MOSI <= \DDS_MOSI_wire\;
    \VAC_MISO_wire\ <= VAC_MISO;
    DDS_MOSI1 <= \DDS_MOSI1_wire\;
    \ICE_IOR_146_wire\ <= ICE_IOR_146;
    VDC_CLK <= \VDC_CLK_wire\;
    \ICE_IOT_222_wire\ <= ICE_IOT_222;
    IAC_CS <= \IAC_CS_wire\;
    \ICE_IOL_18B_wire\ <= ICE_IOL_18B;
    \ICE_IOL_13A_wire\ <= ICE_IOL_13A;
    \ICE_IOB_81_wire\ <= ICE_IOB_81;
    VAC_OSR1 <= \VAC_OSR1_wire\;
    IAC_MOSI <= \IAC_MOSI_wire\;
    DDS_CS1 <= \DDS_CS1_wire\;
    \ICE_IOL_4B_wire\ <= ICE_IOL_4B;
    \ICE_IOB_94_wire\ <= ICE_IOB_94;
    VAC_CS <= \VAC_CS_wire\;
    VAC_CLK <= \VAC_CLK_wire\;
    \ICE_SPI_CE0_wire\ <= ICE_SPI_CE0;
    \ICE_IOR_167_wire\ <= ICE_IOR_167;
    \ICE_IOR_118_wire\ <= ICE_IOR_118;
    \RTD_SDO_wire\ <= RTD_SDO;
    IAC_OSR0 <= \IAC_OSR0_wire\;
    VDC_SCLK <= \VDC_SCLK_wire\;
    VAC_FLT1 <= \VAC_FLT1_wire\;
    \ICE_SPI_MOSI_wire\ <= ICE_SPI_MOSI;
    \ICE_IOR_165_wire\ <= ICE_IOR_165;
    \ICE_IOR_147_wire\ <= ICE_IOR_147;
    \ICE_IOL_14A_wire\ <= ICE_IOL_14A;
    \ICE_IOL_13B_wire\ <= ICE_IOL_13B;
    \ICE_IOB_91_wire\ <= ICE_IOB_91;
    \ICE_GPMO_0_wire\ <= ICE_GPMO_0;
    DDS_RNG_0 <= \DDS_RNG_0_wire\;
    VDC_RNG0 <= \VDC_RNG0_wire\;
    \ICE_SPI_SCLK_wire\ <= ICE_SPI_SCLK;
    \ICE_IOR_152_wire\ <= ICE_IOR_152;
    \ICE_IOL_12A_wire\ <= ICE_IOL_12A;
    \RTD_DRDY_wire\ <= RTD_DRDY;
    ICE_SPI_MISO <= \ICE_SPI_MISO_wire\;
    \ICE_IOT_177_wire\ <= ICE_IOT_177;
    \ICE_IOR_141_wire\ <= ICE_IOR_141;
    \ICE_IOB_80_wire\ <= ICE_IOB_80;
    \ICE_IOB_102_wire\ <= ICE_IOB_102;
    \ICE_GPMO_2_wire\ <= ICE_GPMO_2;
    ICE_GPMI_0 <= \ICE_GPMI_0_wire\;
    \IAC_MISO_wire\ <= IAC_MISO;
    VAC_OSR0 <= \VAC_OSR0_wire\;
    VAC_MOSI <= \VAC_MOSI_wire\;
    TEST_LED <= \TEST_LED_wire\;
    \ICE_IOR_148_wire\ <= ICE_IOR_148;
    STAT_COMM <= \STAT_COMM_wire\;
    \ICE_SYSCLK_wire\ <= ICE_SYSCLK;
    \ICE_IOR_161_wire\ <= ICE_IOR_161;
    \ICE_IOB_95_wire\ <= ICE_IOB_95;
    \ICE_IOB_82_wire\ <= ICE_IOB_82;
    \ICE_IOB_104_wire\ <= ICE_IOB_104;
    IAC_CLK <= \IAC_CLK_wire\;
    DDS_CS <= \DDS_CS_wire\;
    SELIRNG0 <= \SELIRNG0_wire\;
    RTD_SDI <= \RTD_SDI_wire\;
    \ICE_IOT_221_wire\ <= ICE_IOT_221;
    \ICE_IOT_197_wire\ <= ICE_IOT_197;
    DDS_MCLK <= \DDS_MCLK_wire\;
    RTD_SCLK <= \RTD_SCLK_wire\;
    RTD_CS <= \RTD_CS_wire\;
    \ICE_IOR_137_wire\ <= ICE_IOR_137;
    IAC_OSR1 <= \IAC_OSR1_wire\;
    VAC_FLT0 <= \VAC_FLT0_wire\;
    \ICE_IOR_144_wire\ <= ICE_IOR_144;
    \ICE_IOR_128_wire\ <= ICE_IOR_128;
    \ICE_GPMO_1_wire\ <= ICE_GPMO_1;
    IAC_SCLK <= \IAC_SCLK_wire\;
    \EIS_SYNCCLK_wire\ <= EIS_SYNCCLK;
    \ICE_IOR_139_wire\ <= ICE_IOR_139;
    \ICE_IOL_4A_wire\ <= ICE_IOL_4A;
    VAC_SCLK <= \VAC_SCLK_wire\;
    \THERMOSTAT_wire\ <= THERMOSTAT;
    \ICE_IOR_164_wire\ <= ICE_IOR_164;
    \ICE_IOB_103_wire\ <= ICE_IOB_103;
    AMPV_POW <= \AMPV_POW_wire\;
    \VDC_SDO_wire\ <= VDC_SDO;
    \ICE_IOT_174_wire\ <= ICE_IOT_174;
    \ICE_IOR_140_wire\ <= ICE_IOR_140;
    \ICE_IOB_96_wire\ <= ICE_IOB_96;
    CONT_SD <= \CONT_SD_wire\;
    AC_ADC_SYNC <= \AC_ADC_SYNC_wire\;
    SELIRNG1 <= \SELIRNG1_wire\;
    \ICE_IOL_12B_wire\ <= ICE_IOL_12B;
    \ICE_IOR_160_wire\ <= ICE_IOR_160;
    \ICE_IOR_136_wire\ <= ICE_IOR_136;
    DDS_MCLK1 <= \DDS_MCLK1_wire\;
    \ICE_IOT_198_wire\ <= ICE_IOT_198;
    \ICE_IOT_173_wire\ <= ICE_IOT_173;
    \IAC_DRDY_wire\ <= IAC_DRDY;
    \ICE_IOT_178_wire\ <= ICE_IOT_178;
    \ICE_IOR_138_wire\ <= ICE_IOR_138;
    \ICE_IOR_120_wire\ <= ICE_IOR_120;
    IAC_FLT0 <= \IAC_FLT0_wire\;
    DDS_SCK1 <= \DDS_SCK1_wire\;
    \pll_main.zim_pll_inst_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;
    buf_data_iac_19 <= \iac_raw_buf_vac_raw_buf_merged2_physical_RDATA_wire\(13);
    buf_data_vac_19 <= \iac_raw_buf_vac_raw_buf_merged2_physical_RDATA_wire\(9);
    buf_data_iac_18 <= \iac_raw_buf_vac_raw_buf_merged2_physical_RDATA_wire\(5);
    buf_data_vac_18 <= \iac_raw_buf_vac_raw_buf_merged2_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged2_physical_RADDR_wire\ <= '0'&\N__42985\&\N__24526\&\N__20374\&\N__43942\&\N__42238\&\N__39010\&\N__31453\&\N__36502\&\N__43183\&\N__31612\;
    \iac_raw_buf_vac_raw_buf_merged2_physical_WADDR_wire\ <= '0'&\N__40471\&\N__40579\&\N__39409\&\N__39514\&\N__39622\&\N__39730\&\N__39832\&\N__39940\&\N__40045\&\N__40150\;
    \iac_raw_buf_vac_raw_buf_merged2_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged2_physical_WDATA_wire\ <= '0'&'0'&\N__26077\&'0'&'0'&'0'&\N__21073\&'0'&'0'&'0'&\N__27811\&'0'&'0'&'0'&\N__23856\&'0';
    buf_data_iac_9 <= \iac_raw_buf_vac_raw_buf_merged7_physical_RDATA_wire\(13);
    buf_data_vac_9 <= \iac_raw_buf_vac_raw_buf_merged7_physical_RDATA_wire\(9);
    buf_data_iac_8 <= \iac_raw_buf_vac_raw_buf_merged7_physical_RDATA_wire\(5);
    buf_data_vac_8 <= \iac_raw_buf_vac_raw_buf_merged7_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged7_physical_RADDR_wire\ <= '0'&\N__42945\&\N__24480\&\N__20322\&\N__43902\&\N__42201\&\N__38970\&\N__31413\&\N__36468\&\N__43149\&\N__31578\;
    \iac_raw_buf_vac_raw_buf_merged7_physical_WADDR_wire\ <= '0'&\N__40437\&\N__40548\&\N__39369\&\N__39477\&\N__39588\&\N__39696\&\N__39792\&\N__39906\&\N__40011\&\N__40116\;
    \iac_raw_buf_vac_raw_buf_merged7_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged7_physical_WDATA_wire\ <= '0'&'0'&\N__21676\&'0'&'0'&'0'&\N__35284\&'0'&'0'&'0'&\N__24424\&'0'&'0'&'0'&\N__21397\&'0';
    buf_data_iac_21 <= \iac_raw_buf_vac_raw_buf_merged1_physical_RDATA_wire\(13);
    buf_data_vac_21 <= \iac_raw_buf_vac_raw_buf_merged1_physical_RDATA_wire\(9);
    buf_data_iac_20 <= \iac_raw_buf_vac_raw_buf_merged1_physical_RDATA_wire\(5);
    buf_data_vac_20 <= \iac_raw_buf_vac_raw_buf_merged1_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged1_physical_RADDR_wire\ <= '0'&\N__43003\&\N__24544\&\N__20392\&\N__43960\&\N__42256\&\N__39028\&\N__31471\&\N__36520\&\N__43201\&\N__31630\;
    \iac_raw_buf_vac_raw_buf_merged1_physical_WADDR_wire\ <= '0'&\N__40489\&\N__40597\&\N__39427\&\N__39532\&\N__39640\&\N__39748\&\N__39850\&\N__39958\&\N__40063\&\N__40168\;
    \iac_raw_buf_vac_raw_buf_merged1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged1_physical_WDATA_wire\ <= '0'&'0'&\N__27301\&'0'&'0'&'0'&\N__21856\&'0'&'0'&'0'&\N__28138\&'0'&'0'&'0'&\N__25711\&'0';
    buf_data_iac_11 <= \iac_raw_buf_vac_raw_buf_merged6_physical_RDATA_wire\(13);
    buf_data_vac_11 <= \iac_raw_buf_vac_raw_buf_merged6_physical_RDATA_wire\(9);
    buf_data_iac_10 <= \iac_raw_buf_vac_raw_buf_merged6_physical_RDATA_wire\(5);
    buf_data_vac_10 <= \iac_raw_buf_vac_raw_buf_merged6_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged6_physical_RADDR_wire\ <= '0'&\N__42957\&\N__24492\&\N__20334\&\N__43914\&\N__42213\&\N__38982\&\N__31425\&\N__36478\&\N__43159\&\N__31588\;
    \iac_raw_buf_vac_raw_buf_merged6_physical_WADDR_wire\ <= '0'&\N__40447\&\N__40555\&\N__39381\&\N__39489\&\N__39598\&\N__39706\&\N__39804\&\N__39916\&\N__40021\&\N__40126\;
    \iac_raw_buf_vac_raw_buf_merged6_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged6_physical_WDATA_wire\ <= '0'&'0'&\N__33533\&'0'&'0'&'0'&\N__25897\&'0'&'0'&'0'&\N__25969\&'0'&'0'&'0'&\N__24055\&'0';
    buf_data_iac_23 <= \iac_raw_buf_vac_raw_buf_merged0_physical_RDATA_wire\(13);
    buf_data_vac_23 <= \iac_raw_buf_vac_raw_buf_merged0_physical_RDATA_wire\(9);
    buf_data_iac_22 <= \iac_raw_buf_vac_raw_buf_merged0_physical_RDATA_wire\(5);
    buf_data_vac_22 <= \iac_raw_buf_vac_raw_buf_merged0_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged0_physical_RADDR_wire\ <= '0'&\N__43009\&\N__24550\&\N__20398\&\N__43966\&\N__42262\&\N__39034\&\N__31477\&\N__36526\&\N__43207\&\N__31636\;
    \iac_raw_buf_vac_raw_buf_merged0_physical_WADDR_wire\ <= '0'&\N__40495\&\N__40603\&\N__39433\&\N__39538\&\N__39646\&\N__39754\&\N__39856\&\N__39964\&\N__40069\&\N__40174\;
    \iac_raw_buf_vac_raw_buf_merged0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged0_physical_WDATA_wire\ <= '0'&'0'&\N__26275\&'0'&'0'&'0'&\N__24346\&'0'&'0'&'0'&\N__24700\&'0'&'0'&'0'&\N__22711\&'0';
    buf_data_iac_13 <= \iac_raw_buf_vac_raw_buf_merged5_physical_RDATA_wire\(13);
    buf_data_vac_13 <= \iac_raw_buf_vac_raw_buf_merged5_physical_RDATA_wire\(9);
    buf_data_iac_12 <= \iac_raw_buf_vac_raw_buf_merged5_physical_RDATA_wire\(5);
    buf_data_vac_12 <= \iac_raw_buf_vac_raw_buf_merged5_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged5_physical_RADDR_wire\ <= '0'&\N__42967\&\N__24504\&\N__20346\&\N__43924\&\N__42220\&\N__38992\&\N__31435\&\N__36484\&\N__43165\&\N__31594\;
    \iac_raw_buf_vac_raw_buf_merged5_physical_WADDR_wire\ <= '0'&\N__40453\&\N__40561\&\N__39391\&\N__39496\&\N__39604\&\N__39712\&\N__39814\&\N__39922\&\N__40027\&\N__40132\;
    \iac_raw_buf_vac_raw_buf_merged5_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged5_physical_WDATA_wire\ <= '0'&'0'&\N__25812\&'0'&'0'&'0'&\N__21540\&'0'&'0'&'0'&\N__33461\&'0'&'0'&'0'&\N__24097\&'0';
    buf_data_iac_5 <= \iac_raw_buf_vac_raw_buf_merged9_physical_RDATA_wire\(13);
    buf_data_vac_5 <= \iac_raw_buf_vac_raw_buf_merged9_physical_RDATA_wire\(9);
    buf_data_iac_4 <= \iac_raw_buf_vac_raw_buf_merged9_physical_RDATA_wire\(5);
    buf_data_vac_4 <= \iac_raw_buf_vac_raw_buf_merged9_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged9_physical_RADDR_wire\ <= '0'&\N__42954\&\N__24501\&\N__20355\&\N__43911\&\N__42204\&\N__38979\&\N__31422\&\N__36465\&\N__43146\&\N__31575\;
    \iac_raw_buf_vac_raw_buf_merged9_physical_WADDR_wire\ <= '0'&\N__40434\&\N__40539\&\N__39378\&\N__39480\&\N__39585\&\N__39693\&\N__39801\&\N__39903\&\N__40008\&\N__40113\;
    \iac_raw_buf_vac_raw_buf_merged9_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged9_physical_WDATA_wire\ <= '0'&'0'&\N__49078\&'0'&'0'&'0'&\N__38308\&'0'&'0'&'0'&\N__48829\&'0'&'0'&'0'&\N__51331\&'0';
    buf_data_iac_15 <= \iac_raw_buf_vac_raw_buf_merged4_physical_RDATA_wire\(13);
    buf_data_vac_15 <= \iac_raw_buf_vac_raw_buf_merged4_physical_RDATA_wire\(9);
    buf_data_iac_14 <= \iac_raw_buf_vac_raw_buf_merged4_physical_RDATA_wire\(5);
    buf_data_vac_14 <= \iac_raw_buf_vac_raw_buf_merged4_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged4_physical_RADDR_wire\ <= '0'&\N__42973\&\N__24514\&\N__20358\&\N__43930\&\N__42226\&\N__38998\&\N__31441\&\N__36490\&\N__43171\&\N__31600\;
    \iac_raw_buf_vac_raw_buf_merged4_physical_WADDR_wire\ <= '0'&\N__40459\&\N__40567\&\N__39397\&\N__39502\&\N__39610\&\N__39718\&\N__39820\&\N__39928\&\N__40033\&\N__40138\;
    \iac_raw_buf_vac_raw_buf_merged4_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged4_physical_WDATA_wire\ <= '0'&'0'&\N__31990\&'0'&'0'&'0'&\N__20197\&'0'&'0'&'0'&\N__29586\&'0'&'0'&'0'&\N__22681\&'0';
    buf_data_iac_7 <= \iac_raw_buf_vac_raw_buf_merged8_physical_RDATA_wire\(13);
    buf_data_vac_7 <= \iac_raw_buf_vac_raw_buf_merged8_physical_RDATA_wire\(9);
    buf_data_iac_6 <= \iac_raw_buf_vac_raw_buf_merged8_physical_RDATA_wire\(5);
    buf_data_vac_6 <= \iac_raw_buf_vac_raw_buf_merged8_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged8_physical_RADDR_wire\ <= '0'&\N__42966\&\N__24513\&\N__20367\&\N__43923\&\N__42216\&\N__38991\&\N__31434\&\N__36477\&\N__43158\&\N__31587\;
    \iac_raw_buf_vac_raw_buf_merged8_physical_WADDR_wire\ <= '0'&\N__40446\&\N__40551\&\N__39390\&\N__39492\&\N__39597\&\N__39705\&\N__39813\&\N__39915\&\N__40020\&\N__40125\;
    \iac_raw_buf_vac_raw_buf_merged8_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged8_physical_WDATA_wire\ <= '0'&'0'&\N__47881\&'0'&'0'&'0'&\N__47932\&'0'&'0'&'0'&\N__48565\&'0'&'0'&'0'&\N__40864\&'0';
    buf_data_iac_3 <= \iac_raw_buf_vac_raw_buf_merged10_physical_RDATA_wire\(13);
    buf_data_vac_3 <= \iac_raw_buf_vac_raw_buf_merged10_physical_RDATA_wire\(9);
    buf_data_iac_2 <= \iac_raw_buf_vac_raw_buf_merged10_physical_RDATA_wire\(5);
    buf_data_vac_2 <= \iac_raw_buf_vac_raw_buf_merged10_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged10_physical_RADDR_wire\ <= '0'&\N__42997\&\N__24538\&\N__20386\&\N__43954\&\N__42250\&\N__39022\&\N__31465\&\N__36514\&\N__43195\&\N__31624\;
    \iac_raw_buf_vac_raw_buf_merged10_physical_WADDR_wire\ <= '0'&\N__40483\&\N__40591\&\N__39421\&\N__39526\&\N__39634\&\N__39742\&\N__39844\&\N__39952\&\N__40057\&\N__40162\;
    \iac_raw_buf_vac_raw_buf_merged10_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged10_physical_WDATA_wire\ <= '0'&'0'&\N__21046\&'0'&'0'&'0'&\N__21481\&'0'&'0'&'0'&\N__22495\&'0'&'0'&'0'&\N__22435\&'0';
    buf_data_iac_17 <= \iac_raw_buf_vac_raw_buf_merged3_physical_RDATA_wire\(13);
    buf_data_vac_17 <= \iac_raw_buf_vac_raw_buf_merged3_physical_RDATA_wire\(9);
    buf_data_iac_16 <= \iac_raw_buf_vac_raw_buf_merged3_physical_RDATA_wire\(5);
    buf_data_vac_16 <= \iac_raw_buf_vac_raw_buf_merged3_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged3_physical_RADDR_wire\ <= '0'&\N__42979\&\N__24520\&\N__20368\&\N__43936\&\N__42232\&\N__39004\&\N__31447\&\N__36496\&\N__43177\&\N__31606\;
    \iac_raw_buf_vac_raw_buf_merged3_physical_WADDR_wire\ <= '0'&\N__40465\&\N__40573\&\N__39403\&\N__39508\&\N__39616\&\N__39724\&\N__39826\&\N__39934\&\N__40039\&\N__40144\;
    \iac_raw_buf_vac_raw_buf_merged3_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged3_physical_WDATA_wire\ <= '0'&'0'&\N__26038\&'0'&'0'&'0'&\N__22657\&'0'&'0'&'0'&\N__27997\&'0'&'0'&'0'&\N__22595\&'0';
    buf_data_iac_1 <= \iac_raw_buf_vac_raw_buf_merged11_physical_RDATA_wire\(13);
    buf_data_vac_1 <= \iac_raw_buf_vac_raw_buf_merged11_physical_RDATA_wire\(9);
    buf_data_iac_0 <= \iac_raw_buf_vac_raw_buf_merged11_physical_RDATA_wire\(5);
    buf_data_vac_0 <= \iac_raw_buf_vac_raw_buf_merged11_physical_RDATA_wire\(1);
    \iac_raw_buf_vac_raw_buf_merged11_physical_RADDR_wire\ <= '0'&\N__42991\&\N__24532\&\N__20380\&\N__43948\&\N__42244\&\N__39016\&\N__31459\&\N__36508\&\N__43189\&\N__31618\;
    \iac_raw_buf_vac_raw_buf_merged11_physical_WADDR_wire\ <= '0'&\N__40477\&\N__40585\&\N__39415\&\N__39520\&\N__39628\&\N__39736\&\N__39838\&\N__39946\&\N__40051\&\N__40156\;
    \iac_raw_buf_vac_raw_buf_merged11_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \iac_raw_buf_vac_raw_buf_merged11_physical_WDATA_wire\ <= '0'&'0'&\N__23628\&'0'&'0'&'0'&\N__23968\&'0'&'0'&'0'&\N__23458\&'0'&'0'&'0'&\N__23482\&'0';

    \pll_main.zim_pll_inst\ : SB_PLL40_2F_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT_PORTB => "GENCLK_HALF",
            PLLOUT_SELECT_PORTA => "GENCLK",
            FILTER_RANGE => "011",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE_PORTB => '0',
            ENABLE_ICEGATE_PORTA => '0',
            DIVR => "0000",
            DIVQ => "101",
            DIVF => "0011111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => \GNDG0\,
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCOREB => OPEN,
            REFERENCECLK => \N__19018\,
            RESETB => \N__52877\,
            BYPASS => \GNDG0\,
            PLLOUTCOREA => OPEN,
            SDI => \GNDG0\,
            PLLOUTGLOBALB => \clk_16MHz\,
            DYNAMICDELAY => \pll_main.zim_pll_inst_DYNAMICDELAY_wire\,
            LATCHINPUTVALUE => \GNDG0\,
            PLLOUTGLOBALA => \clk_32MHz\,
            SCLK => \GNDG0\
        );

    \iac_raw_buf_vac_raw_buf_merged2_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged2_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged2_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged2_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged2_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged2_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__55158\,
            RE => \N__52860\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged2WCLKN_net\,
            WE => \N__31753\
        );

    \iac_raw_buf_vac_raw_buf_merged7_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged7_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged7_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged7_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged7_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged7_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__55245\,
            RE => \N__52888\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged7WCLKN_net\,
            WE => \N__31751\
        );

    \iac_raw_buf_vac_raw_buf_merged1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged1_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged1_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged1_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged1_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__55093\,
            RE => \N__52873\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged1WCLKN_net\,
            WE => \N__31776\
        );

    \iac_raw_buf_vac_raw_buf_merged6_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged6_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged6_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged6_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged6_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged6_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__55242\,
            RE => \N__52887\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged6WCLKN_net\,
            WE => \N__31719\
        );

    \iac_raw_buf_vac_raw_buf_merged0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged0_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged0_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged0_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged0_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__55079\,
            RE => \N__52886\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged0WCLKN_net\,
            WE => \N__31777\
        );

    \iac_raw_buf_vac_raw_buf_merged5_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged5_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged5_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged5_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged5_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged5_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__55235\,
            RE => \N__52879\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged5WCLKN_net\,
            WE => \N__31750\
        );

    \iac_raw_buf_vac_raw_buf_merged9_physical\ : SB_RAM40_4K
    generic map (
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged9_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged9_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged9_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged9_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged9_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__55225\,
            RE => \N__52836\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged9WCLKN_net\,
            WE => \N__31766\
        );

    \iac_raw_buf_vac_raw_buf_merged4_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged4_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged4_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged4_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged4_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged4_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__55214\,
            RE => \N__52878\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged4WCLKN_net\,
            WE => \N__31726\
        );

    \iac_raw_buf_vac_raw_buf_merged8_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged8_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged8_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged8_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged8_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged8_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__55202\,
            RE => \N__52835\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged8WCLKN_net\,
            WE => \N__31767\
        );

    \iac_raw_buf_vac_raw_buf_merged10_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged10_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged10_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged10_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged10_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged10_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__55110\,
            RE => \N__52837\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged10WCLKN_net\,
            WE => \N__31769\
        );

    \iac_raw_buf_vac_raw_buf_merged3_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged3_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged3_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged3_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged3_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged3_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__55188\,
            RE => \N__52861\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged3WCLKN_net\,
            WE => \N__31752\
        );

    \iac_raw_buf_vac_raw_buf_merged11_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 2,
            READ_MODE => 2,
            INIT_F => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
            INIT_0 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \iac_raw_buf_vac_raw_buf_merged11_physical_RDATA_wire\,
            RADDR => \iac_raw_buf_vac_raw_buf_merged11_physical_RADDR_wire\,
            WADDR => \iac_raw_buf_vac_raw_buf_merged11_physical_WADDR_wire\,
            MASK => \iac_raw_buf_vac_raw_buf_merged11_physical_MASK_wire\,
            WDATA => \iac_raw_buf_vac_raw_buf_merged11_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__55131\,
            RE => \N__52723\,
            WCLKE => 'H',
            WCLK => \INViac_raw_buf_vac_raw_buf_merged11WCLKN_net\,
            WE => \N__31768\
        );

    \ipInertedIOPad_VAC_DRDY_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58652\,
            DIN => \N__58651\,
            DOUT => \N__58650\,
            PACKAGEPIN => \VAC_DRDY_wire\
        );

    \ipInertedIOPad_VAC_DRDY_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58652\,
            PADOUT => \N__58651\,
            PADIN => \N__58650\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \VAC_DRDY\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_FLT1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58643\,
            DIN => \N__58642\,
            DOUT => \N__58641\,
            PACKAGEPIN => \IAC_FLT1_wire\
        );

    \ipInertedIOPad_IAC_FLT1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58643\,
            PADOUT => \N__58642\,
            PADIN => \N__58641\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__28099\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_SCK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58634\,
            DIN => \N__58633\,
            DOUT => \N__58632\,
            PACKAGEPIN => \DDS_SCK_wire\
        );

    \ipInertedIOPad_DDS_SCK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58634\,
            PADOUT => \N__58633\,
            PADIN => \N__58632\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__55915\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_166_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58625\,
            DIN => \N__58624\,
            DOUT => \N__58623\,
            PACKAGEPIN => \ICE_IOR_166_wire\
        );

    \ipInertedIOPad_ICE_IOR_166_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58625\,
            PADOUT => \N__58624\,
            PADIN => \N__58623\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_119_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58616\,
            DIN => \N__58615\,
            DOUT => \N__58614\,
            PACKAGEPIN => \ICE_IOR_119_wire\
        );

    \ipInertedIOPad_ICE_IOR_119_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58616\,
            PADOUT => \N__58615\,
            PADIN => \N__58614\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_MOSI_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58607\,
            DIN => \N__58606\,
            DOUT => \N__58605\,
            PACKAGEPIN => \DDS_MOSI_wire\
        );

    \ipInertedIOPad_DDS_MOSI_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58607\,
            PADOUT => \N__58606\,
            PADIN => \N__58605\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__42901\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_MISO_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58598\,
            DIN => \N__58597\,
            DOUT => \N__58596\,
            PACKAGEPIN => \VAC_MISO_wire\
        );

    \ipInertedIOPad_VAC_MISO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58598\,
            PADOUT => \N__58597\,
            PADIN => \N__58596\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \VAC_MISO\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_MOSI1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58589\,
            DIN => \N__58588\,
            DOUT => \N__58587\,
            PACKAGEPIN => \DDS_MOSI1_wire\
        );

    \ipInertedIOPad_DDS_MOSI1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58589\,
            PADOUT => \N__58588\,
            PADIN => \N__58587\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__21874\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_146_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58580\,
            DIN => \N__58579\,
            DOUT => \N__58578\,
            PACKAGEPIN => \ICE_IOR_146_wire\
        );

    \ipInertedIOPad_ICE_IOR_146_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58580\,
            PADOUT => \N__58579\,
            PADIN => \N__58578\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDC_CLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58571\,
            DIN => \N__58570\,
            DOUT => \N__58569\,
            PACKAGEPIN => \VDC_CLK_wire\
        );

    \ipInertedIOPad_VDC_CLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58571\,
            PADOUT => \N__58570\,
            PADIN => \N__58569\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__32914\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_222_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58562\,
            DIN => \N__58561\,
            DOUT => \N__58560\,
            PACKAGEPIN => \ICE_IOT_222_wire\
        );

    \ipInertedIOPad_ICE_IOT_222_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58562\,
            PADOUT => \N__58561\,
            PADIN => \N__58560\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_CS_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58553\,
            DIN => \N__58552\,
            DOUT => \N__58551\,
            PACKAGEPIN => \IAC_CS_wire\
        );

    \ipInertedIOPad_IAC_CS_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58553\,
            PADOUT => \N__58552\,
            PADIN => \N__58551\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__24847\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_18B_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58544\,
            DIN => \N__58543\,
            DOUT => \N__58542\,
            PACKAGEPIN => \ICE_IOL_18B_wire\
        );

    \ipInertedIOPad_ICE_IOL_18B_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58544\,
            PADOUT => \N__58543\,
            PADIN => \N__58542\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_13A_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58535\,
            DIN => \N__58534\,
            DOUT => \N__58533\,
            PACKAGEPIN => \ICE_IOL_13A_wire\
        );

    \ipInertedIOPad_ICE_IOL_13A_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58535\,
            PADOUT => \N__58534\,
            PADIN => \N__58533\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_81_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58526\,
            DIN => \N__58525\,
            DOUT => \N__58524\,
            PACKAGEPIN => \ICE_IOB_81_wire\
        );

    \ipInertedIOPad_ICE_IOB_81_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58526\,
            PADOUT => \N__58525\,
            PADIN => \N__58524\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_OSR1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58517\,
            DIN => \N__58516\,
            DOUT => \N__58515\,
            PACKAGEPIN => \VAC_OSR1_wire\
        );

    \ipInertedIOPad_VAC_OSR1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58517\,
            PADOUT => \N__58516\,
            PADIN => \N__58515\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__29725\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_MOSI_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58508\,
            DIN => \N__58507\,
            DOUT => \N__58506\,
            PACKAGEPIN => \IAC_MOSI_wire\
        );

    \ipInertedIOPad_IAC_MOSI_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58508\,
            PADOUT => \N__58507\,
            PADIN => \N__58506\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_CS1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58499\,
            DIN => \N__58498\,
            DOUT => \N__58497\,
            PACKAGEPIN => \DDS_CS1_wire\
        );

    \ipInertedIOPad_DDS_CS1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58499\,
            PADOUT => \N__58498\,
            PADIN => \N__58497\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__21631\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_4B_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58490\,
            DIN => \N__58489\,
            DOUT => \N__58488\,
            PACKAGEPIN => \ICE_IOL_4B_wire\
        );

    \ipInertedIOPad_ICE_IOL_4B_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58490\,
            PADOUT => \N__58489\,
            PADIN => \N__58488\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_94_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58481\,
            DIN => \N__58480\,
            DOUT => \N__58479\,
            PACKAGEPIN => \ICE_IOB_94_wire\
        );

    \ipInertedIOPad_ICE_IOB_94_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58481\,
            PADOUT => \N__58480\,
            PADIN => \N__58479\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_CS_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58472\,
            DIN => \N__58471\,
            DOUT => \N__58470\,
            PACKAGEPIN => \VAC_CS_wire\
        );

    \ipInertedIOPad_VAC_CS_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58472\,
            PADOUT => \N__58471\,
            PADIN => \N__58470\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__20254\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_CLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58463\,
            DIN => \N__58462\,
            DOUT => \N__58461\,
            PACKAGEPIN => \VAC_CLK_wire\
        );

    \ipInertedIOPad_VAC_CLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58463\,
            PADOUT => \N__58462\,
            PADIN => \N__58461\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__26148\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_SPI_CE0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58454\,
            DIN => \N__58453\,
            DOUT => \N__58452\,
            PACKAGEPIN => \ICE_SPI_CE0_wire\
        );

    \ipInertedIOPad_ICE_SPI_CE0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58454\,
            PADOUT => \N__58453\,
            PADIN => \N__58452\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \ICE_SPI_CE0\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_167_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58445\,
            DIN => \N__58444\,
            DOUT => \N__58443\,
            PACKAGEPIN => \ICE_IOR_167_wire\
        );

    \ipInertedIOPad_ICE_IOR_167_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58445\,
            PADOUT => \N__58444\,
            PADIN => \N__58443\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_118_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58436\,
            DIN => \N__58435\,
            DOUT => \N__58434\,
            PACKAGEPIN => \ICE_IOR_118_wire\
        );

    \ipInertedIOPad_ICE_IOR_118_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58436\,
            PADOUT => \N__58435\,
            PADIN => \N__58434\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_RTD_SDO_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58427\,
            DIN => \N__58426\,
            DOUT => \N__58425\,
            PACKAGEPIN => \RTD_SDO_wire\
        );

    \ipInertedIOPad_RTD_SDO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58427\,
            PADOUT => \N__58426\,
            PADIN => \N__58425\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \RTD_SDO\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_OSR0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58418\,
            DIN => \N__58417\,
            DOUT => \N__58416\,
            PACKAGEPIN => \IAC_OSR0_wire\
        );

    \ipInertedIOPad_IAC_OSR0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58418\,
            PADOUT => \N__58417\,
            PADIN => \N__58416\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__28225\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDC_SCLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58409\,
            DIN => \N__58408\,
            DOUT => \N__58407\,
            PACKAGEPIN => \VDC_SCLK_wire\
        );

    \ipInertedIOPad_VDC_SCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58409\,
            PADOUT => \N__58408\,
            PADIN => \N__58407\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__26938\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_FLT1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58400\,
            DIN => \N__58399\,
            DOUT => \N__58398\,
            PACKAGEPIN => \VAC_FLT1_wire\
        );

    \ipInertedIOPad_VAC_FLT1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58400\,
            PADOUT => \N__58399\,
            PADIN => \N__58398\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__26221\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_SPI_MOSI_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58391\,
            DIN => \N__58390\,
            DOUT => \N__58389\,
            PACKAGEPIN => \ICE_SPI_MOSI_wire\
        );

    \ipInertedIOPad_ICE_SPI_MOSI_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58391\,
            PADOUT => \N__58390\,
            PADIN => \N__58389\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \ICE_SPI_MOSI\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_165_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58382\,
            DIN => \N__58381\,
            DOUT => \N__58380\,
            PACKAGEPIN => \ICE_IOR_165_wire\
        );

    \ipInertedIOPad_ICE_IOR_165_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58382\,
            PADOUT => \N__58381\,
            PADIN => \N__58380\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_147_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58373\,
            DIN => \N__58372\,
            DOUT => \N__58371\,
            PACKAGEPIN => \ICE_IOR_147_wire\
        );

    \ipInertedIOPad_ICE_IOR_147_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58373\,
            PADOUT => \N__58372\,
            PADIN => \N__58371\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_14A_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58364\,
            DIN => \N__58363\,
            DOUT => \N__58362\,
            PACKAGEPIN => \ICE_IOL_14A_wire\
        );

    \ipInertedIOPad_ICE_IOL_14A_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58364\,
            PADOUT => \N__58363\,
            PADIN => \N__58362\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_13B_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58355\,
            DIN => \N__58354\,
            DOUT => \N__58353\,
            PACKAGEPIN => \ICE_IOL_13B_wire\
        );

    \ipInertedIOPad_ICE_IOL_13B_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58355\,
            PADOUT => \N__58354\,
            PADIN => \N__58353\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_91_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58346\,
            DIN => \N__58345\,
            DOUT => \N__58344\,
            PACKAGEPIN => \ICE_IOB_91_wire\
        );

    \ipInertedIOPad_ICE_IOB_91_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58346\,
            PADOUT => \N__58345\,
            PADIN => \N__58344\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_GPMO_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58337\,
            DIN => \N__58336\,
            DOUT => \N__58335\,
            PACKAGEPIN => \ICE_GPMO_0_wire\
        );

    \ipInertedIOPad_ICE_GPMO_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58337\,
            PADOUT => \N__58336\,
            PADIN => \N__58335\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_RNG_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58328\,
            DIN => \N__58327\,
            DOUT => \N__58326\,
            PACKAGEPIN => \DDS_RNG_0_wire\
        );

    \ipInertedIOPad_DDS_RNG_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58328\,
            PADOUT => \N__58327\,
            PADIN => \N__58326\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__44035\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDC_RNG0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58319\,
            DIN => \N__58318\,
            DOUT => \N__58317\,
            PACKAGEPIN => \VDC_RNG0_wire\
        );

    \ipInertedIOPad_VDC_RNG0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58319\,
            PADOUT => \N__58318\,
            PADIN => \N__58317\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__44767\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_SPI_SCLK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58310\,
            DIN => \N__58309\,
            DOUT => \N__58308\,
            PACKAGEPIN => \ICE_SPI_SCLK_wire\
        );

    \ipInertedIOPad_ICE_SPI_SCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58310\,
            PADOUT => \N__58309\,
            PADIN => \N__58308\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \ICE_SPI_SCLK\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_152_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58301\,
            DIN => \N__58300\,
            DOUT => \N__58299\,
            PACKAGEPIN => \ICE_IOR_152_wire\
        );

    \ipInertedIOPad_ICE_IOR_152_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58301\,
            PADOUT => \N__58300\,
            PADIN => \N__58299\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_12A_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58292\,
            DIN => \N__58291\,
            DOUT => \N__58290\,
            PACKAGEPIN => \ICE_IOL_12A_wire\
        );

    \ipInertedIOPad_ICE_IOL_12A_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58292\,
            PADOUT => \N__58291\,
            PADIN => \N__58290\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_RTD_DRDY_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58283\,
            DIN => \N__58282\,
            DOUT => \N__58281\,
            PACKAGEPIN => \RTD_DRDY_wire\
        );

    \ipInertedIOPad_RTD_DRDY_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58283\,
            PADOUT => \N__58282\,
            PADIN => \N__58281\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \RTD_DRDY\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_SPI_MISO_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58274\,
            DIN => \N__58273\,
            DOUT => \N__58272\,
            PACKAGEPIN => \ICE_SPI_MISO_wire\
        );

    \ipInertedIOPad_ICE_SPI_MISO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58274\,
            PADOUT => \N__58273\,
            PADIN => \N__58272\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__43591\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_177_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58265\,
            DIN => \N__58264\,
            DOUT => \N__58263\,
            PACKAGEPIN => \ICE_IOT_177_wire\
        );

    \ipInertedIOPad_ICE_IOT_177_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58265\,
            PADOUT => \N__58264\,
            PADIN => \N__58263\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_141_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58256\,
            DIN => \N__58255\,
            DOUT => \N__58254\,
            PACKAGEPIN => \ICE_IOR_141_wire\
        );

    \ipInertedIOPad_ICE_IOR_141_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58256\,
            PADOUT => \N__58255\,
            PADIN => \N__58254\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_80_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58247\,
            DIN => \N__58246\,
            DOUT => \N__58245\,
            PACKAGEPIN => \ICE_IOB_80_wire\
        );

    \ipInertedIOPad_ICE_IOB_80_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58247\,
            PADOUT => \N__58246\,
            PADIN => \N__58245\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_102_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58238\,
            DIN => \N__58237\,
            DOUT => \N__58236\,
            PACKAGEPIN => \ICE_IOB_102_wire\
        );

    \ipInertedIOPad_ICE_IOB_102_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58238\,
            PADOUT => \N__58237\,
            PADIN => \N__58236\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_GPMO_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58229\,
            DIN => \N__58228\,
            DOUT => \N__58227\,
            PACKAGEPIN => \ICE_GPMO_2_wire\
        );

    \ipInertedIOPad_ICE_GPMO_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58229\,
            PADOUT => \N__58228\,
            PADIN => \N__58227\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \ICE_GPMO_2\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_GPMI_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58220\,
            DIN => \N__58219\,
            DOUT => \N__58218\,
            PACKAGEPIN => \ICE_GPMI_0_wire\
        );

    \ipInertedIOPad_ICE_GPMI_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58220\,
            PADOUT => \N__58219\,
            PADIN => \N__58218\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__49267\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_MISO_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58211\,
            DIN => \N__58210\,
            DOUT => \N__58209\,
            PACKAGEPIN => \IAC_MISO_wire\
        );

    \ipInertedIOPad_IAC_MISO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58211\,
            PADOUT => \N__58210\,
            PADIN => \N__58209\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \IAC_MISO\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_OSR0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58202\,
            DIN => \N__58201\,
            DOUT => \N__58200\,
            PACKAGEPIN => \VAC_OSR0_wire\
        );

    \ipInertedIOPad_VAC_OSR0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58202\,
            PADOUT => \N__58201\,
            PADIN => \N__58200\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__26113\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_MOSI_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58193\,
            DIN => \N__58192\,
            DOUT => \N__58191\,
            PACKAGEPIN => \VAC_MOSI_wire\
        );

    \ipInertedIOPad_VAC_MOSI_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58193\,
            PADOUT => \N__58192\,
            PADIN => \N__58191\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_TEST_LED_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58184\,
            DIN => \N__58183\,
            DOUT => \N__58182\,
            PACKAGEPIN => \TEST_LED_wire\
        );

    \ipInertedIOPad_TEST_LED_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58184\,
            PADOUT => \N__58183\,
            PADIN => \N__58182\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__40945\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_148_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58175\,
            DIN => \N__58174\,
            DOUT => \N__58173\,
            PACKAGEPIN => \ICE_IOR_148_wire\
        );

    \ipInertedIOPad_ICE_IOR_148_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58175\,
            PADOUT => \N__58174\,
            PADIN => \N__58173\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_STAT_COMM_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58166\,
            DIN => \N__58165\,
            DOUT => \N__58164\,
            PACKAGEPIN => \STAT_COMM_wire\
        );

    \ipInertedIOPad_STAT_COMM_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58166\,
            PADOUT => \N__58165\,
            PADIN => \N__58164\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__19003\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_SYSCLK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58157\,
            DIN => \N__58156\,
            DOUT => \N__58155\,
            PACKAGEPIN => \ICE_SYSCLK_wire\
        );

    \ipInertedIOPad_ICE_SYSCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58157\,
            PADOUT => \N__58156\,
            PADIN => \N__58155\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \ICE_SYSCLK\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_161_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58148\,
            DIN => \N__58147\,
            DOUT => \N__58146\,
            PACKAGEPIN => \ICE_IOR_161_wire\
        );

    \ipInertedIOPad_ICE_IOR_161_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58148\,
            PADOUT => \N__58147\,
            PADIN => \N__58146\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_95_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58139\,
            DIN => \N__58138\,
            DOUT => \N__58137\,
            PACKAGEPIN => \ICE_IOB_95_wire\
        );

    \ipInertedIOPad_ICE_IOB_95_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58139\,
            PADOUT => \N__58138\,
            PADIN => \N__58137\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_82_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58130\,
            DIN => \N__58129\,
            DOUT => \N__58128\,
            PACKAGEPIN => \ICE_IOB_82_wire\
        );

    \ipInertedIOPad_ICE_IOB_82_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58130\,
            PADOUT => \N__58129\,
            PADIN => \N__58128\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_104_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58121\,
            DIN => \N__58120\,
            DOUT => \N__58119\,
            PACKAGEPIN => \ICE_IOB_104_wire\
        );

    \ipInertedIOPad_ICE_IOB_104_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58121\,
            PADOUT => \N__58120\,
            PADIN => \N__58119\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_CLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58112\,
            DIN => \N__58111\,
            DOUT => \N__58110\,
            PACKAGEPIN => \IAC_CLK_wire\
        );

    \ipInertedIOPad_IAC_CLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58112\,
            PADOUT => \N__58111\,
            PADIN => \N__58110\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__26152\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_CS_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58103\,
            DIN => \N__58102\,
            DOUT => \N__58101\,
            PACKAGEPIN => \DDS_CS_wire\
        );

    \ipInertedIOPad_DDS_CS_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58103\,
            PADOUT => \N__58102\,
            PADIN => \N__58101\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__55504\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SELIRNG0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58094\,
            DIN => \N__58093\,
            DOUT => \N__58092\,
            PACKAGEPIN => \SELIRNG0_wire\
        );

    \ipInertedIOPad_SELIRNG0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58094\,
            PADOUT => \N__58093\,
            PADIN => \N__58092\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__38185\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_RTD_SDI_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58085\,
            DIN => \N__58084\,
            DOUT => \N__58083\,
            PACKAGEPIN => \RTD_SDI_wire\
        );

    \ipInertedIOPad_RTD_SDI_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58085\,
            PADOUT => \N__58084\,
            PADIN => \N__58083\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__19798\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_221_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58076\,
            DIN => \N__58075\,
            DOUT => \N__58074\,
            PACKAGEPIN => \ICE_IOT_221_wire\
        );

    \ipInertedIOPad_ICE_IOT_221_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58076\,
            PADOUT => \N__58075\,
            PADIN => \N__58074\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_197_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58067\,
            DIN => \N__58066\,
            DOUT => \N__58065\,
            PACKAGEPIN => \ICE_IOT_197_wire\
        );

    \ipInertedIOPad_ICE_IOT_197_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58067\,
            PADOUT => \N__58066\,
            PADIN => \N__58065\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_MCLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58058\,
            DIN => \N__58057\,
            DOUT => \N__58056\,
            PACKAGEPIN => \DDS_MCLK_wire\
        );

    \ipInertedIOPad_DDS_MCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58058\,
            PADOUT => \N__58057\,
            PADIN => \N__58056\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__55933\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_RTD_SCLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58049\,
            DIN => \N__58048\,
            DOUT => \N__58047\,
            PACKAGEPIN => \RTD_SCLK_wire\
        );

    \ipInertedIOPad_RTD_SCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58049\,
            PADOUT => \N__58048\,
            PADIN => \N__58047\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__19045\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_RTD_CS_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58040\,
            DIN => \N__58039\,
            DOUT => \N__58038\,
            PACKAGEPIN => \RTD_CS_wire\
        );

    \ipInertedIOPad_RTD_CS_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58040\,
            PADOUT => \N__58039\,
            PADIN => \N__58038\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__19099\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_137_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58031\,
            DIN => \N__58030\,
            DOUT => \N__58029\,
            PACKAGEPIN => \ICE_IOR_137_wire\
        );

    \ipInertedIOPad_ICE_IOR_137_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58031\,
            PADOUT => \N__58030\,
            PADIN => \N__58029\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_OSR1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58022\,
            DIN => \N__58021\,
            DOUT => \N__58020\,
            PACKAGEPIN => \IAC_OSR1_wire\
        );

    \ipInertedIOPad_IAC_OSR1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58022\,
            PADOUT => \N__58021\,
            PADIN => \N__58020\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__28060\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_FLT0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__58013\,
            DIN => \N__58012\,
            DOUT => \N__58011\,
            PACKAGEPIN => \VAC_FLT0_wire\
        );

    \ipInertedIOPad_VAC_FLT0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58013\,
            PADOUT => \N__58012\,
            PADIN => \N__58011\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__27880\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_144_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__58004\,
            DIN => \N__58003\,
            DOUT => \N__58002\,
            PACKAGEPIN => \ICE_IOR_144_wire\
        );

    \ipInertedIOPad_ICE_IOR_144_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__58004\,
            PADOUT => \N__58003\,
            PADIN => \N__58002\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_128_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__57995\,
            DIN => \N__57994\,
            DOUT => \N__57993\,
            PACKAGEPIN => \ICE_IOR_128_wire\
        );

    \ipInertedIOPad_ICE_IOR_128_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__57995\,
            PADOUT => \N__57994\,
            PADIN => \N__57993\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_GPMO_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__57986\,
            DIN => \N__57985\,
            DOUT => \N__57984\,
            PACKAGEPIN => \ICE_GPMO_1_wire\
        );

    \ipInertedIOPad_ICE_GPMO_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__57986\,
            PADOUT => \N__57985\,
            PADIN => \N__57984\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_SCLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__57977\,
            DIN => \N__57976\,
            DOUT => \N__57975\,
            PACKAGEPIN => \IAC_SCLK_wire\
        );

    \ipInertedIOPad_IAC_SCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__57977\,
            PADOUT => \N__57976\,
            PADIN => \N__57975\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__26194\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_EIS_SYNCCLK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__57968\,
            DIN => \N__57967\,
            DOUT => \N__57966\,
            PACKAGEPIN => \EIS_SYNCCLK_wire\
        );

    \ipInertedIOPad_EIS_SYNCCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__57968\,
            PADOUT => \N__57967\,
            PADIN => \N__57966\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \EIS_SYNCCLK\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_139_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__57959\,
            DIN => \N__57958\,
            DOUT => \N__57957\,
            PACKAGEPIN => \ICE_IOR_139_wire\
        );

    \ipInertedIOPad_ICE_IOR_139_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__57959\,
            PADOUT => \N__57958\,
            PADIN => \N__57957\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_4A_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__57950\,
            DIN => \N__57949\,
            DOUT => \N__57948\,
            PACKAGEPIN => \ICE_IOL_4A_wire\
        );

    \ipInertedIOPad_ICE_IOL_4A_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__57950\,
            PADOUT => \N__57949\,
            PADIN => \N__57948\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VAC_SCLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__57941\,
            DIN => \N__57940\,
            DOUT => \N__57939\,
            PACKAGEPIN => \VAC_SCLK_wire\
        );

    \ipInertedIOPad_VAC_SCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__57941\,
            PADOUT => \N__57940\,
            PADIN => \N__57939\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__20227\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_THERMOSTAT_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__57932\,
            DIN => \N__57931\,
            DOUT => \N__57930\,
            PACKAGEPIN => \THERMOSTAT_wire\
        );

    \ipInertedIOPad_THERMOSTAT_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__57932\,
            PADOUT => \N__57931\,
            PADIN => \N__57930\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \THERMOSTAT\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_164_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__57923\,
            DIN => \N__57922\,
            DOUT => \N__57921\,
            PACKAGEPIN => \ICE_IOR_164_wire\
        );

    \ipInertedIOPad_ICE_IOR_164_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__57923\,
            PADOUT => \N__57922\,
            PADIN => \N__57921\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_103_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__57914\,
            DIN => \N__57913\,
            DOUT => \N__57912\,
            PACKAGEPIN => \ICE_IOB_103_wire\
        );

    \ipInertedIOPad_ICE_IOB_103_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__57914\,
            PADOUT => \N__57913\,
            PADIN => \N__57912\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_AMPV_POW_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__57905\,
            DIN => \N__57904\,
            DOUT => \N__57903\,
            PACKAGEPIN => \AMPV_POW_wire\
        );

    \ipInertedIOPad_AMPV_POW_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__57905\,
            PADOUT => \N__57904\,
            PADIN => \N__57903\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__30058\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDC_SDO_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__57896\,
            DIN => \N__57895\,
            DOUT => \N__57894\,
            PACKAGEPIN => \VDC_SDO_wire\
        );

    \ipInertedIOPad_VDC_SDO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__57896\,
            PADOUT => \N__57895\,
            PADIN => \N__57894\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \VDC_SDO\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_174_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__57887\,
            DIN => \N__57886\,
            DOUT => \N__57885\,
            PACKAGEPIN => \ICE_IOT_174_wire\
        );

    \ipInertedIOPad_ICE_IOT_174_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__57887\,
            PADOUT => \N__57886\,
            PADIN => \N__57885\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_140_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__57878\,
            DIN => \N__57877\,
            DOUT => \N__57876\,
            PACKAGEPIN => \ICE_IOR_140_wire\
        );

    \ipInertedIOPad_ICE_IOR_140_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__57878\,
            PADOUT => \N__57877\,
            PADIN => \N__57876\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOB_96_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__57869\,
            DIN => \N__57868\,
            DOUT => \N__57867\,
            PACKAGEPIN => \ICE_IOB_96_wire\
        );

    \ipInertedIOPad_ICE_IOB_96_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__57869\,
            PADOUT => \N__57868\,
            PADIN => \N__57867\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_CONT_SD_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__57860\,
            DIN => \N__57859\,
            DOUT => \N__57858\,
            PACKAGEPIN => \CONT_SD_wire\
        );

    \ipInertedIOPad_CONT_SD_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__57860\,
            PADOUT => \N__57859\,
            PADIN => \N__57858\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__50239\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_AC_ADC_SYNC_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__57851\,
            DIN => \N__57850\,
            DOUT => \N__57849\,
            PACKAGEPIN => \AC_ADC_SYNC_wire\
        );

    \ipInertedIOPad_AC_ADC_SYNC_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__57851\,
            PADOUT => \N__57850\,
            PADIN => \N__57849\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__26242\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SELIRNG1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__57842\,
            DIN => \N__57841\,
            DOUT => \N__57840\,
            PACKAGEPIN => \SELIRNG1_wire\
        );

    \ipInertedIOPad_SELIRNG1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__57842\,
            PADOUT => \N__57841\,
            PADIN => \N__57840\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__45511\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOL_12B_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__57833\,
            DIN => \N__57832\,
            DOUT => \N__57831\,
            PACKAGEPIN => \ICE_IOL_12B_wire\
        );

    \ipInertedIOPad_ICE_IOL_12B_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__57833\,
            PADOUT => \N__57832\,
            PADIN => \N__57831\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_160_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__57824\,
            DIN => \N__57823\,
            DOUT => \N__57822\,
            PACKAGEPIN => \ICE_IOR_160_wire\
        );

    \ipInertedIOPad_ICE_IOR_160_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__57824\,
            PADOUT => \N__57823\,
            PADIN => \N__57822\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_136_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__57815\,
            DIN => \N__57814\,
            DOUT => \N__57813\,
            PACKAGEPIN => \ICE_IOR_136_wire\
        );

    \ipInertedIOPad_ICE_IOR_136_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__57815\,
            PADOUT => \N__57814\,
            PADIN => \N__57813\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_MCLK1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__57806\,
            DIN => \N__57805\,
            DOUT => \N__57804\,
            PACKAGEPIN => \DDS_MCLK1_wire\
        );

    \ipInertedIOPad_DDS_MCLK1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__57806\,
            PADOUT => \N__57805\,
            PADIN => \N__57804\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__21649\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_198_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__57797\,
            DIN => \N__57796\,
            DOUT => \N__57795\,
            PACKAGEPIN => \ICE_IOT_198_wire\
        );

    \ipInertedIOPad_ICE_IOT_198_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__57797\,
            PADOUT => \N__57796\,
            PADIN => \N__57795\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_173_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__57788\,
            DIN => \N__57787\,
            DOUT => \N__57786\,
            PACKAGEPIN => \ICE_IOT_173_wire\
        );

    \ipInertedIOPad_ICE_IOT_173_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__57788\,
            PADOUT => \N__57787\,
            PADIN => \N__57786\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_DRDY_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__57779\,
            DIN => \N__57778\,
            DOUT => \N__57777\,
            PACKAGEPIN => \IAC_DRDY_wire\
        );

    \ipInertedIOPad_IAC_DRDY_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__57779\,
            PADOUT => \N__57778\,
            PADIN => \N__57777\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \IAC_DRDY\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOT_178_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__57770\,
            DIN => \N__57769\,
            DOUT => \N__57768\,
            PACKAGEPIN => \ICE_IOT_178_wire\
        );

    \ipInertedIOPad_ICE_IOT_178_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__57770\,
            PADOUT => \N__57769\,
            PADIN => \N__57768\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_138_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__57761\,
            DIN => \N__57760\,
            DOUT => \N__57759\,
            PACKAGEPIN => \ICE_IOR_138_wire\
        );

    \ipInertedIOPad_ICE_IOR_138_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__57761\,
            PADOUT => \N__57760\,
            PADIN => \N__57759\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICE_IOR_120_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__57752\,
            DIN => \N__57751\,
            DOUT => \N__57750\,
            PACKAGEPIN => \ICE_IOR_120_wire\
        );

    \ipInertedIOPad_ICE_IOR_120_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__57752\,
            PADOUT => \N__57751\,
            PADIN => \N__57750\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_IAC_FLT0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__57743\,
            DIN => \N__57742\,
            DOUT => \N__57741\,
            PACKAGEPIN => \IAC_FLT0_wire\
        );

    \ipInertedIOPad_IAC_FLT0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__57743\,
            PADOUT => \N__57742\,
            PADIN => \N__57741\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__28027\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DDS_SCK1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__57734\,
            DIN => \N__57733\,
            DOUT => \N__57732\,
            PACKAGEPIN => \DDS_SCK1_wire\
        );

    \ipInertedIOPad_DDS_SCK1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__57734\,
            PADOUT => \N__57733\,
            PADIN => \N__57732\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__21613\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \I__14461\ : InMux
    port map (
            O => \N__57715\,
            I => \N__57711\
        );

    \I__14460\ : InMux
    port map (
            O => \N__57714\,
            I => \N__57708\
        );

    \I__14459\ : LocalMux
    port map (
            O => \N__57711\,
            I => \N__57705\
        );

    \I__14458\ : LocalMux
    port map (
            O => \N__57708\,
            I => dds0_mclkcnt_0
        );

    \I__14457\ : Odrv4
    port map (
            O => \N__57705\,
            I => dds0_mclkcnt_0
        );

    \I__14456\ : InMux
    port map (
            O => \N__57700\,
            I => \bfn_22_11_0_\
        );

    \I__14455\ : CascadeMux
    port map (
            O => \N__57697\,
            I => \N__57694\
        );

    \I__14454\ : InMux
    port map (
            O => \N__57694\,
            I => \N__57690\
        );

    \I__14453\ : InMux
    port map (
            O => \N__57693\,
            I => \N__57687\
        );

    \I__14452\ : LocalMux
    port map (
            O => \N__57690\,
            I => \N__57684\
        );

    \I__14451\ : LocalMux
    port map (
            O => \N__57687\,
            I => \N__57679\
        );

    \I__14450\ : Span4Mux_h
    port map (
            O => \N__57684\,
            I => \N__57679\
        );

    \I__14449\ : Odrv4
    port map (
            O => \N__57679\,
            I => dds0_mclkcnt_1
        );

    \I__14448\ : InMux
    port map (
            O => \N__57676\,
            I => n19440
        );

    \I__14447\ : CascadeMux
    port map (
            O => \N__57673\,
            I => \N__57670\
        );

    \I__14446\ : InMux
    port map (
            O => \N__57670\,
            I => \N__57666\
        );

    \I__14445\ : InMux
    port map (
            O => \N__57669\,
            I => \N__57663\
        );

    \I__14444\ : LocalMux
    port map (
            O => \N__57666\,
            I => \N__57660\
        );

    \I__14443\ : LocalMux
    port map (
            O => \N__57663\,
            I => dds0_mclkcnt_2
        );

    \I__14442\ : Odrv4
    port map (
            O => \N__57660\,
            I => dds0_mclkcnt_2
        );

    \I__14441\ : InMux
    port map (
            O => \N__57655\,
            I => n19441
        );

    \I__14440\ : InMux
    port map (
            O => \N__57652\,
            I => \N__57648\
        );

    \I__14439\ : InMux
    port map (
            O => \N__57651\,
            I => \N__57645\
        );

    \I__14438\ : LocalMux
    port map (
            O => \N__57648\,
            I => \N__57642\
        );

    \I__14437\ : LocalMux
    port map (
            O => \N__57645\,
            I => dds0_mclkcnt_3
        );

    \I__14436\ : Odrv12
    port map (
            O => \N__57642\,
            I => dds0_mclkcnt_3
        );

    \I__14435\ : InMux
    port map (
            O => \N__57637\,
            I => n19442
        );

    \I__14434\ : InMux
    port map (
            O => \N__57634\,
            I => \N__57630\
        );

    \I__14433\ : InMux
    port map (
            O => \N__57633\,
            I => \N__57627\
        );

    \I__14432\ : LocalMux
    port map (
            O => \N__57630\,
            I => \N__57624\
        );

    \I__14431\ : LocalMux
    port map (
            O => \N__57627\,
            I => dds0_mclkcnt_4
        );

    \I__14430\ : Odrv4
    port map (
            O => \N__57624\,
            I => dds0_mclkcnt_4
        );

    \I__14429\ : InMux
    port map (
            O => \N__57619\,
            I => n19443
        );

    \I__14428\ : InMux
    port map (
            O => \N__57616\,
            I => \N__57612\
        );

    \I__14427\ : InMux
    port map (
            O => \N__57615\,
            I => \N__57609\
        );

    \I__14426\ : LocalMux
    port map (
            O => \N__57612\,
            I => \N__57606\
        );

    \I__14425\ : LocalMux
    port map (
            O => \N__57609\,
            I => dds0_mclkcnt_5
        );

    \I__14424\ : Odrv4
    port map (
            O => \N__57606\,
            I => dds0_mclkcnt_5
        );

    \I__14423\ : InMux
    port map (
            O => \N__57601\,
            I => n19444
        );

    \I__14422\ : InMux
    port map (
            O => \N__57598\,
            I => \N__57595\
        );

    \I__14421\ : LocalMux
    port map (
            O => \N__57595\,
            I => \N__57592\
        );

    \I__14420\ : Odrv4
    port map (
            O => \N__57592\,
            I => n10
        );

    \I__14419\ : InMux
    port map (
            O => \N__57589\,
            I => \N__57583\
        );

    \I__14418\ : InMux
    port map (
            O => \N__57588\,
            I => \N__57583\
        );

    \I__14417\ : LocalMux
    port map (
            O => \N__57583\,
            I => \N__57580\
        );

    \I__14416\ : Span4Mux_h
    port map (
            O => \N__57580\,
            I => \N__57577\
        );

    \I__14415\ : Odrv4
    port map (
            O => \N__57577\,
            I => dds0_mclkcnt_6
        );

    \I__14414\ : InMux
    port map (
            O => \N__57574\,
            I => n19445
        );

    \I__14413\ : InMux
    port map (
            O => \N__57571\,
            I => n19446
        );

    \I__14412\ : InMux
    port map (
            O => \N__57568\,
            I => \N__57564\
        );

    \I__14411\ : InMux
    port map (
            O => \N__57567\,
            I => \N__57561\
        );

    \I__14410\ : LocalMux
    port map (
            O => \N__57564\,
            I => \N__57558\
        );

    \I__14409\ : LocalMux
    port map (
            O => \N__57561\,
            I => dds0_mclkcnt_7
        );

    \I__14408\ : Odrv4
    port map (
            O => \N__57558\,
            I => dds0_mclkcnt_7
        );

    \I__14407\ : InMux
    port map (
            O => \N__57553\,
            I => \N__57544\
        );

    \I__14406\ : InMux
    port map (
            O => \N__57552\,
            I => \N__57526\
        );

    \I__14405\ : InMux
    port map (
            O => \N__57551\,
            I => \N__57526\
        );

    \I__14404\ : InMux
    port map (
            O => \N__57550\,
            I => \N__57516\
        );

    \I__14403\ : InMux
    port map (
            O => \N__57549\,
            I => \N__57516\
        );

    \I__14402\ : InMux
    port map (
            O => \N__57548\,
            I => \N__57513\
        );

    \I__14401\ : InMux
    port map (
            O => \N__57547\,
            I => \N__57510\
        );

    \I__14400\ : LocalMux
    port map (
            O => \N__57544\,
            I => \N__57507\
        );

    \I__14399\ : InMux
    port map (
            O => \N__57543\,
            I => \N__57504\
        );

    \I__14398\ : InMux
    port map (
            O => \N__57542\,
            I => \N__57497\
        );

    \I__14397\ : InMux
    port map (
            O => \N__57541\,
            I => \N__57497\
        );

    \I__14396\ : InMux
    port map (
            O => \N__57540\,
            I => \N__57494\
        );

    \I__14395\ : InMux
    port map (
            O => \N__57539\,
            I => \N__57490\
        );

    \I__14394\ : CascadeMux
    port map (
            O => \N__57538\,
            I => \N__57486\
        );

    \I__14393\ : InMux
    port map (
            O => \N__57537\,
            I => \N__57472\
        );

    \I__14392\ : InMux
    port map (
            O => \N__57536\,
            I => \N__57472\
        );

    \I__14391\ : InMux
    port map (
            O => \N__57535\,
            I => \N__57472\
        );

    \I__14390\ : InMux
    port map (
            O => \N__57534\,
            I => \N__57469\
        );

    \I__14389\ : CascadeMux
    port map (
            O => \N__57533\,
            I => \N__57466\
        );

    \I__14388\ : InMux
    port map (
            O => \N__57532\,
            I => \N__57459\
        );

    \I__14387\ : InMux
    port map (
            O => \N__57531\,
            I => \N__57456\
        );

    \I__14386\ : LocalMux
    port map (
            O => \N__57526\,
            I => \N__57453\
        );

    \I__14385\ : InMux
    port map (
            O => \N__57525\,
            I => \N__57450\
        );

    \I__14384\ : CascadeMux
    port map (
            O => \N__57524\,
            I => \N__57437\
        );

    \I__14383\ : InMux
    port map (
            O => \N__57523\,
            I => \N__57433\
        );

    \I__14382\ : InMux
    port map (
            O => \N__57522\,
            I => \N__57430\
        );

    \I__14381\ : InMux
    port map (
            O => \N__57521\,
            I => \N__57427\
        );

    \I__14380\ : LocalMux
    port map (
            O => \N__57516\,
            I => \N__57422\
        );

    \I__14379\ : LocalMux
    port map (
            O => \N__57513\,
            I => \N__57422\
        );

    \I__14378\ : LocalMux
    port map (
            O => \N__57510\,
            I => \N__57419\
        );

    \I__14377\ : Span4Mux_h
    port map (
            O => \N__57507\,
            I => \N__57414\
        );

    \I__14376\ : LocalMux
    port map (
            O => \N__57504\,
            I => \N__57414\
        );

    \I__14375\ : InMux
    port map (
            O => \N__57503\,
            I => \N__57411\
        );

    \I__14374\ : InMux
    port map (
            O => \N__57502\,
            I => \N__57404\
        );

    \I__14373\ : LocalMux
    port map (
            O => \N__57497\,
            I => \N__57399\
        );

    \I__14372\ : LocalMux
    port map (
            O => \N__57494\,
            I => \N__57399\
        );

    \I__14371\ : InMux
    port map (
            O => \N__57493\,
            I => \N__57396\
        );

    \I__14370\ : LocalMux
    port map (
            O => \N__57490\,
            I => \N__57383\
        );

    \I__14369\ : InMux
    port map (
            O => \N__57489\,
            I => \N__57380\
        );

    \I__14368\ : InMux
    port map (
            O => \N__57486\,
            I => \N__57377\
        );

    \I__14367\ : InMux
    port map (
            O => \N__57485\,
            I => \N__57374\
        );

    \I__14366\ : InMux
    port map (
            O => \N__57484\,
            I => \N__57371\
        );

    \I__14365\ : InMux
    port map (
            O => \N__57483\,
            I => \N__57367\
        );

    \I__14364\ : InMux
    port map (
            O => \N__57482\,
            I => \N__57364\
        );

    \I__14363\ : InMux
    port map (
            O => \N__57481\,
            I => \N__57359\
        );

    \I__14362\ : InMux
    port map (
            O => \N__57480\,
            I => \N__57359\
        );

    \I__14361\ : InMux
    port map (
            O => \N__57479\,
            I => \N__57356\
        );

    \I__14360\ : LocalMux
    port map (
            O => \N__57472\,
            I => \N__57353\
        );

    \I__14359\ : LocalMux
    port map (
            O => \N__57469\,
            I => \N__57350\
        );

    \I__14358\ : InMux
    port map (
            O => \N__57466\,
            I => \N__57347\
        );

    \I__14357\ : CascadeMux
    port map (
            O => \N__57465\,
            I => \N__57342\
        );

    \I__14356\ : InMux
    port map (
            O => \N__57464\,
            I => \N__57334\
        );

    \I__14355\ : InMux
    port map (
            O => \N__57463\,
            I => \N__57334\
        );

    \I__14354\ : InMux
    port map (
            O => \N__57462\,
            I => \N__57334\
        );

    \I__14353\ : LocalMux
    port map (
            O => \N__57459\,
            I => \N__57331\
        );

    \I__14352\ : LocalMux
    port map (
            O => \N__57456\,
            I => \N__57328\
        );

    \I__14351\ : Span4Mux_v
    port map (
            O => \N__57453\,
            I => \N__57323\
        );

    \I__14350\ : LocalMux
    port map (
            O => \N__57450\,
            I => \N__57323\
        );

    \I__14349\ : InMux
    port map (
            O => \N__57449\,
            I => \N__57318\
        );

    \I__14348\ : InMux
    port map (
            O => \N__57448\,
            I => \N__57318\
        );

    \I__14347\ : CascadeMux
    port map (
            O => \N__57447\,
            I => \N__57315\
        );

    \I__14346\ : InMux
    port map (
            O => \N__57446\,
            I => \N__57312\
        );

    \I__14345\ : InMux
    port map (
            O => \N__57445\,
            I => \N__57305\
        );

    \I__14344\ : InMux
    port map (
            O => \N__57444\,
            I => \N__57305\
        );

    \I__14343\ : InMux
    port map (
            O => \N__57443\,
            I => \N__57300\
        );

    \I__14342\ : InMux
    port map (
            O => \N__57442\,
            I => \N__57300\
        );

    \I__14341\ : InMux
    port map (
            O => \N__57441\,
            I => \N__57297\
        );

    \I__14340\ : InMux
    port map (
            O => \N__57440\,
            I => \N__57294\
        );

    \I__14339\ : InMux
    port map (
            O => \N__57437\,
            I => \N__57291\
        );

    \I__14338\ : InMux
    port map (
            O => \N__57436\,
            I => \N__57288\
        );

    \I__14337\ : LocalMux
    port map (
            O => \N__57433\,
            I => \N__57279\
        );

    \I__14336\ : LocalMux
    port map (
            O => \N__57430\,
            I => \N__57279\
        );

    \I__14335\ : LocalMux
    port map (
            O => \N__57427\,
            I => \N__57279\
        );

    \I__14334\ : Span4Mux_h
    port map (
            O => \N__57422\,
            I => \N__57279\
        );

    \I__14333\ : Span4Mux_v
    port map (
            O => \N__57419\,
            I => \N__57274\
        );

    \I__14332\ : Span4Mux_h
    port map (
            O => \N__57414\,
            I => \N__57274\
        );

    \I__14331\ : LocalMux
    port map (
            O => \N__57411\,
            I => \N__57271\
        );

    \I__14330\ : InMux
    port map (
            O => \N__57410\,
            I => \N__57262\
        );

    \I__14329\ : InMux
    port map (
            O => \N__57409\,
            I => \N__57262\
        );

    \I__14328\ : InMux
    port map (
            O => \N__57408\,
            I => \N__57262\
        );

    \I__14327\ : InMux
    port map (
            O => \N__57407\,
            I => \N__57262\
        );

    \I__14326\ : LocalMux
    port map (
            O => \N__57404\,
            I => \N__57259\
        );

    \I__14325\ : Span4Mux_v
    port map (
            O => \N__57399\,
            I => \N__57254\
        );

    \I__14324\ : LocalMux
    port map (
            O => \N__57396\,
            I => \N__57254\
        );

    \I__14323\ : InMux
    port map (
            O => \N__57395\,
            I => \N__57251\
        );

    \I__14322\ : InMux
    port map (
            O => \N__57394\,
            I => \N__57243\
        );

    \I__14321\ : InMux
    port map (
            O => \N__57393\,
            I => \N__57243\
        );

    \I__14320\ : InMux
    port map (
            O => \N__57392\,
            I => \N__57243\
        );

    \I__14319\ : InMux
    port map (
            O => \N__57391\,
            I => \N__57238\
        );

    \I__14318\ : InMux
    port map (
            O => \N__57390\,
            I => \N__57233\
        );

    \I__14317\ : InMux
    port map (
            O => \N__57389\,
            I => \N__57233\
        );

    \I__14316\ : InMux
    port map (
            O => \N__57388\,
            I => \N__57230\
        );

    \I__14315\ : InMux
    port map (
            O => \N__57387\,
            I => \N__57225\
        );

    \I__14314\ : InMux
    port map (
            O => \N__57386\,
            I => \N__57225\
        );

    \I__14313\ : Span4Mux_h
    port map (
            O => \N__57383\,
            I => \N__57220\
        );

    \I__14312\ : LocalMux
    port map (
            O => \N__57380\,
            I => \N__57220\
        );

    \I__14311\ : LocalMux
    port map (
            O => \N__57377\,
            I => \N__57215\
        );

    \I__14310\ : LocalMux
    port map (
            O => \N__57374\,
            I => \N__57215\
        );

    \I__14309\ : LocalMux
    port map (
            O => \N__57371\,
            I => \N__57212\
        );

    \I__14308\ : InMux
    port map (
            O => \N__57370\,
            I => \N__57209\
        );

    \I__14307\ : LocalMux
    port map (
            O => \N__57367\,
            I => \N__57206\
        );

    \I__14306\ : LocalMux
    port map (
            O => \N__57364\,
            I => \N__57193\
        );

    \I__14305\ : LocalMux
    port map (
            O => \N__57359\,
            I => \N__57193\
        );

    \I__14304\ : LocalMux
    port map (
            O => \N__57356\,
            I => \N__57193\
        );

    \I__14303\ : Span4Mux_h
    port map (
            O => \N__57353\,
            I => \N__57193\
        );

    \I__14302\ : Span4Mux_v
    port map (
            O => \N__57350\,
            I => \N__57193\
        );

    \I__14301\ : LocalMux
    port map (
            O => \N__57347\,
            I => \N__57193\
        );

    \I__14300\ : InMux
    port map (
            O => \N__57346\,
            I => \N__57172\
        );

    \I__14299\ : InMux
    port map (
            O => \N__57345\,
            I => \N__57172\
        );

    \I__14298\ : InMux
    port map (
            O => \N__57342\,
            I => \N__57172\
        );

    \I__14297\ : InMux
    port map (
            O => \N__57341\,
            I => \N__57172\
        );

    \I__14296\ : LocalMux
    port map (
            O => \N__57334\,
            I => \N__57163\
        );

    \I__14295\ : Span4Mux_h
    port map (
            O => \N__57331\,
            I => \N__57163\
        );

    \I__14294\ : Span4Mux_v
    port map (
            O => \N__57328\,
            I => \N__57163\
        );

    \I__14293\ : Span4Mux_h
    port map (
            O => \N__57323\,
            I => \N__57163\
        );

    \I__14292\ : LocalMux
    port map (
            O => \N__57318\,
            I => \N__57160\
        );

    \I__14291\ : InMux
    port map (
            O => \N__57315\,
            I => \N__57157\
        );

    \I__14290\ : LocalMux
    port map (
            O => \N__57312\,
            I => \N__57154\
        );

    \I__14289\ : InMux
    port map (
            O => \N__57311\,
            I => \N__57149\
        );

    \I__14288\ : InMux
    port map (
            O => \N__57310\,
            I => \N__57149\
        );

    \I__14287\ : LocalMux
    port map (
            O => \N__57305\,
            I => \N__57142\
        );

    \I__14286\ : LocalMux
    port map (
            O => \N__57300\,
            I => \N__57142\
        );

    \I__14285\ : LocalMux
    port map (
            O => \N__57297\,
            I => \N__57142\
        );

    \I__14284\ : LocalMux
    port map (
            O => \N__57294\,
            I => \N__57135\
        );

    \I__14283\ : LocalMux
    port map (
            O => \N__57291\,
            I => \N__57135\
        );

    \I__14282\ : LocalMux
    port map (
            O => \N__57288\,
            I => \N__57135\
        );

    \I__14281\ : Span4Mux_v
    port map (
            O => \N__57279\,
            I => \N__57126\
        );

    \I__14280\ : Span4Mux_h
    port map (
            O => \N__57274\,
            I => \N__57126\
        );

    \I__14279\ : Span4Mux_h
    port map (
            O => \N__57271\,
            I => \N__57126\
        );

    \I__14278\ : LocalMux
    port map (
            O => \N__57262\,
            I => \N__57126\
        );

    \I__14277\ : Sp12to4
    port map (
            O => \N__57259\,
            I => \N__57119\
        );

    \I__14276\ : Sp12to4
    port map (
            O => \N__57254\,
            I => \N__57119\
        );

    \I__14275\ : LocalMux
    port map (
            O => \N__57251\,
            I => \N__57119\
        );

    \I__14274\ : InMux
    port map (
            O => \N__57250\,
            I => \N__57116\
        );

    \I__14273\ : LocalMux
    port map (
            O => \N__57243\,
            I => \N__57113\
        );

    \I__14272\ : InMux
    port map (
            O => \N__57242\,
            I => \N__57108\
        );

    \I__14271\ : InMux
    port map (
            O => \N__57241\,
            I => \N__57108\
        );

    \I__14270\ : LocalMux
    port map (
            O => \N__57238\,
            I => \N__57091\
        );

    \I__14269\ : LocalMux
    port map (
            O => \N__57233\,
            I => \N__57091\
        );

    \I__14268\ : LocalMux
    port map (
            O => \N__57230\,
            I => \N__57091\
        );

    \I__14267\ : LocalMux
    port map (
            O => \N__57225\,
            I => \N__57091\
        );

    \I__14266\ : Span4Mux_h
    port map (
            O => \N__57220\,
            I => \N__57091\
        );

    \I__14265\ : Span4Mux_h
    port map (
            O => \N__57215\,
            I => \N__57091\
        );

    \I__14264\ : Span4Mux_v
    port map (
            O => \N__57212\,
            I => \N__57091\
        );

    \I__14263\ : LocalMux
    port map (
            O => \N__57209\,
            I => \N__57091\
        );

    \I__14262\ : Span4Mux_v
    port map (
            O => \N__57206\,
            I => \N__57086\
        );

    \I__14261\ : Span4Mux_h
    port map (
            O => \N__57193\,
            I => \N__57086\
        );

    \I__14260\ : InMux
    port map (
            O => \N__57192\,
            I => \N__57081\
        );

    \I__14259\ : InMux
    port map (
            O => \N__57191\,
            I => \N__57081\
        );

    \I__14258\ : InMux
    port map (
            O => \N__57190\,
            I => \N__57074\
        );

    \I__14257\ : InMux
    port map (
            O => \N__57189\,
            I => \N__57074\
        );

    \I__14256\ : InMux
    port map (
            O => \N__57188\,
            I => \N__57074\
        );

    \I__14255\ : InMux
    port map (
            O => \N__57187\,
            I => \N__57071\
        );

    \I__14254\ : InMux
    port map (
            O => \N__57186\,
            I => \N__57064\
        );

    \I__14253\ : InMux
    port map (
            O => \N__57185\,
            I => \N__57064\
        );

    \I__14252\ : InMux
    port map (
            O => \N__57184\,
            I => \N__57064\
        );

    \I__14251\ : InMux
    port map (
            O => \N__57183\,
            I => \N__57061\
        );

    \I__14250\ : InMux
    port map (
            O => \N__57182\,
            I => \N__57058\
        );

    \I__14249\ : InMux
    port map (
            O => \N__57181\,
            I => \N__57055\
        );

    \I__14248\ : LocalMux
    port map (
            O => \N__57172\,
            I => \N__57050\
        );

    \I__14247\ : Span4Mux_v
    port map (
            O => \N__57163\,
            I => \N__57050\
        );

    \I__14246\ : Span12Mux_v
    port map (
            O => \N__57160\,
            I => \N__57045\
        );

    \I__14245\ : LocalMux
    port map (
            O => \N__57157\,
            I => \N__57045\
        );

    \I__14244\ : Span4Mux_v
    port map (
            O => \N__57154\,
            I => \N__57040\
        );

    \I__14243\ : LocalMux
    port map (
            O => \N__57149\,
            I => \N__57040\
        );

    \I__14242\ : Span4Mux_h
    port map (
            O => \N__57142\,
            I => \N__57037\
        );

    \I__14241\ : Span4Mux_v
    port map (
            O => \N__57135\,
            I => \N__57032\
        );

    \I__14240\ : Span4Mux_h
    port map (
            O => \N__57126\,
            I => \N__57032\
        );

    \I__14239\ : Span12Mux_h
    port map (
            O => \N__57119\,
            I => \N__57029\
        );

    \I__14238\ : LocalMux
    port map (
            O => \N__57116\,
            I => \N__57018\
        );

    \I__14237\ : Span4Mux_h
    port map (
            O => \N__57113\,
            I => \N__57018\
        );

    \I__14236\ : LocalMux
    port map (
            O => \N__57108\,
            I => \N__57018\
        );

    \I__14235\ : Span4Mux_v
    port map (
            O => \N__57091\,
            I => \N__57018\
        );

    \I__14234\ : Span4Mux_h
    port map (
            O => \N__57086\,
            I => \N__57018\
        );

    \I__14233\ : LocalMux
    port map (
            O => \N__57081\,
            I => comm_cmd_1
        );

    \I__14232\ : LocalMux
    port map (
            O => \N__57074\,
            I => comm_cmd_1
        );

    \I__14231\ : LocalMux
    port map (
            O => \N__57071\,
            I => comm_cmd_1
        );

    \I__14230\ : LocalMux
    port map (
            O => \N__57064\,
            I => comm_cmd_1
        );

    \I__14229\ : LocalMux
    port map (
            O => \N__57061\,
            I => comm_cmd_1
        );

    \I__14228\ : LocalMux
    port map (
            O => \N__57058\,
            I => comm_cmd_1
        );

    \I__14227\ : LocalMux
    port map (
            O => \N__57055\,
            I => comm_cmd_1
        );

    \I__14226\ : Odrv4
    port map (
            O => \N__57050\,
            I => comm_cmd_1
        );

    \I__14225\ : Odrv12
    port map (
            O => \N__57045\,
            I => comm_cmd_1
        );

    \I__14224\ : Odrv4
    port map (
            O => \N__57040\,
            I => comm_cmd_1
        );

    \I__14223\ : Odrv4
    port map (
            O => \N__57037\,
            I => comm_cmd_1
        );

    \I__14222\ : Odrv4
    port map (
            O => \N__57032\,
            I => comm_cmd_1
        );

    \I__14221\ : Odrv12
    port map (
            O => \N__57029\,
            I => comm_cmd_1
        );

    \I__14220\ : Odrv4
    port map (
            O => \N__57018\,
            I => comm_cmd_1
        );

    \I__14219\ : InMux
    port map (
            O => \N__56989\,
            I => \N__56985\
        );

    \I__14218\ : InMux
    port map (
            O => \N__56988\,
            I => \N__56979\
        );

    \I__14217\ : LocalMux
    port map (
            O => \N__56985\,
            I => \N__56974\
        );

    \I__14216\ : InMux
    port map (
            O => \N__56984\,
            I => \N__56969\
        );

    \I__14215\ : InMux
    port map (
            O => \N__56983\,
            I => \N__56969\
        );

    \I__14214\ : InMux
    port map (
            O => \N__56982\,
            I => \N__56961\
        );

    \I__14213\ : LocalMux
    port map (
            O => \N__56979\,
            I => \N__56946\
        );

    \I__14212\ : InMux
    port map (
            O => \N__56978\,
            I => \N__56942\
        );

    \I__14211\ : CascadeMux
    port map (
            O => \N__56977\,
            I => \N__56935\
        );

    \I__14210\ : Span4Mux_h
    port map (
            O => \N__56974\,
            I => \N__56922\
        );

    \I__14209\ : LocalMux
    port map (
            O => \N__56969\,
            I => \N__56922\
        );

    \I__14208\ : InMux
    port map (
            O => \N__56968\,
            I => \N__56918\
        );

    \I__14207\ : InMux
    port map (
            O => \N__56967\,
            I => \N__56915\
        );

    \I__14206\ : InMux
    port map (
            O => \N__56966\,
            I => \N__56898\
        );

    \I__14205\ : InMux
    port map (
            O => \N__56965\,
            I => \N__56894\
        );

    \I__14204\ : InMux
    port map (
            O => \N__56964\,
            I => \N__56891\
        );

    \I__14203\ : LocalMux
    port map (
            O => \N__56961\,
            I => \N__56880\
        );

    \I__14202\ : InMux
    port map (
            O => \N__56960\,
            I => \N__56875\
        );

    \I__14201\ : InMux
    port map (
            O => \N__56959\,
            I => \N__56875\
        );

    \I__14200\ : InMux
    port map (
            O => \N__56958\,
            I => \N__56868\
        );

    \I__14199\ : InMux
    port map (
            O => \N__56957\,
            I => \N__56868\
        );

    \I__14198\ : InMux
    port map (
            O => \N__56956\,
            I => \N__56868\
        );

    \I__14197\ : InMux
    port map (
            O => \N__56955\,
            I => \N__56860\
        );

    \I__14196\ : InMux
    port map (
            O => \N__56954\,
            I => \N__56860\
        );

    \I__14195\ : InMux
    port map (
            O => \N__56953\,
            I => \N__56855\
        );

    \I__14194\ : InMux
    port map (
            O => \N__56952\,
            I => \N__56855\
        );

    \I__14193\ : InMux
    port map (
            O => \N__56951\,
            I => \N__56848\
        );

    \I__14192\ : InMux
    port map (
            O => \N__56950\,
            I => \N__56848\
        );

    \I__14191\ : InMux
    port map (
            O => \N__56949\,
            I => \N__56848\
        );

    \I__14190\ : Span4Mux_h
    port map (
            O => \N__56946\,
            I => \N__56845\
        );

    \I__14189\ : InMux
    port map (
            O => \N__56945\,
            I => \N__56842\
        );

    \I__14188\ : LocalMux
    port map (
            O => \N__56942\,
            I => \N__56837\
        );

    \I__14187\ : InMux
    port map (
            O => \N__56941\,
            I => \N__56834\
        );

    \I__14186\ : InMux
    port map (
            O => \N__56940\,
            I => \N__56824\
        );

    \I__14185\ : InMux
    port map (
            O => \N__56939\,
            I => \N__56824\
        );

    \I__14184\ : InMux
    port map (
            O => \N__56938\,
            I => \N__56824\
        );

    \I__14183\ : InMux
    port map (
            O => \N__56935\,
            I => \N__56811\
        );

    \I__14182\ : InMux
    port map (
            O => \N__56934\,
            I => \N__56811\
        );

    \I__14181\ : InMux
    port map (
            O => \N__56933\,
            I => \N__56811\
        );

    \I__14180\ : InMux
    port map (
            O => \N__56932\,
            I => \N__56811\
        );

    \I__14179\ : InMux
    port map (
            O => \N__56931\,
            I => \N__56811\
        );

    \I__14178\ : InMux
    port map (
            O => \N__56930\,
            I => \N__56811\
        );

    \I__14177\ : InMux
    port map (
            O => \N__56929\,
            I => \N__56804\
        );

    \I__14176\ : InMux
    port map (
            O => \N__56928\,
            I => \N__56804\
        );

    \I__14175\ : InMux
    port map (
            O => \N__56927\,
            I => \N__56804\
        );

    \I__14174\ : Span4Mux_v
    port map (
            O => \N__56922\,
            I => \N__56794\
        );

    \I__14173\ : InMux
    port map (
            O => \N__56921\,
            I => \N__56791\
        );

    \I__14172\ : LocalMux
    port map (
            O => \N__56918\,
            I => \N__56786\
        );

    \I__14171\ : LocalMux
    port map (
            O => \N__56915\,
            I => \N__56786\
        );

    \I__14170\ : InMux
    port map (
            O => \N__56914\,
            I => \N__56781\
        );

    \I__14169\ : InMux
    port map (
            O => \N__56913\,
            I => \N__56781\
        );

    \I__14168\ : InMux
    port map (
            O => \N__56912\,
            I => \N__56778\
        );

    \I__14167\ : InMux
    port map (
            O => \N__56911\,
            I => \N__56775\
        );

    \I__14166\ : InMux
    port map (
            O => \N__56910\,
            I => \N__56772\
        );

    \I__14165\ : InMux
    port map (
            O => \N__56909\,
            I => \N__56763\
        );

    \I__14164\ : InMux
    port map (
            O => \N__56908\,
            I => \N__56763\
        );

    \I__14163\ : InMux
    port map (
            O => \N__56907\,
            I => \N__56763\
        );

    \I__14162\ : InMux
    port map (
            O => \N__56906\,
            I => \N__56763\
        );

    \I__14161\ : InMux
    port map (
            O => \N__56905\,
            I => \N__56760\
        );

    \I__14160\ : InMux
    port map (
            O => \N__56904\,
            I => \N__56757\
        );

    \I__14159\ : InMux
    port map (
            O => \N__56903\,
            I => \N__56754\
        );

    \I__14158\ : InMux
    port map (
            O => \N__56902\,
            I => \N__56749\
        );

    \I__14157\ : InMux
    port map (
            O => \N__56901\,
            I => \N__56749\
        );

    \I__14156\ : LocalMux
    port map (
            O => \N__56898\,
            I => \N__56746\
        );

    \I__14155\ : InMux
    port map (
            O => \N__56897\,
            I => \N__56743\
        );

    \I__14154\ : LocalMux
    port map (
            O => \N__56894\,
            I => \N__56738\
        );

    \I__14153\ : LocalMux
    port map (
            O => \N__56891\,
            I => \N__56738\
        );

    \I__14152\ : InMux
    port map (
            O => \N__56890\,
            I => \N__56733\
        );

    \I__14151\ : InMux
    port map (
            O => \N__56889\,
            I => \N__56733\
        );

    \I__14150\ : InMux
    port map (
            O => \N__56888\,
            I => \N__56730\
        );

    \I__14149\ : InMux
    port map (
            O => \N__56887\,
            I => \N__56727\
        );

    \I__14148\ : InMux
    port map (
            O => \N__56886\,
            I => \N__56722\
        );

    \I__14147\ : InMux
    port map (
            O => \N__56885\,
            I => \N__56717\
        );

    \I__14146\ : InMux
    port map (
            O => \N__56884\,
            I => \N__56717\
        );

    \I__14145\ : InMux
    port map (
            O => \N__56883\,
            I => \N__56714\
        );

    \I__14144\ : Span4Mux_h
    port map (
            O => \N__56880\,
            I => \N__56707\
        );

    \I__14143\ : LocalMux
    port map (
            O => \N__56875\,
            I => \N__56707\
        );

    \I__14142\ : LocalMux
    port map (
            O => \N__56868\,
            I => \N__56707\
        );

    \I__14141\ : InMux
    port map (
            O => \N__56867\,
            I => \N__56700\
        );

    \I__14140\ : InMux
    port map (
            O => \N__56866\,
            I => \N__56700\
        );

    \I__14139\ : InMux
    port map (
            O => \N__56865\,
            I => \N__56700\
        );

    \I__14138\ : LocalMux
    port map (
            O => \N__56860\,
            I => \N__56695\
        );

    \I__14137\ : LocalMux
    port map (
            O => \N__56855\,
            I => \N__56690\
        );

    \I__14136\ : LocalMux
    port map (
            O => \N__56848\,
            I => \N__56687\
        );

    \I__14135\ : Span4Mux_v
    port map (
            O => \N__56845\,
            I => \N__56678\
        );

    \I__14134\ : LocalMux
    port map (
            O => \N__56842\,
            I => \N__56678\
        );

    \I__14133\ : InMux
    port map (
            O => \N__56841\,
            I => \N__56675\
        );

    \I__14132\ : InMux
    port map (
            O => \N__56840\,
            I => \N__56672\
        );

    \I__14131\ : Span4Mux_v
    port map (
            O => \N__56837\,
            I => \N__56667\
        );

    \I__14130\ : LocalMux
    port map (
            O => \N__56834\,
            I => \N__56667\
        );

    \I__14129\ : InMux
    port map (
            O => \N__56833\,
            I => \N__56662\
        );

    \I__14128\ : InMux
    port map (
            O => \N__56832\,
            I => \N__56662\
        );

    \I__14127\ : InMux
    port map (
            O => \N__56831\,
            I => \N__56659\
        );

    \I__14126\ : LocalMux
    port map (
            O => \N__56824\,
            I => \N__56652\
        );

    \I__14125\ : LocalMux
    port map (
            O => \N__56811\,
            I => \N__56652\
        );

    \I__14124\ : LocalMux
    port map (
            O => \N__56804\,
            I => \N__56652\
        );

    \I__14123\ : InMux
    port map (
            O => \N__56803\,
            I => \N__56649\
        );

    \I__14122\ : InMux
    port map (
            O => \N__56802\,
            I => \N__56646\
        );

    \I__14121\ : InMux
    port map (
            O => \N__56801\,
            I => \N__56643\
        );

    \I__14120\ : InMux
    port map (
            O => \N__56800\,
            I => \N__56625\
        );

    \I__14119\ : InMux
    port map (
            O => \N__56799\,
            I => \N__56625\
        );

    \I__14118\ : InMux
    port map (
            O => \N__56798\,
            I => \N__56625\
        );

    \I__14117\ : InMux
    port map (
            O => \N__56797\,
            I => \N__56625\
        );

    \I__14116\ : Span4Mux_h
    port map (
            O => \N__56794\,
            I => \N__56616\
        );

    \I__14115\ : LocalMux
    port map (
            O => \N__56791\,
            I => \N__56616\
        );

    \I__14114\ : Span4Mux_v
    port map (
            O => \N__56786\,
            I => \N__56616\
        );

    \I__14113\ : LocalMux
    port map (
            O => \N__56781\,
            I => \N__56616\
        );

    \I__14112\ : LocalMux
    port map (
            O => \N__56778\,
            I => \N__56607\
        );

    \I__14111\ : LocalMux
    port map (
            O => \N__56775\,
            I => \N__56607\
        );

    \I__14110\ : LocalMux
    port map (
            O => \N__56772\,
            I => \N__56607\
        );

    \I__14109\ : LocalMux
    port map (
            O => \N__56763\,
            I => \N__56607\
        );

    \I__14108\ : LocalMux
    port map (
            O => \N__56760\,
            I => \N__56598\
        );

    \I__14107\ : LocalMux
    port map (
            O => \N__56757\,
            I => \N__56598\
        );

    \I__14106\ : LocalMux
    port map (
            O => \N__56754\,
            I => \N__56598\
        );

    \I__14105\ : LocalMux
    port map (
            O => \N__56749\,
            I => \N__56598\
        );

    \I__14104\ : Span4Mux_v
    port map (
            O => \N__56746\,
            I => \N__56595\
        );

    \I__14103\ : LocalMux
    port map (
            O => \N__56743\,
            I => \N__56584\
        );

    \I__14102\ : Span4Mux_v
    port map (
            O => \N__56738\,
            I => \N__56584\
        );

    \I__14101\ : LocalMux
    port map (
            O => \N__56733\,
            I => \N__56584\
        );

    \I__14100\ : LocalMux
    port map (
            O => \N__56730\,
            I => \N__56584\
        );

    \I__14099\ : LocalMux
    port map (
            O => \N__56727\,
            I => \N__56584\
        );

    \I__14098\ : InMux
    port map (
            O => \N__56726\,
            I => \N__56579\
        );

    \I__14097\ : InMux
    port map (
            O => \N__56725\,
            I => \N__56579\
        );

    \I__14096\ : LocalMux
    port map (
            O => \N__56722\,
            I => \N__56568\
        );

    \I__14095\ : LocalMux
    port map (
            O => \N__56717\,
            I => \N__56568\
        );

    \I__14094\ : LocalMux
    port map (
            O => \N__56714\,
            I => \N__56568\
        );

    \I__14093\ : Span4Mux_h
    port map (
            O => \N__56707\,
            I => \N__56568\
        );

    \I__14092\ : LocalMux
    port map (
            O => \N__56700\,
            I => \N__56568\
        );

    \I__14091\ : CascadeMux
    port map (
            O => \N__56699\,
            I => \N__56564\
        );

    \I__14090\ : InMux
    port map (
            O => \N__56698\,
            I => \N__56559\
        );

    \I__14089\ : Span4Mux_h
    port map (
            O => \N__56695\,
            I => \N__56556\
        );

    \I__14088\ : InMux
    port map (
            O => \N__56694\,
            I => \N__56551\
        );

    \I__14087\ : InMux
    port map (
            O => \N__56693\,
            I => \N__56551\
        );

    \I__14086\ : Span4Mux_h
    port map (
            O => \N__56690\,
            I => \N__56546\
        );

    \I__14085\ : Span4Mux_h
    port map (
            O => \N__56687\,
            I => \N__56546\
        );

    \I__14084\ : InMux
    port map (
            O => \N__56686\,
            I => \N__56543\
        );

    \I__14083\ : InMux
    port map (
            O => \N__56685\,
            I => \N__56536\
        );

    \I__14082\ : InMux
    port map (
            O => \N__56684\,
            I => \N__56536\
        );

    \I__14081\ : InMux
    port map (
            O => \N__56683\,
            I => \N__56536\
        );

    \I__14080\ : Span4Mux_h
    port map (
            O => \N__56678\,
            I => \N__56533\
        );

    \I__14079\ : LocalMux
    port map (
            O => \N__56675\,
            I => \N__56528\
        );

    \I__14078\ : LocalMux
    port map (
            O => \N__56672\,
            I => \N__56528\
        );

    \I__14077\ : Span4Mux_h
    port map (
            O => \N__56667\,
            I => \N__56517\
        );

    \I__14076\ : LocalMux
    port map (
            O => \N__56662\,
            I => \N__56517\
        );

    \I__14075\ : LocalMux
    port map (
            O => \N__56659\,
            I => \N__56517\
        );

    \I__14074\ : Span4Mux_v
    port map (
            O => \N__56652\,
            I => \N__56517\
        );

    \I__14073\ : LocalMux
    port map (
            O => \N__56649\,
            I => \N__56517\
        );

    \I__14072\ : LocalMux
    port map (
            O => \N__56646\,
            I => \N__56512\
        );

    \I__14071\ : LocalMux
    port map (
            O => \N__56643\,
            I => \N__56512\
        );

    \I__14070\ : InMux
    port map (
            O => \N__56642\,
            I => \N__56509\
        );

    \I__14069\ : InMux
    port map (
            O => \N__56641\,
            I => \N__56502\
        );

    \I__14068\ : InMux
    port map (
            O => \N__56640\,
            I => \N__56502\
        );

    \I__14067\ : InMux
    port map (
            O => \N__56639\,
            I => \N__56502\
        );

    \I__14066\ : InMux
    port map (
            O => \N__56638\,
            I => \N__56499\
        );

    \I__14065\ : InMux
    port map (
            O => \N__56637\,
            I => \N__56490\
        );

    \I__14064\ : InMux
    port map (
            O => \N__56636\,
            I => \N__56490\
        );

    \I__14063\ : InMux
    port map (
            O => \N__56635\,
            I => \N__56490\
        );

    \I__14062\ : InMux
    port map (
            O => \N__56634\,
            I => \N__56490\
        );

    \I__14061\ : LocalMux
    port map (
            O => \N__56625\,
            I => \N__56487\
        );

    \I__14060\ : Span4Mux_v
    port map (
            O => \N__56616\,
            I => \N__56480\
        );

    \I__14059\ : Span4Mux_v
    port map (
            O => \N__56607\,
            I => \N__56480\
        );

    \I__14058\ : Span4Mux_v
    port map (
            O => \N__56598\,
            I => \N__56480\
        );

    \I__14057\ : Span4Mux_h
    port map (
            O => \N__56595\,
            I => \N__56471\
        );

    \I__14056\ : Span4Mux_v
    port map (
            O => \N__56584\,
            I => \N__56471\
        );

    \I__14055\ : LocalMux
    port map (
            O => \N__56579\,
            I => \N__56471\
        );

    \I__14054\ : Span4Mux_v
    port map (
            O => \N__56568\,
            I => \N__56471\
        );

    \I__14053\ : InMux
    port map (
            O => \N__56567\,
            I => \N__56462\
        );

    \I__14052\ : InMux
    port map (
            O => \N__56564\,
            I => \N__56462\
        );

    \I__14051\ : InMux
    port map (
            O => \N__56563\,
            I => \N__56462\
        );

    \I__14050\ : InMux
    port map (
            O => \N__56562\,
            I => \N__56462\
        );

    \I__14049\ : LocalMux
    port map (
            O => \N__56559\,
            I => \N__56451\
        );

    \I__14048\ : Span4Mux_h
    port map (
            O => \N__56556\,
            I => \N__56451\
        );

    \I__14047\ : LocalMux
    port map (
            O => \N__56551\,
            I => \N__56451\
        );

    \I__14046\ : Span4Mux_h
    port map (
            O => \N__56546\,
            I => \N__56451\
        );

    \I__14045\ : LocalMux
    port map (
            O => \N__56543\,
            I => \N__56451\
        );

    \I__14044\ : LocalMux
    port map (
            O => \N__56536\,
            I => \N__56446\
        );

    \I__14043\ : Span4Mux_h
    port map (
            O => \N__56533\,
            I => \N__56446\
        );

    \I__14042\ : Span4Mux_v
    port map (
            O => \N__56528\,
            I => \N__56441\
        );

    \I__14041\ : Span4Mux_h
    port map (
            O => \N__56517\,
            I => \N__56441\
        );

    \I__14040\ : Odrv12
    port map (
            O => \N__56512\,
            I => comm_cmd_0
        );

    \I__14039\ : LocalMux
    port map (
            O => \N__56509\,
            I => comm_cmd_0
        );

    \I__14038\ : LocalMux
    port map (
            O => \N__56502\,
            I => comm_cmd_0
        );

    \I__14037\ : LocalMux
    port map (
            O => \N__56499\,
            I => comm_cmd_0
        );

    \I__14036\ : LocalMux
    port map (
            O => \N__56490\,
            I => comm_cmd_0
        );

    \I__14035\ : Odrv4
    port map (
            O => \N__56487\,
            I => comm_cmd_0
        );

    \I__14034\ : Odrv4
    port map (
            O => \N__56480\,
            I => comm_cmd_0
        );

    \I__14033\ : Odrv4
    port map (
            O => \N__56471\,
            I => comm_cmd_0
        );

    \I__14032\ : LocalMux
    port map (
            O => \N__56462\,
            I => comm_cmd_0
        );

    \I__14031\ : Odrv4
    port map (
            O => \N__56451\,
            I => comm_cmd_0
        );

    \I__14030\ : Odrv4
    port map (
            O => \N__56446\,
            I => comm_cmd_0
        );

    \I__14029\ : Odrv4
    port map (
            O => \N__56441\,
            I => comm_cmd_0
        );

    \I__14028\ : CascadeMux
    port map (
            O => \N__56416\,
            I => \N__56413\
        );

    \I__14027\ : InMux
    port map (
            O => \N__56413\,
            I => \N__56410\
        );

    \I__14026\ : LocalMux
    port map (
            O => \N__56410\,
            I => \N__56407\
        );

    \I__14025\ : Span4Mux_v
    port map (
            O => \N__56407\,
            I => \N__56404\
        );

    \I__14024\ : Odrv4
    port map (
            O => \N__56404\,
            I => n23_adj_1517
        );

    \I__14023\ : InMux
    port map (
            O => \N__56401\,
            I => \N__56398\
        );

    \I__14022\ : LocalMux
    port map (
            O => \N__56398\,
            I => \N__56394\
        );

    \I__14021\ : InMux
    port map (
            O => \N__56397\,
            I => \N__56391\
        );

    \I__14020\ : Span4Mux_h
    port map (
            O => \N__56394\,
            I => \N__56388\
        );

    \I__14019\ : LocalMux
    port map (
            O => \N__56391\,
            I => \N__56382\
        );

    \I__14018\ : Span4Mux_v
    port map (
            O => \N__56388\,
            I => \N__56382\
        );

    \I__14017\ : InMux
    port map (
            O => \N__56387\,
            I => \N__56379\
        );

    \I__14016\ : Odrv4
    port map (
            O => \N__56382\,
            I => req_data_cnt_12
        );

    \I__14015\ : LocalMux
    port map (
            O => \N__56379\,
            I => req_data_cnt_12
        );

    \I__14014\ : InMux
    port map (
            O => \N__56374\,
            I => \N__56371\
        );

    \I__14013\ : LocalMux
    port map (
            O => \N__56371\,
            I => \N__56368\
        );

    \I__14012\ : Span12Mux_v
    port map (
            O => \N__56368\,
            I => \N__56365\
        );

    \I__14011\ : Odrv12
    port map (
            O => \N__56365\,
            I => n20809
        );

    \I__14010\ : InMux
    port map (
            O => \N__56362\,
            I => \N__56359\
        );

    \I__14009\ : LocalMux
    port map (
            O => \N__56359\,
            I => \N__56356\
        );

    \I__14008\ : Odrv4
    port map (
            O => \N__56356\,
            I => n17415
        );

    \I__14007\ : InMux
    port map (
            O => \N__56353\,
            I => \N__56350\
        );

    \I__14006\ : LocalMux
    port map (
            O => \N__56350\,
            I => buf_data_iac_4
        );

    \I__14005\ : InMux
    port map (
            O => \N__56347\,
            I => \N__56331\
        );

    \I__14004\ : InMux
    port map (
            O => \N__56346\,
            I => \N__56326\
        );

    \I__14003\ : InMux
    port map (
            O => \N__56345\,
            I => \N__56326\
        );

    \I__14002\ : InMux
    port map (
            O => \N__56344\,
            I => \N__56321\
        );

    \I__14001\ : InMux
    port map (
            O => \N__56343\,
            I => \N__56321\
        );

    \I__14000\ : CascadeMux
    port map (
            O => \N__56342\,
            I => \N__56318\
        );

    \I__13999\ : CascadeMux
    port map (
            O => \N__56341\,
            I => \N__56312\
        );

    \I__13998\ : InMux
    port map (
            O => \N__56340\,
            I => \N__56301\
        );

    \I__13997\ : InMux
    port map (
            O => \N__56339\,
            I => \N__56301\
        );

    \I__13996\ : InMux
    port map (
            O => \N__56338\,
            I => \N__56301\
        );

    \I__13995\ : InMux
    port map (
            O => \N__56337\,
            I => \N__56296\
        );

    \I__13994\ : InMux
    port map (
            O => \N__56336\,
            I => \N__56296\
        );

    \I__13993\ : InMux
    port map (
            O => \N__56335\,
            I => \N__56291\
        );

    \I__13992\ : InMux
    port map (
            O => \N__56334\,
            I => \N__56291\
        );

    \I__13991\ : LocalMux
    port map (
            O => \N__56331\,
            I => \N__56284\
        );

    \I__13990\ : LocalMux
    port map (
            O => \N__56326\,
            I => \N__56281\
        );

    \I__13989\ : LocalMux
    port map (
            O => \N__56321\,
            I => \N__56278\
        );

    \I__13988\ : InMux
    port map (
            O => \N__56318\,
            I => \N__56275\
        );

    \I__13987\ : InMux
    port map (
            O => \N__56317\,
            I => \N__56266\
        );

    \I__13986\ : InMux
    port map (
            O => \N__56316\,
            I => \N__56261\
        );

    \I__13985\ : InMux
    port map (
            O => \N__56315\,
            I => \N__56253\
        );

    \I__13984\ : InMux
    port map (
            O => \N__56312\,
            I => \N__56248\
        );

    \I__13983\ : InMux
    port map (
            O => \N__56311\,
            I => \N__56248\
        );

    \I__13982\ : InMux
    port map (
            O => \N__56310\,
            I => \N__56245\
        );

    \I__13981\ : InMux
    port map (
            O => \N__56309\,
            I => \N__56240\
        );

    \I__13980\ : InMux
    port map (
            O => \N__56308\,
            I => \N__56240\
        );

    \I__13979\ : LocalMux
    port map (
            O => \N__56301\,
            I => \N__56233\
        );

    \I__13978\ : LocalMux
    port map (
            O => \N__56296\,
            I => \N__56233\
        );

    \I__13977\ : LocalMux
    port map (
            O => \N__56291\,
            I => \N__56233\
        );

    \I__13976\ : InMux
    port map (
            O => \N__56290\,
            I => \N__56228\
        );

    \I__13975\ : InMux
    port map (
            O => \N__56289\,
            I => \N__56228\
        );

    \I__13974\ : InMux
    port map (
            O => \N__56288\,
            I => \N__56225\
        );

    \I__13973\ : InMux
    port map (
            O => \N__56287\,
            I => \N__56222\
        );

    \I__13972\ : Span4Mux_h
    port map (
            O => \N__56284\,
            I => \N__56213\
        );

    \I__13971\ : Span4Mux_h
    port map (
            O => \N__56281\,
            I => \N__56213\
        );

    \I__13970\ : Span4Mux_v
    port map (
            O => \N__56278\,
            I => \N__56213\
        );

    \I__13969\ : LocalMux
    port map (
            O => \N__56275\,
            I => \N__56213\
        );

    \I__13968\ : InMux
    port map (
            O => \N__56274\,
            I => \N__56210\
        );

    \I__13967\ : InMux
    port map (
            O => \N__56273\,
            I => \N__56207\
        );

    \I__13966\ : InMux
    port map (
            O => \N__56272\,
            I => \N__56204\
        );

    \I__13965\ : InMux
    port map (
            O => \N__56271\,
            I => \N__56201\
        );

    \I__13964\ : InMux
    port map (
            O => \N__56270\,
            I => \N__56198\
        );

    \I__13963\ : InMux
    port map (
            O => \N__56269\,
            I => \N__56195\
        );

    \I__13962\ : LocalMux
    port map (
            O => \N__56266\,
            I => \N__56192\
        );

    \I__13961\ : InMux
    port map (
            O => \N__56265\,
            I => \N__56187\
        );

    \I__13960\ : InMux
    port map (
            O => \N__56264\,
            I => \N__56187\
        );

    \I__13959\ : LocalMux
    port map (
            O => \N__56261\,
            I => \N__56184\
        );

    \I__13958\ : InMux
    port map (
            O => \N__56260\,
            I => \N__56181\
        );

    \I__13957\ : InMux
    port map (
            O => \N__56259\,
            I => \N__56176\
        );

    \I__13956\ : InMux
    port map (
            O => \N__56258\,
            I => \N__56176\
        );

    \I__13955\ : InMux
    port map (
            O => \N__56257\,
            I => \N__56173\
        );

    \I__13954\ : InMux
    port map (
            O => \N__56256\,
            I => \N__56170\
        );

    \I__13953\ : LocalMux
    port map (
            O => \N__56253\,
            I => \N__56166\
        );

    \I__13952\ : LocalMux
    port map (
            O => \N__56248\,
            I => \N__56161\
        );

    \I__13951\ : LocalMux
    port map (
            O => \N__56245\,
            I => \N__56161\
        );

    \I__13950\ : LocalMux
    port map (
            O => \N__56240\,
            I => \N__56156\
        );

    \I__13949\ : Span4Mux_v
    port map (
            O => \N__56233\,
            I => \N__56156\
        );

    \I__13948\ : LocalMux
    port map (
            O => \N__56228\,
            I => \N__56147\
        );

    \I__13947\ : LocalMux
    port map (
            O => \N__56225\,
            I => \N__56147\
        );

    \I__13946\ : LocalMux
    port map (
            O => \N__56222\,
            I => \N__56147\
        );

    \I__13945\ : Span4Mux_h
    port map (
            O => \N__56213\,
            I => \N__56147\
        );

    \I__13944\ : LocalMux
    port map (
            O => \N__56210\,
            I => \N__56139\
        );

    \I__13943\ : LocalMux
    port map (
            O => \N__56207\,
            I => \N__56139\
        );

    \I__13942\ : LocalMux
    port map (
            O => \N__56204\,
            I => \N__56134\
        );

    \I__13941\ : LocalMux
    port map (
            O => \N__56201\,
            I => \N__56134\
        );

    \I__13940\ : LocalMux
    port map (
            O => \N__56198\,
            I => \N__56131\
        );

    \I__13939\ : LocalMux
    port map (
            O => \N__56195\,
            I => \N__56118\
        );

    \I__13938\ : Span4Mux_v
    port map (
            O => \N__56192\,
            I => \N__56118\
        );

    \I__13937\ : LocalMux
    port map (
            O => \N__56187\,
            I => \N__56118\
        );

    \I__13936\ : Span4Mux_h
    port map (
            O => \N__56184\,
            I => \N__56118\
        );

    \I__13935\ : LocalMux
    port map (
            O => \N__56181\,
            I => \N__56118\
        );

    \I__13934\ : LocalMux
    port map (
            O => \N__56176\,
            I => \N__56118\
        );

    \I__13933\ : LocalMux
    port map (
            O => \N__56173\,
            I => \N__56115\
        );

    \I__13932\ : LocalMux
    port map (
            O => \N__56170\,
            I => \N__56112\
        );

    \I__13931\ : InMux
    port map (
            O => \N__56169\,
            I => \N__56109\
        );

    \I__13930\ : Span4Mux_v
    port map (
            O => \N__56166\,
            I => \N__56106\
        );

    \I__13929\ : Span12Mux_h
    port map (
            O => \N__56161\,
            I => \N__56103\
        );

    \I__13928\ : Span4Mux_h
    port map (
            O => \N__56156\,
            I => \N__56098\
        );

    \I__13927\ : Span4Mux_v
    port map (
            O => \N__56147\,
            I => \N__56098\
        );

    \I__13926\ : InMux
    port map (
            O => \N__56146\,
            I => \N__56091\
        );

    \I__13925\ : InMux
    port map (
            O => \N__56145\,
            I => \N__56091\
        );

    \I__13924\ : InMux
    port map (
            O => \N__56144\,
            I => \N__56091\
        );

    \I__13923\ : Span4Mux_v
    port map (
            O => \N__56139\,
            I => \N__56082\
        );

    \I__13922\ : Span4Mux_h
    port map (
            O => \N__56134\,
            I => \N__56082\
        );

    \I__13921\ : Span4Mux_v
    port map (
            O => \N__56131\,
            I => \N__56082\
        );

    \I__13920\ : Span4Mux_v
    port map (
            O => \N__56118\,
            I => \N__56082\
        );

    \I__13919\ : Odrv12
    port map (
            O => \N__56115\,
            I => comm_cmd_3
        );

    \I__13918\ : Odrv4
    port map (
            O => \N__56112\,
            I => comm_cmd_3
        );

    \I__13917\ : LocalMux
    port map (
            O => \N__56109\,
            I => comm_cmd_3
        );

    \I__13916\ : Odrv4
    port map (
            O => \N__56106\,
            I => comm_cmd_3
        );

    \I__13915\ : Odrv12
    port map (
            O => \N__56103\,
            I => comm_cmd_3
        );

    \I__13914\ : Odrv4
    port map (
            O => \N__56098\,
            I => comm_cmd_3
        );

    \I__13913\ : LocalMux
    port map (
            O => \N__56091\,
            I => comm_cmd_3
        );

    \I__13912\ : Odrv4
    port map (
            O => \N__56082\,
            I => comm_cmd_3
        );

    \I__13911\ : InMux
    port map (
            O => \N__56065\,
            I => \N__56062\
        );

    \I__13910\ : LocalMux
    port map (
            O => \N__56062\,
            I => \N__56059\
        );

    \I__13909\ : Span4Mux_h
    port map (
            O => \N__56059\,
            I => \N__56056\
        );

    \I__13908\ : Odrv4
    port map (
            O => \N__56056\,
            I => n22_adj_1606
        );

    \I__13907\ : InMux
    port map (
            O => \N__56053\,
            I => \N__56050\
        );

    \I__13906\ : LocalMux
    port map (
            O => \N__56050\,
            I => \N__56047\
        );

    \I__13905\ : Span12Mux_v
    port map (
            O => \N__56047\,
            I => \N__56044\
        );

    \I__13904\ : Odrv12
    port map (
            O => \N__56044\,
            I => n30_adj_1608
        );

    \I__13903\ : InMux
    port map (
            O => \N__56041\,
            I => \N__56037\
        );

    \I__13902\ : InMux
    port map (
            O => \N__56040\,
            I => \N__56034\
        );

    \I__13901\ : LocalMux
    port map (
            O => \N__56037\,
            I => \N__56031\
        );

    \I__13900\ : LocalMux
    port map (
            O => \N__56034\,
            I => \N__56019\
        );

    \I__13899\ : Glb2LocalMux
    port map (
            O => \N__56031\,
            I => \N__55984\
        );

    \I__13898\ : ClkMux
    port map (
            O => \N__56030\,
            I => \N__55984\
        );

    \I__13897\ : ClkMux
    port map (
            O => \N__56029\,
            I => \N__55984\
        );

    \I__13896\ : ClkMux
    port map (
            O => \N__56028\,
            I => \N__55984\
        );

    \I__13895\ : ClkMux
    port map (
            O => \N__56027\,
            I => \N__55984\
        );

    \I__13894\ : ClkMux
    port map (
            O => \N__56026\,
            I => \N__55984\
        );

    \I__13893\ : ClkMux
    port map (
            O => \N__56025\,
            I => \N__55984\
        );

    \I__13892\ : ClkMux
    port map (
            O => \N__56024\,
            I => \N__55984\
        );

    \I__13891\ : ClkMux
    port map (
            O => \N__56023\,
            I => \N__55984\
        );

    \I__13890\ : ClkMux
    port map (
            O => \N__56022\,
            I => \N__55984\
        );

    \I__13889\ : Glb2LocalMux
    port map (
            O => \N__56019\,
            I => \N__55984\
        );

    \I__13888\ : ClkMux
    port map (
            O => \N__56018\,
            I => \N__55984\
        );

    \I__13887\ : ClkMux
    port map (
            O => \N__56017\,
            I => \N__55984\
        );

    \I__13886\ : ClkMux
    port map (
            O => \N__56016\,
            I => \N__55984\
        );

    \I__13885\ : ClkMux
    port map (
            O => \N__56015\,
            I => \N__55984\
        );

    \I__13884\ : GlobalMux
    port map (
            O => \N__55984\,
            I => \clk_16MHz\
        );

    \I__13883\ : InMux
    port map (
            O => \N__55981\,
            I => \N__55978\
        );

    \I__13882\ : LocalMux
    port map (
            O => \N__55978\,
            I => \N__55974\
        );

    \I__13881\ : InMux
    port map (
            O => \N__55977\,
            I => \N__55971\
        );

    \I__13880\ : Odrv12
    port map (
            O => \N__55974\,
            I => dds0_mclk
        );

    \I__13879\ : LocalMux
    port map (
            O => \N__55971\,
            I => dds0_mclk
        );

    \I__13878\ : InMux
    port map (
            O => \N__55966\,
            I => \N__55963\
        );

    \I__13877\ : LocalMux
    port map (
            O => \N__55963\,
            I => \N__55959\
        );

    \I__13876\ : InMux
    port map (
            O => \N__55962\,
            I => \N__55956\
        );

    \I__13875\ : Span4Mux_h
    port map (
            O => \N__55959\,
            I => \N__55953\
        );

    \I__13874\ : LocalMux
    port map (
            O => \N__55956\,
            I => \N__55950\
        );

    \I__13873\ : Span4Mux_h
    port map (
            O => \N__55953\,
            I => \N__55944\
        );

    \I__13872\ : Span4Mux_h
    port map (
            O => \N__55950\,
            I => \N__55944\
        );

    \I__13871\ : InMux
    port map (
            O => \N__55949\,
            I => \N__55941\
        );

    \I__13870\ : Span4Mux_h
    port map (
            O => \N__55944\,
            I => \N__55938\
        );

    \I__13869\ : LocalMux
    port map (
            O => \N__55941\,
            I => buf_control_6
        );

    \I__13868\ : Odrv4
    port map (
            O => \N__55938\,
            I => buf_control_6
        );

    \I__13867\ : IoInMux
    port map (
            O => \N__55933\,
            I => \N__55930\
        );

    \I__13866\ : LocalMux
    port map (
            O => \N__55930\,
            I => \N__55927\
        );

    \I__13865\ : Span4Mux_s3_v
    port map (
            O => \N__55927\,
            I => \N__55924\
        );

    \I__13864\ : Sp12to4
    port map (
            O => \N__55924\,
            I => \N__55921\
        );

    \I__13863\ : Span12Mux_s8_h
    port map (
            O => \N__55921\,
            I => \N__55918\
        );

    \I__13862\ : Odrv12
    port map (
            O => \N__55918\,
            I => \DDS_MCLK\
        );

    \I__13861\ : IoInMux
    port map (
            O => \N__55915\,
            I => \N__55912\
        );

    \I__13860\ : LocalMux
    port map (
            O => \N__55912\,
            I => \N__55909\
        );

    \I__13859\ : Span4Mux_s1_v
    port map (
            O => \N__55909\,
            I => \N__55906\
        );

    \I__13858\ : Sp12to4
    port map (
            O => \N__55906\,
            I => \N__55902\
        );

    \I__13857\ : CascadeMux
    port map (
            O => \N__55905\,
            I => \N__55899\
        );

    \I__13856\ : Span12Mux_s8_h
    port map (
            O => \N__55902\,
            I => \N__55896\
        );

    \I__13855\ : InMux
    port map (
            O => \N__55899\,
            I => \N__55893\
        );

    \I__13854\ : Odrv12
    port map (
            O => \N__55896\,
            I => \DDS_SCK\
        );

    \I__13853\ : LocalMux
    port map (
            O => \N__55893\,
            I => \DDS_SCK\
        );

    \I__13852\ : CascadeMux
    port map (
            O => \N__55888\,
            I => \N__55875\
        );

    \I__13851\ : InMux
    port map (
            O => \N__55887\,
            I => \N__55863\
        );

    \I__13850\ : InMux
    port map (
            O => \N__55886\,
            I => \N__55845\
        );

    \I__13849\ : InMux
    port map (
            O => \N__55885\,
            I => \N__55845\
        );

    \I__13848\ : InMux
    port map (
            O => \N__55884\,
            I => \N__55845\
        );

    \I__13847\ : InMux
    port map (
            O => \N__55883\,
            I => \N__55845\
        );

    \I__13846\ : InMux
    port map (
            O => \N__55882\,
            I => \N__55845\
        );

    \I__13845\ : InMux
    port map (
            O => \N__55881\,
            I => \N__55845\
        );

    \I__13844\ : InMux
    port map (
            O => \N__55880\,
            I => \N__55845\
        );

    \I__13843\ : InMux
    port map (
            O => \N__55879\,
            I => \N__55840\
        );

    \I__13842\ : InMux
    port map (
            O => \N__55878\,
            I => \N__55840\
        );

    \I__13841\ : InMux
    port map (
            O => \N__55875\,
            I => \N__55833\
        );

    \I__13840\ : InMux
    port map (
            O => \N__55874\,
            I => \N__55833\
        );

    \I__13839\ : InMux
    port map (
            O => \N__55873\,
            I => \N__55833\
        );

    \I__13838\ : InMux
    port map (
            O => \N__55872\,
            I => \N__55827\
        );

    \I__13837\ : InMux
    port map (
            O => \N__55871\,
            I => \N__55827\
        );

    \I__13836\ : InMux
    port map (
            O => \N__55870\,
            I => \N__55816\
        );

    \I__13835\ : InMux
    port map (
            O => \N__55869\,
            I => \N__55816\
        );

    \I__13834\ : InMux
    port map (
            O => \N__55868\,
            I => \N__55816\
        );

    \I__13833\ : InMux
    port map (
            O => \N__55867\,
            I => \N__55816\
        );

    \I__13832\ : InMux
    port map (
            O => \N__55866\,
            I => \N__55816\
        );

    \I__13831\ : LocalMux
    port map (
            O => \N__55863\,
            I => \N__55813\
        );

    \I__13830\ : InMux
    port map (
            O => \N__55862\,
            I => \N__55810\
        );

    \I__13829\ : InMux
    port map (
            O => \N__55861\,
            I => \N__55807\
        );

    \I__13828\ : InMux
    port map (
            O => \N__55860\,
            I => \N__55804\
        );

    \I__13827\ : LocalMux
    port map (
            O => \N__55845\,
            I => \N__55801\
        );

    \I__13826\ : LocalMux
    port map (
            O => \N__55840\,
            I => \N__55796\
        );

    \I__13825\ : LocalMux
    port map (
            O => \N__55833\,
            I => \N__55796\
        );

    \I__13824\ : InMux
    port map (
            O => \N__55832\,
            I => \N__55792\
        );

    \I__13823\ : LocalMux
    port map (
            O => \N__55827\,
            I => \N__55787\
        );

    \I__13822\ : LocalMux
    port map (
            O => \N__55816\,
            I => \N__55787\
        );

    \I__13821\ : Span4Mux_h
    port map (
            O => \N__55813\,
            I => \N__55784\
        );

    \I__13820\ : LocalMux
    port map (
            O => \N__55810\,
            I => \N__55781\
        );

    \I__13819\ : LocalMux
    port map (
            O => \N__55807\,
            I => \N__55776\
        );

    \I__13818\ : LocalMux
    port map (
            O => \N__55804\,
            I => \N__55776\
        );

    \I__13817\ : Span4Mux_v
    port map (
            O => \N__55801\,
            I => \N__55771\
        );

    \I__13816\ : Span4Mux_v
    port map (
            O => \N__55796\,
            I => \N__55771\
        );

    \I__13815\ : InMux
    port map (
            O => \N__55795\,
            I => \N__55768\
        );

    \I__13814\ : LocalMux
    port map (
            O => \N__55792\,
            I => \N__55765\
        );

    \I__13813\ : Span4Mux_v
    port map (
            O => \N__55787\,
            I => \N__55760\
        );

    \I__13812\ : Span4Mux_h
    port map (
            O => \N__55784\,
            I => \N__55760\
        );

    \I__13811\ : Span4Mux_v
    port map (
            O => \N__55781\,
            I => \N__55753\
        );

    \I__13810\ : Span4Mux_v
    port map (
            O => \N__55776\,
            I => \N__55753\
        );

    \I__13809\ : Span4Mux_h
    port map (
            O => \N__55771\,
            I => \N__55753\
        );

    \I__13808\ : LocalMux
    port map (
            O => \N__55768\,
            I => dds_state_2
        );

    \I__13807\ : Odrv4
    port map (
            O => \N__55765\,
            I => dds_state_2
        );

    \I__13806\ : Odrv4
    port map (
            O => \N__55760\,
            I => dds_state_2
        );

    \I__13805\ : Odrv4
    port map (
            O => \N__55753\,
            I => dds_state_2
        );

    \I__13804\ : InMux
    port map (
            O => \N__55744\,
            I => \N__55741\
        );

    \I__13803\ : LocalMux
    port map (
            O => \N__55741\,
            I => \N__55734\
        );

    \I__13802\ : InMux
    port map (
            O => \N__55740\,
            I => \N__55731\
        );

    \I__13801\ : InMux
    port map (
            O => \N__55739\,
            I => \N__55728\
        );

    \I__13800\ : InMux
    port map (
            O => \N__55738\,
            I => \N__55725\
        );

    \I__13799\ : InMux
    port map (
            O => \N__55737\,
            I => \N__55722\
        );

    \I__13798\ : Span4Mux_v
    port map (
            O => \N__55734\,
            I => \N__55713\
        );

    \I__13797\ : LocalMux
    port map (
            O => \N__55731\,
            I => \N__55713\
        );

    \I__13796\ : LocalMux
    port map (
            O => \N__55728\,
            I => \N__55713\
        );

    \I__13795\ : LocalMux
    port map (
            O => \N__55725\,
            I => \N__55713\
        );

    \I__13794\ : LocalMux
    port map (
            O => \N__55722\,
            I => \N__55708\
        );

    \I__13793\ : Span4Mux_h
    port map (
            O => \N__55713\,
            I => \N__55705\
        );

    \I__13792\ : InMux
    port map (
            O => \N__55712\,
            I => \N__55700\
        );

    \I__13791\ : InMux
    port map (
            O => \N__55711\,
            I => \N__55700\
        );

    \I__13790\ : Span4Mux_v
    port map (
            O => \N__55708\,
            I => \N__55697\
        );

    \I__13789\ : Span4Mux_h
    port map (
            O => \N__55705\,
            I => \N__55690\
        );

    \I__13788\ : LocalMux
    port map (
            O => \N__55700\,
            I => \N__55690\
        );

    \I__13787\ : Span4Mux_h
    port map (
            O => \N__55697\,
            I => \N__55687\
        );

    \I__13786\ : InMux
    port map (
            O => \N__55696\,
            I => \N__55682\
        );

    \I__13785\ : InMux
    port map (
            O => \N__55695\,
            I => \N__55682\
        );

    \I__13784\ : Span4Mux_v
    port map (
            O => \N__55690\,
            I => \N__55679\
        );

    \I__13783\ : Odrv4
    port map (
            O => \N__55687\,
            I => dds_state_0
        );

    \I__13782\ : LocalMux
    port map (
            O => \N__55682\,
            I => dds_state_0
        );

    \I__13781\ : Odrv4
    port map (
            O => \N__55679\,
            I => dds_state_0
        );

    \I__13780\ : CEMux
    port map (
            O => \N__55672\,
            I => \N__55669\
        );

    \I__13779\ : LocalMux
    port map (
            O => \N__55669\,
            I => \N__55656\
        );

    \I__13778\ : InMux
    port map (
            O => \N__55668\,
            I => \N__55640\
        );

    \I__13777\ : InMux
    port map (
            O => \N__55667\,
            I => \N__55640\
        );

    \I__13776\ : InMux
    port map (
            O => \N__55666\,
            I => \N__55640\
        );

    \I__13775\ : InMux
    port map (
            O => \N__55665\,
            I => \N__55640\
        );

    \I__13774\ : InMux
    port map (
            O => \N__55664\,
            I => \N__55640\
        );

    \I__13773\ : InMux
    port map (
            O => \N__55663\,
            I => \N__55640\
        );

    \I__13772\ : InMux
    port map (
            O => \N__55662\,
            I => \N__55640\
        );

    \I__13771\ : InMux
    port map (
            O => \N__55661\,
            I => \N__55635\
        );

    \I__13770\ : InMux
    port map (
            O => \N__55660\,
            I => \N__55635\
        );

    \I__13769\ : SRMux
    port map (
            O => \N__55659\,
            I => \N__55623\
        );

    \I__13768\ : Span4Mux_v
    port map (
            O => \N__55656\,
            I => \N__55617\
        );

    \I__13767\ : InMux
    port map (
            O => \N__55655\,
            I => \N__55614\
        );

    \I__13766\ : LocalMux
    port map (
            O => \N__55640\,
            I => \N__55608\
        );

    \I__13765\ : LocalMux
    port map (
            O => \N__55635\,
            I => \N__55608\
        );

    \I__13764\ : InMux
    port map (
            O => \N__55634\,
            I => \N__55603\
        );

    \I__13763\ : InMux
    port map (
            O => \N__55633\,
            I => \N__55603\
        );

    \I__13762\ : InMux
    port map (
            O => \N__55632\,
            I => \N__55592\
        );

    \I__13761\ : InMux
    port map (
            O => \N__55631\,
            I => \N__55592\
        );

    \I__13760\ : InMux
    port map (
            O => \N__55630\,
            I => \N__55592\
        );

    \I__13759\ : InMux
    port map (
            O => \N__55629\,
            I => \N__55592\
        );

    \I__13758\ : InMux
    port map (
            O => \N__55628\,
            I => \N__55592\
        );

    \I__13757\ : InMux
    port map (
            O => \N__55627\,
            I => \N__55589\
        );

    \I__13756\ : InMux
    port map (
            O => \N__55626\,
            I => \N__55586\
        );

    \I__13755\ : LocalMux
    port map (
            O => \N__55623\,
            I => \N__55582\
        );

    \I__13754\ : InMux
    port map (
            O => \N__55622\,
            I => \N__55579\
        );

    \I__13753\ : InMux
    port map (
            O => \N__55621\,
            I => \N__55574\
        );

    \I__13752\ : InMux
    port map (
            O => \N__55620\,
            I => \N__55574\
        );

    \I__13751\ : Span4Mux_h
    port map (
            O => \N__55617\,
            I => \N__55571\
        );

    \I__13750\ : LocalMux
    port map (
            O => \N__55614\,
            I => \N__55568\
        );

    \I__13749\ : InMux
    port map (
            O => \N__55613\,
            I => \N__55563\
        );

    \I__13748\ : Span4Mux_h
    port map (
            O => \N__55608\,
            I => \N__55556\
        );

    \I__13747\ : LocalMux
    port map (
            O => \N__55603\,
            I => \N__55556\
        );

    \I__13746\ : LocalMux
    port map (
            O => \N__55592\,
            I => \N__55556\
        );

    \I__13745\ : LocalMux
    port map (
            O => \N__55589\,
            I => \N__55553\
        );

    \I__13744\ : LocalMux
    port map (
            O => \N__55586\,
            I => \N__55550\
        );

    \I__13743\ : InMux
    port map (
            O => \N__55585\,
            I => \N__55547\
        );

    \I__13742\ : Span4Mux_h
    port map (
            O => \N__55582\,
            I => \N__55540\
        );

    \I__13741\ : LocalMux
    port map (
            O => \N__55579\,
            I => \N__55540\
        );

    \I__13740\ : LocalMux
    port map (
            O => \N__55574\,
            I => \N__55540\
        );

    \I__13739\ : Span4Mux_h
    port map (
            O => \N__55571\,
            I => \N__55537\
        );

    \I__13738\ : Span12Mux_h
    port map (
            O => \N__55568\,
            I => \N__55534\
        );

    \I__13737\ : InMux
    port map (
            O => \N__55567\,
            I => \N__55529\
        );

    \I__13736\ : InMux
    port map (
            O => \N__55566\,
            I => \N__55529\
        );

    \I__13735\ : LocalMux
    port map (
            O => \N__55563\,
            I => \N__55524\
        );

    \I__13734\ : Span4Mux_h
    port map (
            O => \N__55556\,
            I => \N__55524\
        );

    \I__13733\ : Span4Mux_v
    port map (
            O => \N__55553\,
            I => \N__55515\
        );

    \I__13732\ : Span4Mux_h
    port map (
            O => \N__55550\,
            I => \N__55515\
        );

    \I__13731\ : LocalMux
    port map (
            O => \N__55547\,
            I => \N__55515\
        );

    \I__13730\ : Span4Mux_h
    port map (
            O => \N__55540\,
            I => \N__55515\
        );

    \I__13729\ : Odrv4
    port map (
            O => \N__55537\,
            I => dds_state_1
        );

    \I__13728\ : Odrv12
    port map (
            O => \N__55534\,
            I => dds_state_1
        );

    \I__13727\ : LocalMux
    port map (
            O => \N__55529\,
            I => dds_state_1
        );

    \I__13726\ : Odrv4
    port map (
            O => \N__55524\,
            I => dds_state_1
        );

    \I__13725\ : Odrv4
    port map (
            O => \N__55515\,
            I => dds_state_1
        );

    \I__13724\ : IoInMux
    port map (
            O => \N__55504\,
            I => \N__55501\
        );

    \I__13723\ : LocalMux
    port map (
            O => \N__55501\,
            I => \N__55498\
        );

    \I__13722\ : Span4Mux_s0_v
    port map (
            O => \N__55498\,
            I => \N__55495\
        );

    \I__13721\ : Span4Mux_h
    port map (
            O => \N__55495\,
            I => \N__55492\
        );

    \I__13720\ : Span4Mux_v
    port map (
            O => \N__55492\,
            I => \N__55489\
        );

    \I__13719\ : Span4Mux_v
    port map (
            O => \N__55489\,
            I => \N__55486\
        );

    \I__13718\ : Odrv4
    port map (
            O => \N__55486\,
            I => \DDS_CS\
        );

    \I__13717\ : CEMux
    port map (
            O => \N__55483\,
            I => \N__55480\
        );

    \I__13716\ : LocalMux
    port map (
            O => \N__55480\,
            I => \N__55477\
        );

    \I__13715\ : Odrv4
    port map (
            O => \N__55477\,
            I => \SIG_DDS.n9_adj_1385\
        );

    \I__13714\ : InMux
    port map (
            O => \N__55474\,
            I => \N__55469\
        );

    \I__13713\ : CascadeMux
    port map (
            O => \N__55473\,
            I => \N__55466\
        );

    \I__13712\ : InMux
    port map (
            O => \N__55472\,
            I => \N__55455\
        );

    \I__13711\ : LocalMux
    port map (
            O => \N__55469\,
            I => \N__55452\
        );

    \I__13710\ : InMux
    port map (
            O => \N__55466\,
            I => \N__55443\
        );

    \I__13709\ : InMux
    port map (
            O => \N__55465\,
            I => \N__55443\
        );

    \I__13708\ : InMux
    port map (
            O => \N__55464\,
            I => \N__55443\
        );

    \I__13707\ : InMux
    port map (
            O => \N__55463\,
            I => \N__55443\
        );

    \I__13706\ : InMux
    port map (
            O => \N__55462\,
            I => \N__55438\
        );

    \I__13705\ : InMux
    port map (
            O => \N__55461\,
            I => \N__55438\
        );

    \I__13704\ : InMux
    port map (
            O => \N__55460\,
            I => \N__55432\
        );

    \I__13703\ : InMux
    port map (
            O => \N__55459\,
            I => \N__55432\
        );

    \I__13702\ : InMux
    port map (
            O => \N__55458\,
            I => \N__55418\
        );

    \I__13701\ : LocalMux
    port map (
            O => \N__55455\,
            I => \N__55415\
        );

    \I__13700\ : Span4Mux_v
    port map (
            O => \N__55452\,
            I => \N__55410\
        );

    \I__13699\ : LocalMux
    port map (
            O => \N__55443\,
            I => \N__55410\
        );

    \I__13698\ : LocalMux
    port map (
            O => \N__55438\,
            I => \N__55398\
        );

    \I__13697\ : SRMux
    port map (
            O => \N__55437\,
            I => \N__55395\
        );

    \I__13696\ : LocalMux
    port map (
            O => \N__55432\,
            I => \N__55392\
        );

    \I__13695\ : SRMux
    port map (
            O => \N__55431\,
            I => \N__55389\
        );

    \I__13694\ : InMux
    port map (
            O => \N__55430\,
            I => \N__55384\
        );

    \I__13693\ : InMux
    port map (
            O => \N__55429\,
            I => \N__55384\
        );

    \I__13692\ : InMux
    port map (
            O => \N__55428\,
            I => \N__55379\
        );

    \I__13691\ : InMux
    port map (
            O => \N__55427\,
            I => \N__55362\
        );

    \I__13690\ : InMux
    port map (
            O => \N__55426\,
            I => \N__55362\
        );

    \I__13689\ : InMux
    port map (
            O => \N__55425\,
            I => \N__55362\
        );

    \I__13688\ : InMux
    port map (
            O => \N__55424\,
            I => \N__55362\
        );

    \I__13687\ : InMux
    port map (
            O => \N__55423\,
            I => \N__55362\
        );

    \I__13686\ : InMux
    port map (
            O => \N__55422\,
            I => \N__55362\
        );

    \I__13685\ : InMux
    port map (
            O => \N__55421\,
            I => \N__55362\
        );

    \I__13684\ : LocalMux
    port map (
            O => \N__55418\,
            I => \N__55355\
        );

    \I__13683\ : Span4Mux_h
    port map (
            O => \N__55415\,
            I => \N__55355\
        );

    \I__13682\ : Span4Mux_h
    port map (
            O => \N__55410\,
            I => \N__55355\
        );

    \I__13681\ : InMux
    port map (
            O => \N__55409\,
            I => \N__55350\
        );

    \I__13680\ : InMux
    port map (
            O => \N__55408\,
            I => \N__55350\
        );

    \I__13679\ : InMux
    port map (
            O => \N__55407\,
            I => \N__55347\
        );

    \I__13678\ : InMux
    port map (
            O => \N__55406\,
            I => \N__55342\
        );

    \I__13677\ : InMux
    port map (
            O => \N__55405\,
            I => \N__55342\
        );

    \I__13676\ : InMux
    port map (
            O => \N__55404\,
            I => \N__55333\
        );

    \I__13675\ : InMux
    port map (
            O => \N__55403\,
            I => \N__55333\
        );

    \I__13674\ : InMux
    port map (
            O => \N__55402\,
            I => \N__55333\
        );

    \I__13673\ : InMux
    port map (
            O => \N__55401\,
            I => \N__55333\
        );

    \I__13672\ : Span4Mux_v
    port map (
            O => \N__55398\,
            I => \N__55328\
        );

    \I__13671\ : LocalMux
    port map (
            O => \N__55395\,
            I => \N__55328\
        );

    \I__13670\ : Span4Mux_v
    port map (
            O => \N__55392\,
            I => \N__55321\
        );

    \I__13669\ : LocalMux
    port map (
            O => \N__55389\,
            I => \N__55321\
        );

    \I__13668\ : LocalMux
    port map (
            O => \N__55384\,
            I => \N__55321\
        );

    \I__13667\ : SRMux
    port map (
            O => \N__55383\,
            I => \N__55318\
        );

    \I__13666\ : InMux
    port map (
            O => \N__55382\,
            I => \N__55315\
        );

    \I__13665\ : LocalMux
    port map (
            O => \N__55379\,
            I => \N__55312\
        );

    \I__13664\ : InMux
    port map (
            O => \N__55378\,
            I => \N__55307\
        );

    \I__13663\ : InMux
    port map (
            O => \N__55377\,
            I => \N__55307\
        );

    \I__13662\ : LocalMux
    port map (
            O => \N__55362\,
            I => \N__55304\
        );

    \I__13661\ : Span4Mux_v
    port map (
            O => \N__55355\,
            I => \N__55299\
        );

    \I__13660\ : LocalMux
    port map (
            O => \N__55350\,
            I => \N__55299\
        );

    \I__13659\ : LocalMux
    port map (
            O => \N__55347\,
            I => \N__55294\
        );

    \I__13658\ : LocalMux
    port map (
            O => \N__55342\,
            I => \N__55294\
        );

    \I__13657\ : LocalMux
    port map (
            O => \N__55333\,
            I => \N__55291\
        );

    \I__13656\ : Span4Mux_h
    port map (
            O => \N__55328\,
            I => \N__55284\
        );

    \I__13655\ : Span4Mux_h
    port map (
            O => \N__55321\,
            I => \N__55284\
        );

    \I__13654\ : LocalMux
    port map (
            O => \N__55318\,
            I => \N__55284\
        );

    \I__13653\ : LocalMux
    port map (
            O => \N__55315\,
            I => \N__55281\
        );

    \I__13652\ : Span4Mux_v
    port map (
            O => \N__55312\,
            I => \N__55274\
        );

    \I__13651\ : LocalMux
    port map (
            O => \N__55307\,
            I => \N__55274\
        );

    \I__13650\ : Span4Mux_h
    port map (
            O => \N__55304\,
            I => \N__55274\
        );

    \I__13649\ : Span4Mux_h
    port map (
            O => \N__55299\,
            I => \N__55271\
        );

    \I__13648\ : Span4Mux_h
    port map (
            O => \N__55294\,
            I => \N__55268\
        );

    \I__13647\ : Span4Mux_v
    port map (
            O => \N__55291\,
            I => \N__55263\
        );

    \I__13646\ : Span4Mux_h
    port map (
            O => \N__55284\,
            I => \N__55263\
        );

    \I__13645\ : Span4Mux_h
    port map (
            O => \N__55281\,
            I => \N__55258\
        );

    \I__13644\ : Span4Mux_h
    port map (
            O => \N__55274\,
            I => \N__55258\
        );

    \I__13643\ : Span4Mux_h
    port map (
            O => \N__55271\,
            I => \N__55255\
        );

    \I__13642\ : Odrv4
    port map (
            O => \N__55268\,
            I => comm_clear
        );

    \I__13641\ : Odrv4
    port map (
            O => \N__55263\,
            I => comm_clear
        );

    \I__13640\ : Odrv4
    port map (
            O => \N__55258\,
            I => comm_clear
        );

    \I__13639\ : Odrv4
    port map (
            O => \N__55255\,
            I => comm_clear
        );

    \I__13638\ : ClkMux
    port map (
            O => \N__55246\,
            I => \N__54727\
        );

    \I__13637\ : ClkMux
    port map (
            O => \N__55245\,
            I => \N__54727\
        );

    \I__13636\ : ClkMux
    port map (
            O => \N__55244\,
            I => \N__54727\
        );

    \I__13635\ : ClkMux
    port map (
            O => \N__55243\,
            I => \N__54727\
        );

    \I__13634\ : ClkMux
    port map (
            O => \N__55242\,
            I => \N__54727\
        );

    \I__13633\ : ClkMux
    port map (
            O => \N__55241\,
            I => \N__54727\
        );

    \I__13632\ : ClkMux
    port map (
            O => \N__55240\,
            I => \N__54727\
        );

    \I__13631\ : ClkMux
    port map (
            O => \N__55239\,
            I => \N__54727\
        );

    \I__13630\ : ClkMux
    port map (
            O => \N__55238\,
            I => \N__54727\
        );

    \I__13629\ : ClkMux
    port map (
            O => \N__55237\,
            I => \N__54727\
        );

    \I__13628\ : ClkMux
    port map (
            O => \N__55236\,
            I => \N__54727\
        );

    \I__13627\ : ClkMux
    port map (
            O => \N__55235\,
            I => \N__54727\
        );

    \I__13626\ : ClkMux
    port map (
            O => \N__55234\,
            I => \N__54727\
        );

    \I__13625\ : ClkMux
    port map (
            O => \N__55233\,
            I => \N__54727\
        );

    \I__13624\ : ClkMux
    port map (
            O => \N__55232\,
            I => \N__54727\
        );

    \I__13623\ : ClkMux
    port map (
            O => \N__55231\,
            I => \N__54727\
        );

    \I__13622\ : ClkMux
    port map (
            O => \N__55230\,
            I => \N__54727\
        );

    \I__13621\ : ClkMux
    port map (
            O => \N__55229\,
            I => \N__54727\
        );

    \I__13620\ : ClkMux
    port map (
            O => \N__55228\,
            I => \N__54727\
        );

    \I__13619\ : ClkMux
    port map (
            O => \N__55227\,
            I => \N__54727\
        );

    \I__13618\ : ClkMux
    port map (
            O => \N__55226\,
            I => \N__54727\
        );

    \I__13617\ : ClkMux
    port map (
            O => \N__55225\,
            I => \N__54727\
        );

    \I__13616\ : ClkMux
    port map (
            O => \N__55224\,
            I => \N__54727\
        );

    \I__13615\ : ClkMux
    port map (
            O => \N__55223\,
            I => \N__54727\
        );

    \I__13614\ : ClkMux
    port map (
            O => \N__55222\,
            I => \N__54727\
        );

    \I__13613\ : ClkMux
    port map (
            O => \N__55221\,
            I => \N__54727\
        );

    \I__13612\ : ClkMux
    port map (
            O => \N__55220\,
            I => \N__54727\
        );

    \I__13611\ : ClkMux
    port map (
            O => \N__55219\,
            I => \N__54727\
        );

    \I__13610\ : ClkMux
    port map (
            O => \N__55218\,
            I => \N__54727\
        );

    \I__13609\ : ClkMux
    port map (
            O => \N__55217\,
            I => \N__54727\
        );

    \I__13608\ : ClkMux
    port map (
            O => \N__55216\,
            I => \N__54727\
        );

    \I__13607\ : ClkMux
    port map (
            O => \N__55215\,
            I => \N__54727\
        );

    \I__13606\ : ClkMux
    port map (
            O => \N__55214\,
            I => \N__54727\
        );

    \I__13605\ : ClkMux
    port map (
            O => \N__55213\,
            I => \N__54727\
        );

    \I__13604\ : ClkMux
    port map (
            O => \N__55212\,
            I => \N__54727\
        );

    \I__13603\ : ClkMux
    port map (
            O => \N__55211\,
            I => \N__54727\
        );

    \I__13602\ : ClkMux
    port map (
            O => \N__55210\,
            I => \N__54727\
        );

    \I__13601\ : ClkMux
    port map (
            O => \N__55209\,
            I => \N__54727\
        );

    \I__13600\ : ClkMux
    port map (
            O => \N__55208\,
            I => \N__54727\
        );

    \I__13599\ : ClkMux
    port map (
            O => \N__55207\,
            I => \N__54727\
        );

    \I__13598\ : ClkMux
    port map (
            O => \N__55206\,
            I => \N__54727\
        );

    \I__13597\ : ClkMux
    port map (
            O => \N__55205\,
            I => \N__54727\
        );

    \I__13596\ : ClkMux
    port map (
            O => \N__55204\,
            I => \N__54727\
        );

    \I__13595\ : ClkMux
    port map (
            O => \N__55203\,
            I => \N__54727\
        );

    \I__13594\ : ClkMux
    port map (
            O => \N__55202\,
            I => \N__54727\
        );

    \I__13593\ : ClkMux
    port map (
            O => \N__55201\,
            I => \N__54727\
        );

    \I__13592\ : ClkMux
    port map (
            O => \N__55200\,
            I => \N__54727\
        );

    \I__13591\ : ClkMux
    port map (
            O => \N__55199\,
            I => \N__54727\
        );

    \I__13590\ : ClkMux
    port map (
            O => \N__55198\,
            I => \N__54727\
        );

    \I__13589\ : ClkMux
    port map (
            O => \N__55197\,
            I => \N__54727\
        );

    \I__13588\ : ClkMux
    port map (
            O => \N__55196\,
            I => \N__54727\
        );

    \I__13587\ : ClkMux
    port map (
            O => \N__55195\,
            I => \N__54727\
        );

    \I__13586\ : ClkMux
    port map (
            O => \N__55194\,
            I => \N__54727\
        );

    \I__13585\ : ClkMux
    port map (
            O => \N__55193\,
            I => \N__54727\
        );

    \I__13584\ : ClkMux
    port map (
            O => \N__55192\,
            I => \N__54727\
        );

    \I__13583\ : ClkMux
    port map (
            O => \N__55191\,
            I => \N__54727\
        );

    \I__13582\ : ClkMux
    port map (
            O => \N__55190\,
            I => \N__54727\
        );

    \I__13581\ : ClkMux
    port map (
            O => \N__55189\,
            I => \N__54727\
        );

    \I__13580\ : ClkMux
    port map (
            O => \N__55188\,
            I => \N__54727\
        );

    \I__13579\ : ClkMux
    port map (
            O => \N__55187\,
            I => \N__54727\
        );

    \I__13578\ : ClkMux
    port map (
            O => \N__55186\,
            I => \N__54727\
        );

    \I__13577\ : ClkMux
    port map (
            O => \N__55185\,
            I => \N__54727\
        );

    \I__13576\ : ClkMux
    port map (
            O => \N__55184\,
            I => \N__54727\
        );

    \I__13575\ : ClkMux
    port map (
            O => \N__55183\,
            I => \N__54727\
        );

    \I__13574\ : ClkMux
    port map (
            O => \N__55182\,
            I => \N__54727\
        );

    \I__13573\ : ClkMux
    port map (
            O => \N__55181\,
            I => \N__54727\
        );

    \I__13572\ : ClkMux
    port map (
            O => \N__55180\,
            I => \N__54727\
        );

    \I__13571\ : ClkMux
    port map (
            O => \N__55179\,
            I => \N__54727\
        );

    \I__13570\ : ClkMux
    port map (
            O => \N__55178\,
            I => \N__54727\
        );

    \I__13569\ : ClkMux
    port map (
            O => \N__55177\,
            I => \N__54727\
        );

    \I__13568\ : ClkMux
    port map (
            O => \N__55176\,
            I => \N__54727\
        );

    \I__13567\ : ClkMux
    port map (
            O => \N__55175\,
            I => \N__54727\
        );

    \I__13566\ : ClkMux
    port map (
            O => \N__55174\,
            I => \N__54727\
        );

    \I__13565\ : ClkMux
    port map (
            O => \N__55173\,
            I => \N__54727\
        );

    \I__13564\ : ClkMux
    port map (
            O => \N__55172\,
            I => \N__54727\
        );

    \I__13563\ : ClkMux
    port map (
            O => \N__55171\,
            I => \N__54727\
        );

    \I__13562\ : ClkMux
    port map (
            O => \N__55170\,
            I => \N__54727\
        );

    \I__13561\ : ClkMux
    port map (
            O => \N__55169\,
            I => \N__54727\
        );

    \I__13560\ : ClkMux
    port map (
            O => \N__55168\,
            I => \N__54727\
        );

    \I__13559\ : ClkMux
    port map (
            O => \N__55167\,
            I => \N__54727\
        );

    \I__13558\ : ClkMux
    port map (
            O => \N__55166\,
            I => \N__54727\
        );

    \I__13557\ : ClkMux
    port map (
            O => \N__55165\,
            I => \N__54727\
        );

    \I__13556\ : ClkMux
    port map (
            O => \N__55164\,
            I => \N__54727\
        );

    \I__13555\ : ClkMux
    port map (
            O => \N__55163\,
            I => \N__54727\
        );

    \I__13554\ : ClkMux
    port map (
            O => \N__55162\,
            I => \N__54727\
        );

    \I__13553\ : ClkMux
    port map (
            O => \N__55161\,
            I => \N__54727\
        );

    \I__13552\ : ClkMux
    port map (
            O => \N__55160\,
            I => \N__54727\
        );

    \I__13551\ : ClkMux
    port map (
            O => \N__55159\,
            I => \N__54727\
        );

    \I__13550\ : ClkMux
    port map (
            O => \N__55158\,
            I => \N__54727\
        );

    \I__13549\ : ClkMux
    port map (
            O => \N__55157\,
            I => \N__54727\
        );

    \I__13548\ : ClkMux
    port map (
            O => \N__55156\,
            I => \N__54727\
        );

    \I__13547\ : ClkMux
    port map (
            O => \N__55155\,
            I => \N__54727\
        );

    \I__13546\ : ClkMux
    port map (
            O => \N__55154\,
            I => \N__54727\
        );

    \I__13545\ : ClkMux
    port map (
            O => \N__55153\,
            I => \N__54727\
        );

    \I__13544\ : ClkMux
    port map (
            O => \N__55152\,
            I => \N__54727\
        );

    \I__13543\ : ClkMux
    port map (
            O => \N__55151\,
            I => \N__54727\
        );

    \I__13542\ : ClkMux
    port map (
            O => \N__55150\,
            I => \N__54727\
        );

    \I__13541\ : ClkMux
    port map (
            O => \N__55149\,
            I => \N__54727\
        );

    \I__13540\ : ClkMux
    port map (
            O => \N__55148\,
            I => \N__54727\
        );

    \I__13539\ : ClkMux
    port map (
            O => \N__55147\,
            I => \N__54727\
        );

    \I__13538\ : ClkMux
    port map (
            O => \N__55146\,
            I => \N__54727\
        );

    \I__13537\ : ClkMux
    port map (
            O => \N__55145\,
            I => \N__54727\
        );

    \I__13536\ : ClkMux
    port map (
            O => \N__55144\,
            I => \N__54727\
        );

    \I__13535\ : ClkMux
    port map (
            O => \N__55143\,
            I => \N__54727\
        );

    \I__13534\ : ClkMux
    port map (
            O => \N__55142\,
            I => \N__54727\
        );

    \I__13533\ : ClkMux
    port map (
            O => \N__55141\,
            I => \N__54727\
        );

    \I__13532\ : ClkMux
    port map (
            O => \N__55140\,
            I => \N__54727\
        );

    \I__13531\ : ClkMux
    port map (
            O => \N__55139\,
            I => \N__54727\
        );

    \I__13530\ : ClkMux
    port map (
            O => \N__55138\,
            I => \N__54727\
        );

    \I__13529\ : ClkMux
    port map (
            O => \N__55137\,
            I => \N__54727\
        );

    \I__13528\ : ClkMux
    port map (
            O => \N__55136\,
            I => \N__54727\
        );

    \I__13527\ : ClkMux
    port map (
            O => \N__55135\,
            I => \N__54727\
        );

    \I__13526\ : ClkMux
    port map (
            O => \N__55134\,
            I => \N__54727\
        );

    \I__13525\ : ClkMux
    port map (
            O => \N__55133\,
            I => \N__54727\
        );

    \I__13524\ : ClkMux
    port map (
            O => \N__55132\,
            I => \N__54727\
        );

    \I__13523\ : ClkMux
    port map (
            O => \N__55131\,
            I => \N__54727\
        );

    \I__13522\ : ClkMux
    port map (
            O => \N__55130\,
            I => \N__54727\
        );

    \I__13521\ : ClkMux
    port map (
            O => \N__55129\,
            I => \N__54727\
        );

    \I__13520\ : ClkMux
    port map (
            O => \N__55128\,
            I => \N__54727\
        );

    \I__13519\ : ClkMux
    port map (
            O => \N__55127\,
            I => \N__54727\
        );

    \I__13518\ : ClkMux
    port map (
            O => \N__55126\,
            I => \N__54727\
        );

    \I__13517\ : ClkMux
    port map (
            O => \N__55125\,
            I => \N__54727\
        );

    \I__13516\ : ClkMux
    port map (
            O => \N__55124\,
            I => \N__54727\
        );

    \I__13515\ : ClkMux
    port map (
            O => \N__55123\,
            I => \N__54727\
        );

    \I__13514\ : ClkMux
    port map (
            O => \N__55122\,
            I => \N__54727\
        );

    \I__13513\ : ClkMux
    port map (
            O => \N__55121\,
            I => \N__54727\
        );

    \I__13512\ : ClkMux
    port map (
            O => \N__55120\,
            I => \N__54727\
        );

    \I__13511\ : ClkMux
    port map (
            O => \N__55119\,
            I => \N__54727\
        );

    \I__13510\ : ClkMux
    port map (
            O => \N__55118\,
            I => \N__54727\
        );

    \I__13509\ : ClkMux
    port map (
            O => \N__55117\,
            I => \N__54727\
        );

    \I__13508\ : ClkMux
    port map (
            O => \N__55116\,
            I => \N__54727\
        );

    \I__13507\ : ClkMux
    port map (
            O => \N__55115\,
            I => \N__54727\
        );

    \I__13506\ : ClkMux
    port map (
            O => \N__55114\,
            I => \N__54727\
        );

    \I__13505\ : ClkMux
    port map (
            O => \N__55113\,
            I => \N__54727\
        );

    \I__13504\ : ClkMux
    port map (
            O => \N__55112\,
            I => \N__54727\
        );

    \I__13503\ : ClkMux
    port map (
            O => \N__55111\,
            I => \N__54727\
        );

    \I__13502\ : ClkMux
    port map (
            O => \N__55110\,
            I => \N__54727\
        );

    \I__13501\ : ClkMux
    port map (
            O => \N__55109\,
            I => \N__54727\
        );

    \I__13500\ : ClkMux
    port map (
            O => \N__55108\,
            I => \N__54727\
        );

    \I__13499\ : ClkMux
    port map (
            O => \N__55107\,
            I => \N__54727\
        );

    \I__13498\ : ClkMux
    port map (
            O => \N__55106\,
            I => \N__54727\
        );

    \I__13497\ : ClkMux
    port map (
            O => \N__55105\,
            I => \N__54727\
        );

    \I__13496\ : ClkMux
    port map (
            O => \N__55104\,
            I => \N__54727\
        );

    \I__13495\ : ClkMux
    port map (
            O => \N__55103\,
            I => \N__54727\
        );

    \I__13494\ : ClkMux
    port map (
            O => \N__55102\,
            I => \N__54727\
        );

    \I__13493\ : ClkMux
    port map (
            O => \N__55101\,
            I => \N__54727\
        );

    \I__13492\ : ClkMux
    port map (
            O => \N__55100\,
            I => \N__54727\
        );

    \I__13491\ : ClkMux
    port map (
            O => \N__55099\,
            I => \N__54727\
        );

    \I__13490\ : ClkMux
    port map (
            O => \N__55098\,
            I => \N__54727\
        );

    \I__13489\ : ClkMux
    port map (
            O => \N__55097\,
            I => \N__54727\
        );

    \I__13488\ : ClkMux
    port map (
            O => \N__55096\,
            I => \N__54727\
        );

    \I__13487\ : ClkMux
    port map (
            O => \N__55095\,
            I => \N__54727\
        );

    \I__13486\ : ClkMux
    port map (
            O => \N__55094\,
            I => \N__54727\
        );

    \I__13485\ : ClkMux
    port map (
            O => \N__55093\,
            I => \N__54727\
        );

    \I__13484\ : ClkMux
    port map (
            O => \N__55092\,
            I => \N__54727\
        );

    \I__13483\ : ClkMux
    port map (
            O => \N__55091\,
            I => \N__54727\
        );

    \I__13482\ : ClkMux
    port map (
            O => \N__55090\,
            I => \N__54727\
        );

    \I__13481\ : ClkMux
    port map (
            O => \N__55089\,
            I => \N__54727\
        );

    \I__13480\ : ClkMux
    port map (
            O => \N__55088\,
            I => \N__54727\
        );

    \I__13479\ : ClkMux
    port map (
            O => \N__55087\,
            I => \N__54727\
        );

    \I__13478\ : ClkMux
    port map (
            O => \N__55086\,
            I => \N__54727\
        );

    \I__13477\ : ClkMux
    port map (
            O => \N__55085\,
            I => \N__54727\
        );

    \I__13476\ : ClkMux
    port map (
            O => \N__55084\,
            I => \N__54727\
        );

    \I__13475\ : ClkMux
    port map (
            O => \N__55083\,
            I => \N__54727\
        );

    \I__13474\ : ClkMux
    port map (
            O => \N__55082\,
            I => \N__54727\
        );

    \I__13473\ : ClkMux
    port map (
            O => \N__55081\,
            I => \N__54727\
        );

    \I__13472\ : ClkMux
    port map (
            O => \N__55080\,
            I => \N__54727\
        );

    \I__13471\ : ClkMux
    port map (
            O => \N__55079\,
            I => \N__54727\
        );

    \I__13470\ : ClkMux
    port map (
            O => \N__55078\,
            I => \N__54727\
        );

    \I__13469\ : ClkMux
    port map (
            O => \N__55077\,
            I => \N__54727\
        );

    \I__13468\ : ClkMux
    port map (
            O => \N__55076\,
            I => \N__54727\
        );

    \I__13467\ : ClkMux
    port map (
            O => \N__55075\,
            I => \N__54727\
        );

    \I__13466\ : ClkMux
    port map (
            O => \N__55074\,
            I => \N__54727\
        );

    \I__13465\ : GlobalMux
    port map (
            O => \N__54727\,
            I => \clk_32MHz\
        );

    \I__13464\ : InMux
    port map (
            O => \N__54724\,
            I => \N__54706\
        );

    \I__13463\ : InMux
    port map (
            O => \N__54723\,
            I => \N__54696\
        );

    \I__13462\ : InMux
    port map (
            O => \N__54722\,
            I => \N__54690\
        );

    \I__13461\ : InMux
    port map (
            O => \N__54721\,
            I => \N__54687\
        );

    \I__13460\ : InMux
    port map (
            O => \N__54720\,
            I => \N__54684\
        );

    \I__13459\ : InMux
    port map (
            O => \N__54719\,
            I => \N__54681\
        );

    \I__13458\ : InMux
    port map (
            O => \N__54718\,
            I => \N__54676\
        );

    \I__13457\ : InMux
    port map (
            O => \N__54717\,
            I => \N__54676\
        );

    \I__13456\ : CascadeMux
    port map (
            O => \N__54716\,
            I => \N__54653\
        );

    \I__13455\ : CascadeMux
    port map (
            O => \N__54715\,
            I => \N__54650\
        );

    \I__13454\ : CascadeMux
    port map (
            O => \N__54714\,
            I => \N__54646\
        );

    \I__13453\ : CascadeMux
    port map (
            O => \N__54713\,
            I => \N__54642\
        );

    \I__13452\ : CascadeMux
    port map (
            O => \N__54712\,
            I => \N__54639\
        );

    \I__13451\ : CascadeMux
    port map (
            O => \N__54711\,
            I => \N__54636\
        );

    \I__13450\ : InMux
    port map (
            O => \N__54710\,
            I => \N__54632\
        );

    \I__13449\ : InMux
    port map (
            O => \N__54709\,
            I => \N__54629\
        );

    \I__13448\ : LocalMux
    port map (
            O => \N__54706\,
            I => \N__54626\
        );

    \I__13447\ : InMux
    port map (
            O => \N__54705\,
            I => \N__54620\
        );

    \I__13446\ : InMux
    port map (
            O => \N__54704\,
            I => \N__54617\
        );

    \I__13445\ : InMux
    port map (
            O => \N__54703\,
            I => \N__54612\
        );

    \I__13444\ : InMux
    port map (
            O => \N__54702\,
            I => \N__54612\
        );

    \I__13443\ : InMux
    port map (
            O => \N__54701\,
            I => \N__54604\
        );

    \I__13442\ : InMux
    port map (
            O => \N__54700\,
            I => \N__54604\
        );

    \I__13441\ : InMux
    port map (
            O => \N__54699\,
            I => \N__54601\
        );

    \I__13440\ : LocalMux
    port map (
            O => \N__54696\,
            I => \N__54593\
        );

    \I__13439\ : CascadeMux
    port map (
            O => \N__54695\,
            I => \N__54585\
        );

    \I__13438\ : CascadeMux
    port map (
            O => \N__54694\,
            I => \N__54581\
        );

    \I__13437\ : CascadeMux
    port map (
            O => \N__54693\,
            I => \N__54577\
        );

    \I__13436\ : LocalMux
    port map (
            O => \N__54690\,
            I => \N__54571\
        );

    \I__13435\ : LocalMux
    port map (
            O => \N__54687\,
            I => \N__54571\
        );

    \I__13434\ : LocalMux
    port map (
            O => \N__54684\,
            I => \N__54564\
        );

    \I__13433\ : LocalMux
    port map (
            O => \N__54681\,
            I => \N__54564\
        );

    \I__13432\ : LocalMux
    port map (
            O => \N__54676\,
            I => \N__54564\
        );

    \I__13431\ : InMux
    port map (
            O => \N__54675\,
            I => \N__54558\
        );

    \I__13430\ : InMux
    port map (
            O => \N__54674\,
            I => \N__54555\
        );

    \I__13429\ : InMux
    port map (
            O => \N__54673\,
            I => \N__54550\
        );

    \I__13428\ : InMux
    port map (
            O => \N__54672\,
            I => \N__54550\
        );

    \I__13427\ : InMux
    port map (
            O => \N__54671\,
            I => \N__54545\
        );

    \I__13426\ : InMux
    port map (
            O => \N__54670\,
            I => \N__54545\
        );

    \I__13425\ : CascadeMux
    port map (
            O => \N__54669\,
            I => \N__54541\
        );

    \I__13424\ : InMux
    port map (
            O => \N__54668\,
            I => \N__54538\
        );

    \I__13423\ : InMux
    port map (
            O => \N__54667\,
            I => \N__54522\
        );

    \I__13422\ : InMux
    port map (
            O => \N__54666\,
            I => \N__54522\
        );

    \I__13421\ : InMux
    port map (
            O => \N__54665\,
            I => \N__54522\
        );

    \I__13420\ : InMux
    port map (
            O => \N__54664\,
            I => \N__54522\
        );

    \I__13419\ : InMux
    port map (
            O => \N__54663\,
            I => \N__54522\
        );

    \I__13418\ : InMux
    port map (
            O => \N__54662\,
            I => \N__54522\
        );

    \I__13417\ : InMux
    port map (
            O => \N__54661\,
            I => \N__54511\
        );

    \I__13416\ : InMux
    port map (
            O => \N__54660\,
            I => \N__54511\
        );

    \I__13415\ : InMux
    port map (
            O => \N__54659\,
            I => \N__54511\
        );

    \I__13414\ : InMux
    port map (
            O => \N__54658\,
            I => \N__54511\
        );

    \I__13413\ : InMux
    port map (
            O => \N__54657\,
            I => \N__54511\
        );

    \I__13412\ : InMux
    port map (
            O => \N__54656\,
            I => \N__54508\
        );

    \I__13411\ : InMux
    port map (
            O => \N__54653\,
            I => \N__54495\
        );

    \I__13410\ : InMux
    port map (
            O => \N__54650\,
            I => \N__54495\
        );

    \I__13409\ : InMux
    port map (
            O => \N__54649\,
            I => \N__54495\
        );

    \I__13408\ : InMux
    port map (
            O => \N__54646\,
            I => \N__54495\
        );

    \I__13407\ : InMux
    port map (
            O => \N__54645\,
            I => \N__54495\
        );

    \I__13406\ : InMux
    port map (
            O => \N__54642\,
            I => \N__54495\
        );

    \I__13405\ : InMux
    port map (
            O => \N__54639\,
            I => \N__54490\
        );

    \I__13404\ : InMux
    port map (
            O => \N__54636\,
            I => \N__54490\
        );

    \I__13403\ : InMux
    port map (
            O => \N__54635\,
            I => \N__54482\
        );

    \I__13402\ : LocalMux
    port map (
            O => \N__54632\,
            I => \N__54475\
        );

    \I__13401\ : LocalMux
    port map (
            O => \N__54629\,
            I => \N__54475\
        );

    \I__13400\ : Span4Mux_h
    port map (
            O => \N__54626\,
            I => \N__54475\
        );

    \I__13399\ : InMux
    port map (
            O => \N__54625\,
            I => \N__54472\
        );

    \I__13398\ : InMux
    port map (
            O => \N__54624\,
            I => \N__54467\
        );

    \I__13397\ : InMux
    port map (
            O => \N__54623\,
            I => \N__54467\
        );

    \I__13396\ : LocalMux
    port map (
            O => \N__54620\,
            I => \N__54460\
        );

    \I__13395\ : LocalMux
    port map (
            O => \N__54617\,
            I => \N__54460\
        );

    \I__13394\ : LocalMux
    port map (
            O => \N__54612\,
            I => \N__54460\
        );

    \I__13393\ : InMux
    port map (
            O => \N__54611\,
            I => \N__54455\
        );

    \I__13392\ : InMux
    port map (
            O => \N__54610\,
            I => \N__54455\
        );

    \I__13391\ : SRMux
    port map (
            O => \N__54609\,
            I => \N__54452\
        );

    \I__13390\ : LocalMux
    port map (
            O => \N__54604\,
            I => \N__54448\
        );

    \I__13389\ : LocalMux
    port map (
            O => \N__54601\,
            I => \N__54445\
        );

    \I__13388\ : InMux
    port map (
            O => \N__54600\,
            I => \N__54442\
        );

    \I__13387\ : CascadeMux
    port map (
            O => \N__54599\,
            I => \N__54437\
        );

    \I__13386\ : CascadeMux
    port map (
            O => \N__54598\,
            I => \N__54434\
        );

    \I__13385\ : InMux
    port map (
            O => \N__54597\,
            I => \N__54430\
        );

    \I__13384\ : InMux
    port map (
            O => \N__54596\,
            I => \N__54427\
        );

    \I__13383\ : Span4Mux_h
    port map (
            O => \N__54593\,
            I => \N__54424\
        );

    \I__13382\ : InMux
    port map (
            O => \N__54592\,
            I => \N__54421\
        );

    \I__13381\ : InMux
    port map (
            O => \N__54591\,
            I => \N__54416\
        );

    \I__13380\ : InMux
    port map (
            O => \N__54590\,
            I => \N__54416\
        );

    \I__13379\ : InMux
    port map (
            O => \N__54589\,
            I => \N__54399\
        );

    \I__13378\ : InMux
    port map (
            O => \N__54588\,
            I => \N__54399\
        );

    \I__13377\ : InMux
    port map (
            O => \N__54585\,
            I => \N__54399\
        );

    \I__13376\ : InMux
    port map (
            O => \N__54584\,
            I => \N__54399\
        );

    \I__13375\ : InMux
    port map (
            O => \N__54581\,
            I => \N__54399\
        );

    \I__13374\ : InMux
    port map (
            O => \N__54580\,
            I => \N__54399\
        );

    \I__13373\ : InMux
    port map (
            O => \N__54577\,
            I => \N__54399\
        );

    \I__13372\ : InMux
    port map (
            O => \N__54576\,
            I => \N__54399\
        );

    \I__13371\ : Span4Mux_v
    port map (
            O => \N__54571\,
            I => \N__54394\
        );

    \I__13370\ : Span4Mux_v
    port map (
            O => \N__54564\,
            I => \N__54394\
        );

    \I__13369\ : InMux
    port map (
            O => \N__54563\,
            I => \N__54389\
        );

    \I__13368\ : InMux
    port map (
            O => \N__54562\,
            I => \N__54389\
        );

    \I__13367\ : InMux
    port map (
            O => \N__54561\,
            I => \N__54384\
        );

    \I__13366\ : LocalMux
    port map (
            O => \N__54558\,
            I => \N__54381\
        );

    \I__13365\ : LocalMux
    port map (
            O => \N__54555\,
            I => \N__54376\
        );

    \I__13364\ : LocalMux
    port map (
            O => \N__54550\,
            I => \N__54376\
        );

    \I__13363\ : LocalMux
    port map (
            O => \N__54545\,
            I => \N__54373\
        );

    \I__13362\ : InMux
    port map (
            O => \N__54544\,
            I => \N__54369\
        );

    \I__13361\ : InMux
    port map (
            O => \N__54541\,
            I => \N__54364\
        );

    \I__13360\ : LocalMux
    port map (
            O => \N__54538\,
            I => \N__54361\
        );

    \I__13359\ : InMux
    port map (
            O => \N__54537\,
            I => \N__54358\
        );

    \I__13358\ : InMux
    port map (
            O => \N__54536\,
            I => \N__54355\
        );

    \I__13357\ : InMux
    port map (
            O => \N__54535\,
            I => \N__54352\
        );

    \I__13356\ : LocalMux
    port map (
            O => \N__54522\,
            I => \N__54341\
        );

    \I__13355\ : LocalMux
    port map (
            O => \N__54511\,
            I => \N__54341\
        );

    \I__13354\ : LocalMux
    port map (
            O => \N__54508\,
            I => \N__54341\
        );

    \I__13353\ : LocalMux
    port map (
            O => \N__54495\,
            I => \N__54341\
        );

    \I__13352\ : LocalMux
    port map (
            O => \N__54490\,
            I => \N__54341\
        );

    \I__13351\ : InMux
    port map (
            O => \N__54489\,
            I => \N__54336\
        );

    \I__13350\ : InMux
    port map (
            O => \N__54488\,
            I => \N__54336\
        );

    \I__13349\ : InMux
    port map (
            O => \N__54487\,
            I => \N__54329\
        );

    \I__13348\ : InMux
    port map (
            O => \N__54486\,
            I => \N__54329\
        );

    \I__13347\ : InMux
    port map (
            O => \N__54485\,
            I => \N__54329\
        );

    \I__13346\ : LocalMux
    port map (
            O => \N__54482\,
            I => \N__54318\
        );

    \I__13345\ : Span4Mux_h
    port map (
            O => \N__54475\,
            I => \N__54318\
        );

    \I__13344\ : LocalMux
    port map (
            O => \N__54472\,
            I => \N__54318\
        );

    \I__13343\ : LocalMux
    port map (
            O => \N__54467\,
            I => \N__54318\
        );

    \I__13342\ : Span4Mux_v
    port map (
            O => \N__54460\,
            I => \N__54318\
        );

    \I__13341\ : LocalMux
    port map (
            O => \N__54455\,
            I => \N__54315\
        );

    \I__13340\ : LocalMux
    port map (
            O => \N__54452\,
            I => \N__54312\
        );

    \I__13339\ : InMux
    port map (
            O => \N__54451\,
            I => \N__54309\
        );

    \I__13338\ : Span4Mux_h
    port map (
            O => \N__54448\,
            I => \N__54306\
        );

    \I__13337\ : Span4Mux_h
    port map (
            O => \N__54445\,
            I => \N__54301\
        );

    \I__13336\ : LocalMux
    port map (
            O => \N__54442\,
            I => \N__54301\
        );

    \I__13335\ : InMux
    port map (
            O => \N__54441\,
            I => \N__54298\
        );

    \I__13334\ : InMux
    port map (
            O => \N__54440\,
            I => \N__54295\
        );

    \I__13333\ : InMux
    port map (
            O => \N__54437\,
            I => \N__54288\
        );

    \I__13332\ : InMux
    port map (
            O => \N__54434\,
            I => \N__54288\
        );

    \I__13331\ : InMux
    port map (
            O => \N__54433\,
            I => \N__54288\
        );

    \I__13330\ : LocalMux
    port map (
            O => \N__54430\,
            I => \N__54285\
        );

    \I__13329\ : LocalMux
    port map (
            O => \N__54427\,
            I => \N__54280\
        );

    \I__13328\ : Span4Mux_h
    port map (
            O => \N__54424\,
            I => \N__54280\
        );

    \I__13327\ : LocalMux
    port map (
            O => \N__54421\,
            I => \N__54275\
        );

    \I__13326\ : LocalMux
    port map (
            O => \N__54416\,
            I => \N__54275\
        );

    \I__13325\ : LocalMux
    port map (
            O => \N__54399\,
            I => \N__54268\
        );

    \I__13324\ : Span4Mux_h
    port map (
            O => \N__54394\,
            I => \N__54268\
        );

    \I__13323\ : LocalMux
    port map (
            O => \N__54389\,
            I => \N__54268\
        );

    \I__13322\ : InMux
    port map (
            O => \N__54388\,
            I => \N__54263\
        );

    \I__13321\ : InMux
    port map (
            O => \N__54387\,
            I => \N__54263\
        );

    \I__13320\ : LocalMux
    port map (
            O => \N__54384\,
            I => \N__54260\
        );

    \I__13319\ : Span4Mux_v
    port map (
            O => \N__54381\,
            I => \N__54253\
        );

    \I__13318\ : Span4Mux_h
    port map (
            O => \N__54376\,
            I => \N__54253\
        );

    \I__13317\ : Span4Mux_v
    port map (
            O => \N__54373\,
            I => \N__54253\
        );

    \I__13316\ : InMux
    port map (
            O => \N__54372\,
            I => \N__54250\
        );

    \I__13315\ : LocalMux
    port map (
            O => \N__54369\,
            I => \N__54246\
        );

    \I__13314\ : CascadeMux
    port map (
            O => \N__54368\,
            I => \N__54241\
        );

    \I__13313\ : InMux
    port map (
            O => \N__54367\,
            I => \N__54235\
        );

    \I__13312\ : LocalMux
    port map (
            O => \N__54364\,
            I => \N__54228\
        );

    \I__13311\ : Span4Mux_v
    port map (
            O => \N__54361\,
            I => \N__54228\
        );

    \I__13310\ : LocalMux
    port map (
            O => \N__54358\,
            I => \N__54228\
        );

    \I__13309\ : LocalMux
    port map (
            O => \N__54355\,
            I => \N__54223\
        );

    \I__13308\ : LocalMux
    port map (
            O => \N__54352\,
            I => \N__54223\
        );

    \I__13307\ : Span4Mux_v
    port map (
            O => \N__54341\,
            I => \N__54220\
        );

    \I__13306\ : LocalMux
    port map (
            O => \N__54336\,
            I => \N__54211\
        );

    \I__13305\ : LocalMux
    port map (
            O => \N__54329\,
            I => \N__54211\
        );

    \I__13304\ : Span4Mux_v
    port map (
            O => \N__54318\,
            I => \N__54211\
        );

    \I__13303\ : Span4Mux_v
    port map (
            O => \N__54315\,
            I => \N__54211\
        );

    \I__13302\ : Span4Mux_v
    port map (
            O => \N__54312\,
            I => \N__54200\
        );

    \I__13301\ : LocalMux
    port map (
            O => \N__54309\,
            I => \N__54200\
        );

    \I__13300\ : Span4Mux_h
    port map (
            O => \N__54306\,
            I => \N__54200\
        );

    \I__13299\ : Span4Mux_h
    port map (
            O => \N__54301\,
            I => \N__54200\
        );

    \I__13298\ : LocalMux
    port map (
            O => \N__54298\,
            I => \N__54200\
        );

    \I__13297\ : LocalMux
    port map (
            O => \N__54295\,
            I => \N__54193\
        );

    \I__13296\ : LocalMux
    port map (
            O => \N__54288\,
            I => \N__54193\
        );

    \I__13295\ : Span4Mux_h
    port map (
            O => \N__54285\,
            I => \N__54193\
        );

    \I__13294\ : Sp12to4
    port map (
            O => \N__54280\,
            I => \N__54184\
        );

    \I__13293\ : Sp12to4
    port map (
            O => \N__54275\,
            I => \N__54184\
        );

    \I__13292\ : Sp12to4
    port map (
            O => \N__54268\,
            I => \N__54184\
        );

    \I__13291\ : LocalMux
    port map (
            O => \N__54263\,
            I => \N__54184\
        );

    \I__13290\ : Span4Mux_h
    port map (
            O => \N__54260\,
            I => \N__54177\
        );

    \I__13289\ : Span4Mux_v
    port map (
            O => \N__54253\,
            I => \N__54177\
        );

    \I__13288\ : LocalMux
    port map (
            O => \N__54250\,
            I => \N__54177\
        );

    \I__13287\ : InMux
    port map (
            O => \N__54249\,
            I => \N__54172\
        );

    \I__13286\ : Span4Mux_h
    port map (
            O => \N__54246\,
            I => \N__54169\
        );

    \I__13285\ : InMux
    port map (
            O => \N__54245\,
            I => \N__54166\
        );

    \I__13284\ : InMux
    port map (
            O => \N__54244\,
            I => \N__54157\
        );

    \I__13283\ : InMux
    port map (
            O => \N__54241\,
            I => \N__54157\
        );

    \I__13282\ : InMux
    port map (
            O => \N__54240\,
            I => \N__54157\
        );

    \I__13281\ : InMux
    port map (
            O => \N__54239\,
            I => \N__54157\
        );

    \I__13280\ : InMux
    port map (
            O => \N__54238\,
            I => \N__54154\
        );

    \I__13279\ : LocalMux
    port map (
            O => \N__54235\,
            I => \N__54143\
        );

    \I__13278\ : Span4Mux_v
    port map (
            O => \N__54228\,
            I => \N__54143\
        );

    \I__13277\ : Span4Mux_v
    port map (
            O => \N__54223\,
            I => \N__54143\
        );

    \I__13276\ : Span4Mux_h
    port map (
            O => \N__54220\,
            I => \N__54143\
        );

    \I__13275\ : Span4Mux_v
    port map (
            O => \N__54211\,
            I => \N__54143\
        );

    \I__13274\ : Sp12to4
    port map (
            O => \N__54200\,
            I => \N__54138\
        );

    \I__13273\ : Sp12to4
    port map (
            O => \N__54193\,
            I => \N__54138\
        );

    \I__13272\ : Span12Mux_v
    port map (
            O => \N__54184\,
            I => \N__54135\
        );

    \I__13271\ : Span4Mux_h
    port map (
            O => \N__54177\,
            I => \N__54132\
        );

    \I__13270\ : InMux
    port map (
            O => \N__54176\,
            I => \N__54127\
        );

    \I__13269\ : InMux
    port map (
            O => \N__54175\,
            I => \N__54127\
        );

    \I__13268\ : LocalMux
    port map (
            O => \N__54172\,
            I => comm_state_3
        );

    \I__13267\ : Odrv4
    port map (
            O => \N__54169\,
            I => comm_state_3
        );

    \I__13266\ : LocalMux
    port map (
            O => \N__54166\,
            I => comm_state_3
        );

    \I__13265\ : LocalMux
    port map (
            O => \N__54157\,
            I => comm_state_3
        );

    \I__13264\ : LocalMux
    port map (
            O => \N__54154\,
            I => comm_state_3
        );

    \I__13263\ : Odrv4
    port map (
            O => \N__54143\,
            I => comm_state_3
        );

    \I__13262\ : Odrv12
    port map (
            O => \N__54138\,
            I => comm_state_3
        );

    \I__13261\ : Odrv12
    port map (
            O => \N__54135\,
            I => comm_state_3
        );

    \I__13260\ : Odrv4
    port map (
            O => \N__54132\,
            I => comm_state_3
        );

    \I__13259\ : LocalMux
    port map (
            O => \N__54127\,
            I => comm_state_3
        );

    \I__13258\ : InMux
    port map (
            O => \N__54106\,
            I => \N__54076\
        );

    \I__13257\ : InMux
    port map (
            O => \N__54105\,
            I => \N__54067\
        );

    \I__13256\ : InMux
    port map (
            O => \N__54104\,
            I => \N__54067\
        );

    \I__13255\ : InMux
    port map (
            O => \N__54103\,
            I => \N__54067\
        );

    \I__13254\ : InMux
    port map (
            O => \N__54102\,
            I => \N__54067\
        );

    \I__13253\ : InMux
    port map (
            O => \N__54101\,
            I => \N__54064\
        );

    \I__13252\ : InMux
    port map (
            O => \N__54100\,
            I => \N__54061\
        );

    \I__13251\ : InMux
    port map (
            O => \N__54099\,
            I => \N__54052\
        );

    \I__13250\ : InMux
    port map (
            O => \N__54098\,
            I => \N__54052\
        );

    \I__13249\ : InMux
    port map (
            O => \N__54097\,
            I => \N__54052\
        );

    \I__13248\ : InMux
    port map (
            O => \N__54096\,
            I => \N__54052\
        );

    \I__13247\ : InMux
    port map (
            O => \N__54095\,
            I => \N__54048\
        );

    \I__13246\ : InMux
    port map (
            O => \N__54094\,
            I => \N__54045\
        );

    \I__13245\ : InMux
    port map (
            O => \N__54093\,
            I => \N__54042\
        );

    \I__13244\ : InMux
    port map (
            O => \N__54092\,
            I => \N__54039\
        );

    \I__13243\ : InMux
    port map (
            O => \N__54091\,
            I => \N__54036\
        );

    \I__13242\ : InMux
    port map (
            O => \N__54090\,
            I => \N__54028\
        );

    \I__13241\ : InMux
    port map (
            O => \N__54089\,
            I => \N__54010\
        );

    \I__13240\ : InMux
    port map (
            O => \N__54088\,
            I => \N__54010\
        );

    \I__13239\ : InMux
    port map (
            O => \N__54087\,
            I => \N__54010\
        );

    \I__13238\ : InMux
    port map (
            O => \N__54086\,
            I => \N__54010\
        );

    \I__13237\ : InMux
    port map (
            O => \N__54085\,
            I => \N__54010\
        );

    \I__13236\ : InMux
    port map (
            O => \N__54084\,
            I => \N__54010\
        );

    \I__13235\ : InMux
    port map (
            O => \N__54083\,
            I => \N__54010\
        );

    \I__13234\ : InMux
    port map (
            O => \N__54082\,
            I => \N__54010\
        );

    \I__13233\ : InMux
    port map (
            O => \N__54081\,
            I => \N__54005\
        );

    \I__13232\ : InMux
    port map (
            O => \N__54080\,
            I => \N__54005\
        );

    \I__13231\ : InMux
    port map (
            O => \N__54079\,
            I => \N__54002\
        );

    \I__13230\ : LocalMux
    port map (
            O => \N__54076\,
            I => \N__53997\
        );

    \I__13229\ : LocalMux
    port map (
            O => \N__54067\,
            I => \N__53988\
        );

    \I__13228\ : LocalMux
    port map (
            O => \N__54064\,
            I => \N__53988\
        );

    \I__13227\ : LocalMux
    port map (
            O => \N__54061\,
            I => \N__53988\
        );

    \I__13226\ : LocalMux
    port map (
            O => \N__54052\,
            I => \N__53988\
        );

    \I__13225\ : InMux
    port map (
            O => \N__54051\,
            I => \N__53972\
        );

    \I__13224\ : LocalMux
    port map (
            O => \N__54048\,
            I => \N__53967\
        );

    \I__13223\ : LocalMux
    port map (
            O => \N__54045\,
            I => \N__53967\
        );

    \I__13222\ : LocalMux
    port map (
            O => \N__54042\,
            I => \N__53964\
        );

    \I__13221\ : LocalMux
    port map (
            O => \N__54039\,
            I => \N__53961\
        );

    \I__13220\ : LocalMux
    port map (
            O => \N__54036\,
            I => \N__53958\
        );

    \I__13219\ : InMux
    port map (
            O => \N__54035\,
            I => \N__53953\
        );

    \I__13218\ : InMux
    port map (
            O => \N__54034\,
            I => \N__53950\
        );

    \I__13217\ : InMux
    port map (
            O => \N__54033\,
            I => \N__53932\
        );

    \I__13216\ : InMux
    port map (
            O => \N__54032\,
            I => \N__53929\
        );

    \I__13215\ : InMux
    port map (
            O => \N__54031\,
            I => \N__53926\
        );

    \I__13214\ : LocalMux
    port map (
            O => \N__54028\,
            I => \N__53923\
        );

    \I__13213\ : InMux
    port map (
            O => \N__54027\,
            I => \N__53920\
        );

    \I__13212\ : LocalMux
    port map (
            O => \N__54010\,
            I => \N__53913\
        );

    \I__13211\ : LocalMux
    port map (
            O => \N__54005\,
            I => \N__53913\
        );

    \I__13210\ : LocalMux
    port map (
            O => \N__54002\,
            I => \N__53913\
        );

    \I__13209\ : CascadeMux
    port map (
            O => \N__54001\,
            I => \N__53910\
        );

    \I__13208\ : InMux
    port map (
            O => \N__54000\,
            I => \N__53905\
        );

    \I__13207\ : Span4Mux_v
    port map (
            O => \N__53997\,
            I => \N__53895\
        );

    \I__13206\ : Span4Mux_v
    port map (
            O => \N__53988\,
            I => \N__53895\
        );

    \I__13205\ : InMux
    port map (
            O => \N__53987\,
            I => \N__53892\
        );

    \I__13204\ : InMux
    port map (
            O => \N__53986\,
            I => \N__53889\
        );

    \I__13203\ : InMux
    port map (
            O => \N__53985\,
            I => \N__53886\
        );

    \I__13202\ : InMux
    port map (
            O => \N__53984\,
            I => \N__53878\
        );

    \I__13201\ : InMux
    port map (
            O => \N__53983\,
            I => \N__53875\
        );

    \I__13200\ : InMux
    port map (
            O => \N__53982\,
            I => \N__53854\
        );

    \I__13199\ : InMux
    port map (
            O => \N__53981\,
            I => \N__53854\
        );

    \I__13198\ : InMux
    port map (
            O => \N__53980\,
            I => \N__53854\
        );

    \I__13197\ : InMux
    port map (
            O => \N__53979\,
            I => \N__53854\
        );

    \I__13196\ : InMux
    port map (
            O => \N__53978\,
            I => \N__53854\
        );

    \I__13195\ : InMux
    port map (
            O => \N__53977\,
            I => \N__53854\
        );

    \I__13194\ : InMux
    port map (
            O => \N__53976\,
            I => \N__53854\
        );

    \I__13193\ : InMux
    port map (
            O => \N__53975\,
            I => \N__53854\
        );

    \I__13192\ : LocalMux
    port map (
            O => \N__53972\,
            I => \N__53851\
        );

    \I__13191\ : Span4Mux_v
    port map (
            O => \N__53967\,
            I => \N__53848\
        );

    \I__13190\ : Span4Mux_v
    port map (
            O => \N__53964\,
            I => \N__53843\
        );

    \I__13189\ : Span4Mux_v
    port map (
            O => \N__53961\,
            I => \N__53843\
        );

    \I__13188\ : Span4Mux_v
    port map (
            O => \N__53958\,
            I => \N__53840\
        );

    \I__13187\ : InMux
    port map (
            O => \N__53957\,
            I => \N__53834\
        );

    \I__13186\ : InMux
    port map (
            O => \N__53956\,
            I => \N__53831\
        );

    \I__13185\ : LocalMux
    port map (
            O => \N__53953\,
            I => \N__53823\
        );

    \I__13184\ : LocalMux
    port map (
            O => \N__53950\,
            I => \N__53823\
        );

    \I__13183\ : InMux
    port map (
            O => \N__53949\,
            I => \N__53806\
        );

    \I__13182\ : InMux
    port map (
            O => \N__53948\,
            I => \N__53806\
        );

    \I__13181\ : InMux
    port map (
            O => \N__53947\,
            I => \N__53806\
        );

    \I__13180\ : InMux
    port map (
            O => \N__53946\,
            I => \N__53806\
        );

    \I__13179\ : InMux
    port map (
            O => \N__53945\,
            I => \N__53806\
        );

    \I__13178\ : InMux
    port map (
            O => \N__53944\,
            I => \N__53806\
        );

    \I__13177\ : InMux
    port map (
            O => \N__53943\,
            I => \N__53806\
        );

    \I__13176\ : InMux
    port map (
            O => \N__53942\,
            I => \N__53806\
        );

    \I__13175\ : InMux
    port map (
            O => \N__53941\,
            I => \N__53791\
        );

    \I__13174\ : InMux
    port map (
            O => \N__53940\,
            I => \N__53791\
        );

    \I__13173\ : InMux
    port map (
            O => \N__53939\,
            I => \N__53791\
        );

    \I__13172\ : InMux
    port map (
            O => \N__53938\,
            I => \N__53791\
        );

    \I__13171\ : InMux
    port map (
            O => \N__53937\,
            I => \N__53791\
        );

    \I__13170\ : InMux
    port map (
            O => \N__53936\,
            I => \N__53791\
        );

    \I__13169\ : InMux
    port map (
            O => \N__53935\,
            I => \N__53791\
        );

    \I__13168\ : LocalMux
    port map (
            O => \N__53932\,
            I => \N__53780\
        );

    \I__13167\ : LocalMux
    port map (
            O => \N__53929\,
            I => \N__53780\
        );

    \I__13166\ : LocalMux
    port map (
            O => \N__53926\,
            I => \N__53780\
        );

    \I__13165\ : Span4Mux_v
    port map (
            O => \N__53923\,
            I => \N__53780\
        );

    \I__13164\ : LocalMux
    port map (
            O => \N__53920\,
            I => \N__53780\
        );

    \I__13163\ : Span4Mux_v
    port map (
            O => \N__53913\,
            I => \N__53777\
        );

    \I__13162\ : InMux
    port map (
            O => \N__53910\,
            I => \N__53774\
        );

    \I__13161\ : InMux
    port map (
            O => \N__53909\,
            I => \N__53771\
        );

    \I__13160\ : InMux
    port map (
            O => \N__53908\,
            I => \N__53768\
        );

    \I__13159\ : LocalMux
    port map (
            O => \N__53905\,
            I => \N__53765\
        );

    \I__13158\ : InMux
    port map (
            O => \N__53904\,
            I => \N__53756\
        );

    \I__13157\ : InMux
    port map (
            O => \N__53903\,
            I => \N__53756\
        );

    \I__13156\ : InMux
    port map (
            O => \N__53902\,
            I => \N__53756\
        );

    \I__13155\ : InMux
    port map (
            O => \N__53901\,
            I => \N__53756\
        );

    \I__13154\ : InMux
    port map (
            O => \N__53900\,
            I => \N__53753\
        );

    \I__13153\ : Span4Mux_h
    port map (
            O => \N__53895\,
            I => \N__53750\
        );

    \I__13152\ : LocalMux
    port map (
            O => \N__53892\,
            I => \N__53743\
        );

    \I__13151\ : LocalMux
    port map (
            O => \N__53889\,
            I => \N__53743\
        );

    \I__13150\ : LocalMux
    port map (
            O => \N__53886\,
            I => \N__53743\
        );

    \I__13149\ : InMux
    port map (
            O => \N__53885\,
            I => \N__53733\
        );

    \I__13148\ : InMux
    port map (
            O => \N__53884\,
            I => \N__53733\
        );

    \I__13147\ : InMux
    port map (
            O => \N__53883\,
            I => \N__53733\
        );

    \I__13146\ : InMux
    port map (
            O => \N__53882\,
            I => \N__53728\
        );

    \I__13145\ : InMux
    port map (
            O => \N__53881\,
            I => \N__53728\
        );

    \I__13144\ : LocalMux
    port map (
            O => \N__53878\,
            I => \N__53723\
        );

    \I__13143\ : LocalMux
    port map (
            O => \N__53875\,
            I => \N__53723\
        );

    \I__13142\ : InMux
    port map (
            O => \N__53874\,
            I => \N__53720\
        );

    \I__13141\ : InMux
    port map (
            O => \N__53873\,
            I => \N__53713\
        );

    \I__13140\ : InMux
    port map (
            O => \N__53872\,
            I => \N__53713\
        );

    \I__13139\ : InMux
    port map (
            O => \N__53871\,
            I => \N__53713\
        );

    \I__13138\ : LocalMux
    port map (
            O => \N__53854\,
            I => \N__53704\
        );

    \I__13137\ : Span4Mux_v
    port map (
            O => \N__53851\,
            I => \N__53704\
        );

    \I__13136\ : Span4Mux_h
    port map (
            O => \N__53848\,
            I => \N__53704\
        );

    \I__13135\ : Span4Mux_h
    port map (
            O => \N__53843\,
            I => \N__53704\
        );

    \I__13134\ : Span4Mux_h
    port map (
            O => \N__53840\,
            I => \N__53701\
        );

    \I__13133\ : InMux
    port map (
            O => \N__53839\,
            I => \N__53696\
        );

    \I__13132\ : InMux
    port map (
            O => \N__53838\,
            I => \N__53696\
        );

    \I__13131\ : InMux
    port map (
            O => \N__53837\,
            I => \N__53693\
        );

    \I__13130\ : LocalMux
    port map (
            O => \N__53834\,
            I => \N__53688\
        );

    \I__13129\ : LocalMux
    port map (
            O => \N__53831\,
            I => \N__53688\
        );

    \I__13128\ : CascadeMux
    port map (
            O => \N__53830\,
            I => \N__53682\
        );

    \I__13127\ : InMux
    port map (
            O => \N__53829\,
            I => \N__53676\
        );

    \I__13126\ : InMux
    port map (
            O => \N__53828\,
            I => \N__53673\
        );

    \I__13125\ : Span4Mux_v
    port map (
            O => \N__53823\,
            I => \N__53670\
        );

    \I__13124\ : LocalMux
    port map (
            O => \N__53806\,
            I => \N__53659\
        );

    \I__13123\ : LocalMux
    port map (
            O => \N__53791\,
            I => \N__53659\
        );

    \I__13122\ : Span4Mux_v
    port map (
            O => \N__53780\,
            I => \N__53659\
        );

    \I__13121\ : Span4Mux_h
    port map (
            O => \N__53777\,
            I => \N__53659\
        );

    \I__13120\ : LocalMux
    port map (
            O => \N__53774\,
            I => \N__53659\
        );

    \I__13119\ : LocalMux
    port map (
            O => \N__53771\,
            I => \N__53645\
        );

    \I__13118\ : LocalMux
    port map (
            O => \N__53768\,
            I => \N__53645\
        );

    \I__13117\ : Sp12to4
    port map (
            O => \N__53765\,
            I => \N__53645\
        );

    \I__13116\ : LocalMux
    port map (
            O => \N__53756\,
            I => \N__53645\
        );

    \I__13115\ : LocalMux
    port map (
            O => \N__53753\,
            I => \N__53638\
        );

    \I__13114\ : Span4Mux_h
    port map (
            O => \N__53750\,
            I => \N__53638\
        );

    \I__13113\ : Span4Mux_v
    port map (
            O => \N__53743\,
            I => \N__53638\
        );

    \I__13112\ : InMux
    port map (
            O => \N__53742\,
            I => \N__53630\
        );

    \I__13111\ : InMux
    port map (
            O => \N__53741\,
            I => \N__53630\
        );

    \I__13110\ : InMux
    port map (
            O => \N__53740\,
            I => \N__53630\
        );

    \I__13109\ : LocalMux
    port map (
            O => \N__53733\,
            I => \N__53623\
        );

    \I__13108\ : LocalMux
    port map (
            O => \N__53728\,
            I => \N__53623\
        );

    \I__13107\ : Span4Mux_v
    port map (
            O => \N__53723\,
            I => \N__53623\
        );

    \I__13106\ : LocalMux
    port map (
            O => \N__53720\,
            I => \N__53608\
        );

    \I__13105\ : LocalMux
    port map (
            O => \N__53713\,
            I => \N__53608\
        );

    \I__13104\ : Span4Mux_h
    port map (
            O => \N__53704\,
            I => \N__53608\
        );

    \I__13103\ : Span4Mux_h
    port map (
            O => \N__53701\,
            I => \N__53608\
        );

    \I__13102\ : LocalMux
    port map (
            O => \N__53696\,
            I => \N__53608\
        );

    \I__13101\ : LocalMux
    port map (
            O => \N__53693\,
            I => \N__53608\
        );

    \I__13100\ : Span4Mux_v
    port map (
            O => \N__53688\,
            I => \N__53608\
        );

    \I__13099\ : InMux
    port map (
            O => \N__53687\,
            I => \N__53601\
        );

    \I__13098\ : InMux
    port map (
            O => \N__53686\,
            I => \N__53601\
        );

    \I__13097\ : InMux
    port map (
            O => \N__53685\,
            I => \N__53601\
        );

    \I__13096\ : InMux
    port map (
            O => \N__53682\,
            I => \N__53592\
        );

    \I__13095\ : InMux
    port map (
            O => \N__53681\,
            I => \N__53592\
        );

    \I__13094\ : InMux
    port map (
            O => \N__53680\,
            I => \N__53592\
        );

    \I__13093\ : InMux
    port map (
            O => \N__53679\,
            I => \N__53592\
        );

    \I__13092\ : LocalMux
    port map (
            O => \N__53676\,
            I => \N__53587\
        );

    \I__13091\ : LocalMux
    port map (
            O => \N__53673\,
            I => \N__53587\
        );

    \I__13090\ : Span4Mux_h
    port map (
            O => \N__53670\,
            I => \N__53582\
        );

    \I__13089\ : Span4Mux_v
    port map (
            O => \N__53659\,
            I => \N__53582\
        );

    \I__13088\ : InMux
    port map (
            O => \N__53658\,
            I => \N__53571\
        );

    \I__13087\ : InMux
    port map (
            O => \N__53657\,
            I => \N__53571\
        );

    \I__13086\ : InMux
    port map (
            O => \N__53656\,
            I => \N__53571\
        );

    \I__13085\ : InMux
    port map (
            O => \N__53655\,
            I => \N__53571\
        );

    \I__13084\ : InMux
    port map (
            O => \N__53654\,
            I => \N__53571\
        );

    \I__13083\ : Span12Mux_v
    port map (
            O => \N__53645\,
            I => \N__53568\
        );

    \I__13082\ : Span4Mux_v
    port map (
            O => \N__53638\,
            I => \N__53565\
        );

    \I__13081\ : InMux
    port map (
            O => \N__53637\,
            I => \N__53562\
        );

    \I__13080\ : LocalMux
    port map (
            O => \N__53630\,
            I => \N__53555\
        );

    \I__13079\ : Span4Mux_v
    port map (
            O => \N__53623\,
            I => \N__53555\
        );

    \I__13078\ : Span4Mux_v
    port map (
            O => \N__53608\,
            I => \N__53555\
        );

    \I__13077\ : LocalMux
    port map (
            O => \N__53601\,
            I => comm_state_1
        );

    \I__13076\ : LocalMux
    port map (
            O => \N__53592\,
            I => comm_state_1
        );

    \I__13075\ : Odrv12
    port map (
            O => \N__53587\,
            I => comm_state_1
        );

    \I__13074\ : Odrv4
    port map (
            O => \N__53582\,
            I => comm_state_1
        );

    \I__13073\ : LocalMux
    port map (
            O => \N__53571\,
            I => comm_state_1
        );

    \I__13072\ : Odrv12
    port map (
            O => \N__53568\,
            I => comm_state_1
        );

    \I__13071\ : Odrv4
    port map (
            O => \N__53565\,
            I => comm_state_1
        );

    \I__13070\ : LocalMux
    port map (
            O => \N__53562\,
            I => comm_state_1
        );

    \I__13069\ : Odrv4
    port map (
            O => \N__53555\,
            I => comm_state_1
        );

    \I__13068\ : InMux
    port map (
            O => \N__53536\,
            I => \N__53533\
        );

    \I__13067\ : LocalMux
    port map (
            O => \N__53533\,
            I => \N__53526\
        );

    \I__13066\ : CascadeMux
    port map (
            O => \N__53532\,
            I => \N__53523\
        );

    \I__13065\ : CascadeMux
    port map (
            O => \N__53531\,
            I => \N__53518\
        );

    \I__13064\ : InMux
    port map (
            O => \N__53530\,
            I => \N__53513\
        );

    \I__13063\ : InMux
    port map (
            O => \N__53529\,
            I => \N__53513\
        );

    \I__13062\ : Span4Mux_h
    port map (
            O => \N__53526\,
            I => \N__53506\
        );

    \I__13061\ : InMux
    port map (
            O => \N__53523\,
            I => \N__53503\
        );

    \I__13060\ : InMux
    port map (
            O => \N__53522\,
            I => \N__53500\
        );

    \I__13059\ : CascadeMux
    port map (
            O => \N__53521\,
            I => \N__53482\
        );

    \I__13058\ : InMux
    port map (
            O => \N__53518\,
            I => \N__53479\
        );

    \I__13057\ : LocalMux
    port map (
            O => \N__53513\,
            I => \N__53476\
        );

    \I__13056\ : InMux
    port map (
            O => \N__53512\,
            I => \N__53467\
        );

    \I__13055\ : InMux
    port map (
            O => \N__53511\,
            I => \N__53467\
        );

    \I__13054\ : InMux
    port map (
            O => \N__53510\,
            I => \N__53467\
        );

    \I__13053\ : InMux
    port map (
            O => \N__53509\,
            I => \N__53463\
        );

    \I__13052\ : Span4Mux_h
    port map (
            O => \N__53506\,
            I => \N__53454\
        );

    \I__13051\ : LocalMux
    port map (
            O => \N__53503\,
            I => \N__53454\
        );

    \I__13050\ : LocalMux
    port map (
            O => \N__53500\,
            I => \N__53454\
        );

    \I__13049\ : InMux
    port map (
            O => \N__53499\,
            I => \N__53451\
        );

    \I__13048\ : InMux
    port map (
            O => \N__53498\,
            I => \N__53439\
        );

    \I__13047\ : InMux
    port map (
            O => \N__53497\,
            I => \N__53439\
        );

    \I__13046\ : InMux
    port map (
            O => \N__53496\,
            I => \N__53439\
        );

    \I__13045\ : InMux
    port map (
            O => \N__53495\,
            I => \N__53439\
        );

    \I__13044\ : InMux
    port map (
            O => \N__53494\,
            I => \N__53432\
        );

    \I__13043\ : InMux
    port map (
            O => \N__53493\,
            I => \N__53432\
        );

    \I__13042\ : InMux
    port map (
            O => \N__53492\,
            I => \N__53421\
        );

    \I__13041\ : InMux
    port map (
            O => \N__53491\,
            I => \N__53421\
        );

    \I__13040\ : InMux
    port map (
            O => \N__53490\,
            I => \N__53421\
        );

    \I__13039\ : InMux
    port map (
            O => \N__53489\,
            I => \N__53421\
        );

    \I__13038\ : InMux
    port map (
            O => \N__53488\,
            I => \N__53421\
        );

    \I__13037\ : InMux
    port map (
            O => \N__53487\,
            I => \N__53418\
        );

    \I__13036\ : InMux
    port map (
            O => \N__53486\,
            I => \N__53414\
        );

    \I__13035\ : InMux
    port map (
            O => \N__53485\,
            I => \N__53411\
        );

    \I__13034\ : InMux
    port map (
            O => \N__53482\,
            I => \N__53408\
        );

    \I__13033\ : LocalMux
    port map (
            O => \N__53479\,
            I => \N__53403\
        );

    \I__13032\ : Span4Mux_v
    port map (
            O => \N__53476\,
            I => \N__53403\
        );

    \I__13031\ : InMux
    port map (
            O => \N__53475\,
            I => \N__53398\
        );

    \I__13030\ : InMux
    port map (
            O => \N__53474\,
            I => \N__53398\
        );

    \I__13029\ : LocalMux
    port map (
            O => \N__53467\,
            I => \N__53395\
        );

    \I__13028\ : InMux
    port map (
            O => \N__53466\,
            I => \N__53392\
        );

    \I__13027\ : LocalMux
    port map (
            O => \N__53463\,
            I => \N__53389\
        );

    \I__13026\ : InMux
    port map (
            O => \N__53462\,
            I => \N__53384\
        );

    \I__13025\ : InMux
    port map (
            O => \N__53461\,
            I => \N__53384\
        );

    \I__13024\ : Span4Mux_v
    port map (
            O => \N__53454\,
            I => \N__53379\
        );

    \I__13023\ : LocalMux
    port map (
            O => \N__53451\,
            I => \N__53379\
        );

    \I__13022\ : InMux
    port map (
            O => \N__53450\,
            I => \N__53372\
        );

    \I__13021\ : InMux
    port map (
            O => \N__53449\,
            I => \N__53372\
        );

    \I__13020\ : InMux
    port map (
            O => \N__53448\,
            I => \N__53372\
        );

    \I__13019\ : LocalMux
    port map (
            O => \N__53439\,
            I => \N__53368\
        );

    \I__13018\ : InMux
    port map (
            O => \N__53438\,
            I => \N__53365\
        );

    \I__13017\ : InMux
    port map (
            O => \N__53437\,
            I => \N__53362\
        );

    \I__13016\ : LocalMux
    port map (
            O => \N__53432\,
            I => \N__53358\
        );

    \I__13015\ : LocalMux
    port map (
            O => \N__53421\,
            I => \N__53353\
        );

    \I__13014\ : LocalMux
    port map (
            O => \N__53418\,
            I => \N__53353\
        );

    \I__13013\ : InMux
    port map (
            O => \N__53417\,
            I => \N__53350\
        );

    \I__13012\ : LocalMux
    port map (
            O => \N__53414\,
            I => \N__53345\
        );

    \I__13011\ : LocalMux
    port map (
            O => \N__53411\,
            I => \N__53345\
        );

    \I__13010\ : LocalMux
    port map (
            O => \N__53408\,
            I => \N__53340\
        );

    \I__13009\ : Span4Mux_h
    port map (
            O => \N__53403\,
            I => \N__53340\
        );

    \I__13008\ : LocalMux
    port map (
            O => \N__53398\,
            I => \N__53337\
        );

    \I__13007\ : Span4Mux_v
    port map (
            O => \N__53395\,
            I => \N__53332\
        );

    \I__13006\ : LocalMux
    port map (
            O => \N__53392\,
            I => \N__53332\
        );

    \I__13005\ : Sp12to4
    port map (
            O => \N__53389\,
            I => \N__53327\
        );

    \I__13004\ : LocalMux
    port map (
            O => \N__53384\,
            I => \N__53327\
        );

    \I__13003\ : Span4Mux_h
    port map (
            O => \N__53379\,
            I => \N__53324\
        );

    \I__13002\ : LocalMux
    port map (
            O => \N__53372\,
            I => \N__53321\
        );

    \I__13001\ : InMux
    port map (
            O => \N__53371\,
            I => \N__53318\
        );

    \I__13000\ : Span4Mux_h
    port map (
            O => \N__53368\,
            I => \N__53311\
        );

    \I__12999\ : LocalMux
    port map (
            O => \N__53365\,
            I => \N__53311\
        );

    \I__12998\ : LocalMux
    port map (
            O => \N__53362\,
            I => \N__53311\
        );

    \I__12997\ : InMux
    port map (
            O => \N__53361\,
            I => \N__53308\
        );

    \I__12996\ : Span4Mux_v
    port map (
            O => \N__53358\,
            I => \N__53303\
        );

    \I__12995\ : Span4Mux_v
    port map (
            O => \N__53353\,
            I => \N__53303\
        );

    \I__12994\ : LocalMux
    port map (
            O => \N__53350\,
            I => \N__53300\
        );

    \I__12993\ : Span4Mux_v
    port map (
            O => \N__53345\,
            I => \N__53291\
        );

    \I__12992\ : Span4Mux_h
    port map (
            O => \N__53340\,
            I => \N__53291\
        );

    \I__12991\ : Span4Mux_v
    port map (
            O => \N__53337\,
            I => \N__53291\
        );

    \I__12990\ : Span4Mux_v
    port map (
            O => \N__53332\,
            I => \N__53291\
        );

    \I__12989\ : Span12Mux_v
    port map (
            O => \N__53327\,
            I => \N__53288\
        );

    \I__12988\ : Span4Mux_h
    port map (
            O => \N__53324\,
            I => \N__53285\
        );

    \I__12987\ : Odrv12
    port map (
            O => \N__53321\,
            I => comm_state_0
        );

    \I__12986\ : LocalMux
    port map (
            O => \N__53318\,
            I => comm_state_0
        );

    \I__12985\ : Odrv4
    port map (
            O => \N__53311\,
            I => comm_state_0
        );

    \I__12984\ : LocalMux
    port map (
            O => \N__53308\,
            I => comm_state_0
        );

    \I__12983\ : Odrv4
    port map (
            O => \N__53303\,
            I => comm_state_0
        );

    \I__12982\ : Odrv4
    port map (
            O => \N__53300\,
            I => comm_state_0
        );

    \I__12981\ : Odrv4
    port map (
            O => \N__53291\,
            I => comm_state_0
        );

    \I__12980\ : Odrv12
    port map (
            O => \N__53288\,
            I => comm_state_0
        );

    \I__12979\ : Odrv4
    port map (
            O => \N__53285\,
            I => comm_state_0
        );

    \I__12978\ : CEMux
    port map (
            O => \N__53266\,
            I => \N__53263\
        );

    \I__12977\ : LocalMux
    port map (
            O => \N__53263\,
            I => n11347
        );

    \I__12976\ : InMux
    port map (
            O => \N__53260\,
            I => \N__53255\
        );

    \I__12975\ : InMux
    port map (
            O => \N__53259\,
            I => \N__53250\
        );

    \I__12974\ : InMux
    port map (
            O => \N__53258\,
            I => \N__53250\
        );

    \I__12973\ : LocalMux
    port map (
            O => \N__53255\,
            I => \N__53247\
        );

    \I__12972\ : LocalMux
    port map (
            O => \N__53250\,
            I => \N__53244\
        );

    \I__12971\ : Span4Mux_v
    port map (
            O => \N__53247\,
            I => \N__53239\
        );

    \I__12970\ : Span4Mux_v
    port map (
            O => \N__53244\,
            I => \N__53239\
        );

    \I__12969\ : Span4Mux_h
    port map (
            O => \N__53239\,
            I => \N__53236\
        );

    \I__12968\ : Odrv4
    port map (
            O => \N__53236\,
            I => comm_tx_buf_0
        );

    \I__12967\ : InMux
    port map (
            O => \N__53233\,
            I => \N__53230\
        );

    \I__12966\ : LocalMux
    port map (
            O => \N__53230\,
            I => \N__53225\
        );

    \I__12965\ : InMux
    port map (
            O => \N__53229\,
            I => \N__53222\
        );

    \I__12964\ : InMux
    port map (
            O => \N__53228\,
            I => \N__53219\
        );

    \I__12963\ : Odrv4
    port map (
            O => \N__53225\,
            I => \comm_spi.n22650\
        );

    \I__12962\ : LocalMux
    port map (
            O => \N__53222\,
            I => \comm_spi.n22650\
        );

    \I__12961\ : LocalMux
    port map (
            O => \N__53219\,
            I => \comm_spi.n22650\
        );

    \I__12960\ : SRMux
    port map (
            O => \N__53212\,
            I => \N__53209\
        );

    \I__12959\ : LocalMux
    port map (
            O => \N__53209\,
            I => \N__53206\
        );

    \I__12958\ : Span4Mux_v
    port map (
            O => \N__53206\,
            I => \N__53203\
        );

    \I__12957\ : Odrv4
    port map (
            O => \N__53203\,
            I => \comm_spi.data_tx_7__N_764\
        );

    \I__12956\ : InMux
    port map (
            O => \N__53200\,
            I => \N__53194\
        );

    \I__12955\ : InMux
    port map (
            O => \N__53199\,
            I => \N__53194\
        );

    \I__12954\ : LocalMux
    port map (
            O => \N__53194\,
            I => \N__53190\
        );

    \I__12953\ : InMux
    port map (
            O => \N__53193\,
            I => \N__53187\
        );

    \I__12952\ : Span4Mux_v
    port map (
            O => \N__53190\,
            I => \N__53184\
        );

    \I__12951\ : LocalMux
    port map (
            O => \N__53187\,
            I => \N__53181\
        );

    \I__12950\ : Odrv4
    port map (
            O => \N__53184\,
            I => comm_tx_buf_1
        );

    \I__12949\ : Odrv4
    port map (
            O => \N__53181\,
            I => comm_tx_buf_1
        );

    \I__12948\ : SRMux
    port map (
            O => \N__53176\,
            I => \N__53173\
        );

    \I__12947\ : LocalMux
    port map (
            O => \N__53173\,
            I => \N__53170\
        );

    \I__12946\ : Sp12to4
    port map (
            O => \N__53170\,
            I => \N__53167\
        );

    \I__12945\ : Odrv12
    port map (
            O => \N__53167\,
            I => \comm_spi.data_tx_7__N_784\
        );

    \I__12944\ : InMux
    port map (
            O => \N__53164\,
            I => \N__53161\
        );

    \I__12943\ : LocalMux
    port map (
            O => \N__53161\,
            I => \N__53157\
        );

    \I__12942\ : InMux
    port map (
            O => \N__53160\,
            I => \N__53154\
        );

    \I__12941\ : Span4Mux_h
    port map (
            O => \N__53157\,
            I => \N__53149\
        );

    \I__12940\ : LocalMux
    port map (
            O => \N__53154\,
            I => \N__53149\
        );

    \I__12939\ : Span4Mux_v
    port map (
            O => \N__53149\,
            I => \N__53145\
        );

    \I__12938\ : InMux
    port map (
            O => \N__53148\,
            I => \N__53142\
        );

    \I__12937\ : Span4Mux_h
    port map (
            O => \N__53145\,
            I => \N__53139\
        );

    \I__12936\ : LocalMux
    port map (
            O => \N__53142\,
            I => \N__53136\
        );

    \I__12935\ : Odrv4
    port map (
            O => \N__53139\,
            I => comm_tx_buf_4
        );

    \I__12934\ : Odrv4
    port map (
            O => \N__53136\,
            I => comm_tx_buf_4
        );

    \I__12933\ : SRMux
    port map (
            O => \N__53131\,
            I => \N__53128\
        );

    \I__12932\ : LocalMux
    port map (
            O => \N__53128\,
            I => \N__53125\
        );

    \I__12931\ : Span4Mux_v
    port map (
            O => \N__53125\,
            I => \N__53122\
        );

    \I__12930\ : Odrv4
    port map (
            O => \N__53122\,
            I => \comm_spi.data_tx_7__N_775\
        );

    \I__12929\ : CascadeMux
    port map (
            O => \N__53119\,
            I => \n20502_cascade_\
        );

    \I__12928\ : InMux
    port map (
            O => \N__53116\,
            I => \N__53113\
        );

    \I__12927\ : LocalMux
    port map (
            O => \N__53113\,
            I => n12_adj_1583
        );

    \I__12926\ : InMux
    port map (
            O => \N__53110\,
            I => \N__53107\
        );

    \I__12925\ : LocalMux
    port map (
            O => \N__53107\,
            I => n20502
        );

    \I__12924\ : InMux
    port map (
            O => \N__53104\,
            I => \N__53100\
        );

    \I__12923\ : InMux
    port map (
            O => \N__53103\,
            I => \N__53097\
        );

    \I__12922\ : LocalMux
    port map (
            O => \N__53100\,
            I => \N__53094\
        );

    \I__12921\ : LocalMux
    port map (
            O => \N__53097\,
            I => secclk_cnt_19
        );

    \I__12920\ : Odrv12
    port map (
            O => \N__53094\,
            I => secclk_cnt_19
        );

    \I__12919\ : InMux
    port map (
            O => \N__53089\,
            I => \N__53085\
        );

    \I__12918\ : InMux
    port map (
            O => \N__53088\,
            I => \N__53082\
        );

    \I__12917\ : LocalMux
    port map (
            O => \N__53085\,
            I => \N__53079\
        );

    \I__12916\ : LocalMux
    port map (
            O => \N__53082\,
            I => secclk_cnt_21
        );

    \I__12915\ : Odrv12
    port map (
            O => \N__53079\,
            I => secclk_cnt_21
        );

    \I__12914\ : CascadeMux
    port map (
            O => \N__53074\,
            I => \N__53071\
        );

    \I__12913\ : InMux
    port map (
            O => \N__53071\,
            I => \N__53068\
        );

    \I__12912\ : LocalMux
    port map (
            O => \N__53068\,
            I => \N__53064\
        );

    \I__12911\ : InMux
    port map (
            O => \N__53067\,
            I => \N__53061\
        );

    \I__12910\ : Span4Mux_v
    port map (
            O => \N__53064\,
            I => \N__53058\
        );

    \I__12909\ : LocalMux
    port map (
            O => \N__53061\,
            I => secclk_cnt_12
        );

    \I__12908\ : Odrv4
    port map (
            O => \N__53058\,
            I => secclk_cnt_12
        );

    \I__12907\ : InMux
    port map (
            O => \N__53053\,
            I => \N__53049\
        );

    \I__12906\ : InMux
    port map (
            O => \N__53052\,
            I => \N__53046\
        );

    \I__12905\ : LocalMux
    port map (
            O => \N__53049\,
            I => \N__53043\
        );

    \I__12904\ : LocalMux
    port map (
            O => \N__53046\,
            I => secclk_cnt_22
        );

    \I__12903\ : Odrv12
    port map (
            O => \N__53043\,
            I => secclk_cnt_22
        );

    \I__12902\ : InMux
    port map (
            O => \N__53038\,
            I => \N__53035\
        );

    \I__12901\ : LocalMux
    port map (
            O => \N__53035\,
            I => \N__53032\
        );

    \I__12900\ : Span4Mux_h
    port map (
            O => \N__53032\,
            I => \N__53029\
        );

    \I__12899\ : Odrv4
    port map (
            O => \N__53029\,
            I => n14_adj_1578
        );

    \I__12898\ : CascadeMux
    port map (
            O => \N__53026\,
            I => \N__53022\
        );

    \I__12897\ : CascadeMux
    port map (
            O => \N__53025\,
            I => \N__53019\
        );

    \I__12896\ : InMux
    port map (
            O => \N__53022\,
            I => \N__53015\
        );

    \I__12895\ : InMux
    port map (
            O => \N__53019\,
            I => \N__53012\
        );

    \I__12894\ : CascadeMux
    port map (
            O => \N__53018\,
            I => \N__53009\
        );

    \I__12893\ : LocalMux
    port map (
            O => \N__53015\,
            I => \N__53006\
        );

    \I__12892\ : LocalMux
    port map (
            O => \N__53012\,
            I => \N__53002\
        );

    \I__12891\ : InMux
    port map (
            O => \N__53009\,
            I => \N__52999\
        );

    \I__12890\ : Span4Mux_h
    port map (
            O => \N__53006\,
            I => \N__52996\
        );

    \I__12889\ : CascadeMux
    port map (
            O => \N__53005\,
            I => \N__52993\
        );

    \I__12888\ : Span4Mux_h
    port map (
            O => \N__53002\,
            I => \N__52990\
        );

    \I__12887\ : LocalMux
    port map (
            O => \N__52999\,
            I => \N__52985\
        );

    \I__12886\ : Span4Mux_h
    port map (
            O => \N__52996\,
            I => \N__52985\
        );

    \I__12885\ : InMux
    port map (
            O => \N__52993\,
            I => \N__52982\
        );

    \I__12884\ : Span4Mux_h
    port map (
            O => \N__52990\,
            I => \N__52979\
        );

    \I__12883\ : Span4Mux_h
    port map (
            O => \N__52985\,
            I => \N__52976\
        );

    \I__12882\ : LocalMux
    port map (
            O => \N__52982\,
            I => trig_dds0
        );

    \I__12881\ : Odrv4
    port map (
            O => \N__52979\,
            I => trig_dds0
        );

    \I__12880\ : Odrv4
    port map (
            O => \N__52976\,
            I => trig_dds0
        );

    \I__12879\ : InMux
    port map (
            O => \N__52969\,
            I => \N__52966\
        );

    \I__12878\ : LocalMux
    port map (
            O => \N__52966\,
            I => \N__52963\
        );

    \I__12877\ : Odrv12
    port map (
            O => \N__52963\,
            I => \comm_spi.n14582\
        );

    \I__12876\ : InMux
    port map (
            O => \N__52960\,
            I => \N__52957\
        );

    \I__12875\ : LocalMux
    port map (
            O => \N__52957\,
            I => \N__52954\
        );

    \I__12874\ : Span4Mux_v
    port map (
            O => \N__52954\,
            I => \N__52949\
        );

    \I__12873\ : InMux
    port map (
            O => \N__52953\,
            I => \N__52946\
        );

    \I__12872\ : InMux
    port map (
            O => \N__52952\,
            I => \N__52943\
        );

    \I__12871\ : Sp12to4
    port map (
            O => \N__52949\,
            I => \N__52938\
        );

    \I__12870\ : LocalMux
    port map (
            O => \N__52946\,
            I => \N__52933\
        );

    \I__12869\ : LocalMux
    port map (
            O => \N__52943\,
            I => \N__52933\
        );

    \I__12868\ : InMux
    port map (
            O => \N__52942\,
            I => \N__52930\
        );

    \I__12867\ : InMux
    port map (
            O => \N__52941\,
            I => \N__52927\
        );

    \I__12866\ : Span12Mux_h
    port map (
            O => \N__52938\,
            I => \N__52924\
        );

    \I__12865\ : Sp12to4
    port map (
            O => \N__52933\,
            I => \N__52917\
        );

    \I__12864\ : LocalMux
    port map (
            O => \N__52930\,
            I => \N__52917\
        );

    \I__12863\ : LocalMux
    port map (
            O => \N__52927\,
            I => \N__52917\
        );

    \I__12862\ : Span12Mux_v
    port map (
            O => \N__52924\,
            I => \N__52914\
        );

    \I__12861\ : Span12Mux_v
    port map (
            O => \N__52917\,
            I => \N__52911\
        );

    \I__12860\ : Odrv12
    port map (
            O => \N__52914\,
            I => \ICE_SPI_SCLK\
        );

    \I__12859\ : Odrv12
    port map (
            O => \N__52911\,
            I => \ICE_SPI_SCLK\
        );

    \I__12858\ : SRMux
    port map (
            O => \N__52906\,
            I => \N__52903\
        );

    \I__12857\ : LocalMux
    port map (
            O => \N__52903\,
            I => \N__52900\
        );

    \I__12856\ : Odrv4
    port map (
            O => \N__52900\,
            I => \comm_spi.iclk_N_755\
        );

    \I__12855\ : SRMux
    port map (
            O => \N__52897\,
            I => \N__52894\
        );

    \I__12854\ : LocalMux
    port map (
            O => \N__52894\,
            I => \N__52891\
        );

    \I__12853\ : Odrv4
    port map (
            O => \N__52891\,
            I => \comm_spi.data_tx_7__N_765\
        );

    \I__12852\ : SRMux
    port map (
            O => \N__52888\,
            I => \N__52883\
        );

    \I__12851\ : SRMux
    port map (
            O => \N__52887\,
            I => \N__52880\
        );

    \I__12850\ : SRMux
    port map (
            O => \N__52886\,
            I => \N__52874\
        );

    \I__12849\ : LocalMux
    port map (
            O => \N__52883\,
            I => \N__52868\
        );

    \I__12848\ : LocalMux
    port map (
            O => \N__52880\,
            I => \N__52868\
        );

    \I__12847\ : SRMux
    port map (
            O => \N__52879\,
            I => \N__52865\
        );

    \I__12846\ : SRMux
    port map (
            O => \N__52878\,
            I => \N__52862\
        );

    \I__12845\ : IoInMux
    port map (
            O => \N__52877\,
            I => \N__52857\
        );

    \I__12844\ : LocalMux
    port map (
            O => \N__52874\,
            I => \N__52854\
        );

    \I__12843\ : SRMux
    port map (
            O => \N__52873\,
            I => \N__52851\
        );

    \I__12842\ : Span4Mux_v
    port map (
            O => \N__52868\,
            I => \N__52844\
        );

    \I__12841\ : LocalMux
    port map (
            O => \N__52865\,
            I => \N__52844\
        );

    \I__12840\ : LocalMux
    port map (
            O => \N__52862\,
            I => \N__52844\
        );

    \I__12839\ : SRMux
    port map (
            O => \N__52861\,
            I => \N__52841\
        );

    \I__12838\ : SRMux
    port map (
            O => \N__52860\,
            I => \N__52838\
        );

    \I__12837\ : LocalMux
    port map (
            O => \N__52857\,
            I => \N__52832\
        );

    \I__12836\ : Span4Mux_v
    port map (
            O => \N__52854\,
            I => \N__52823\
        );

    \I__12835\ : LocalMux
    port map (
            O => \N__52851\,
            I => \N__52823\
        );

    \I__12834\ : Span4Mux_v
    port map (
            O => \N__52844\,
            I => \N__52816\
        );

    \I__12833\ : LocalMux
    port map (
            O => \N__52841\,
            I => \N__52816\
        );

    \I__12832\ : LocalMux
    port map (
            O => \N__52838\,
            I => \N__52816\
        );

    \I__12831\ : SRMux
    port map (
            O => \N__52837\,
            I => \N__52813\
        );

    \I__12830\ : SRMux
    port map (
            O => \N__52836\,
            I => \N__52806\
        );

    \I__12829\ : SRMux
    port map (
            O => \N__52835\,
            I => \N__52796\
        );

    \I__12828\ : Span4Mux_s0_v
    port map (
            O => \N__52832\,
            I => \N__52788\
        );

    \I__12827\ : CascadeMux
    port map (
            O => \N__52831\,
            I => \N__52785\
        );

    \I__12826\ : CascadeMux
    port map (
            O => \N__52830\,
            I => \N__52781\
        );

    \I__12825\ : CascadeMux
    port map (
            O => \N__52829\,
            I => \N__52777\
        );

    \I__12824\ : CascadeMux
    port map (
            O => \N__52828\,
            I => \N__52773\
        );

    \I__12823\ : Span4Mux_h
    port map (
            O => \N__52823\,
            I => \N__52766\
        );

    \I__12822\ : Span4Mux_v
    port map (
            O => \N__52816\,
            I => \N__52766\
        );

    \I__12821\ : LocalMux
    port map (
            O => \N__52813\,
            I => \N__52766\
        );

    \I__12820\ : CascadeMux
    port map (
            O => \N__52812\,
            I => \N__52763\
        );

    \I__12819\ : CascadeMux
    port map (
            O => \N__52811\,
            I => \N__52759\
        );

    \I__12818\ : CascadeMux
    port map (
            O => \N__52810\,
            I => \N__52755\
        );

    \I__12817\ : CascadeMux
    port map (
            O => \N__52809\,
            I => \N__52751\
        );

    \I__12816\ : LocalMux
    port map (
            O => \N__52806\,
            I => \N__52744\
        );

    \I__12815\ : InMux
    port map (
            O => \N__52805\,
            I => \N__52737\
        );

    \I__12814\ : InMux
    port map (
            O => \N__52804\,
            I => \N__52737\
        );

    \I__12813\ : InMux
    port map (
            O => \N__52803\,
            I => \N__52737\
        );

    \I__12812\ : InMux
    port map (
            O => \N__52802\,
            I => \N__52728\
        );

    \I__12811\ : InMux
    port map (
            O => \N__52801\,
            I => \N__52728\
        );

    \I__12810\ : InMux
    port map (
            O => \N__52800\,
            I => \N__52728\
        );

    \I__12809\ : InMux
    port map (
            O => \N__52799\,
            I => \N__52728\
        );

    \I__12808\ : LocalMux
    port map (
            O => \N__52796\,
            I => \N__52725\
        );

    \I__12807\ : InMux
    port map (
            O => \N__52795\,
            I => \N__52720\
        );

    \I__12806\ : CascadeMux
    port map (
            O => \N__52794\,
            I => \N__52716\
        );

    \I__12805\ : CascadeMux
    port map (
            O => \N__52793\,
            I => \N__52712\
        );

    \I__12804\ : CascadeMux
    port map (
            O => \N__52792\,
            I => \N__52708\
        );

    \I__12803\ : CascadeMux
    port map (
            O => \N__52791\,
            I => \N__52704\
        );

    \I__12802\ : Span4Mux_v
    port map (
            O => \N__52788\,
            I => \N__52701\
        );

    \I__12801\ : InMux
    port map (
            O => \N__52785\,
            I => \N__52686\
        );

    \I__12800\ : InMux
    port map (
            O => \N__52784\,
            I => \N__52686\
        );

    \I__12799\ : InMux
    port map (
            O => \N__52781\,
            I => \N__52686\
        );

    \I__12798\ : InMux
    port map (
            O => \N__52780\,
            I => \N__52686\
        );

    \I__12797\ : InMux
    port map (
            O => \N__52777\,
            I => \N__52686\
        );

    \I__12796\ : InMux
    port map (
            O => \N__52776\,
            I => \N__52686\
        );

    \I__12795\ : InMux
    port map (
            O => \N__52773\,
            I => \N__52686\
        );

    \I__12794\ : Span4Mux_v
    port map (
            O => \N__52766\,
            I => \N__52683\
        );

    \I__12793\ : InMux
    port map (
            O => \N__52763\,
            I => \N__52668\
        );

    \I__12792\ : InMux
    port map (
            O => \N__52762\,
            I => \N__52668\
        );

    \I__12791\ : InMux
    port map (
            O => \N__52759\,
            I => \N__52668\
        );

    \I__12790\ : InMux
    port map (
            O => \N__52758\,
            I => \N__52668\
        );

    \I__12789\ : InMux
    port map (
            O => \N__52755\,
            I => \N__52668\
        );

    \I__12788\ : InMux
    port map (
            O => \N__52754\,
            I => \N__52668\
        );

    \I__12787\ : InMux
    port map (
            O => \N__52751\,
            I => \N__52668\
        );

    \I__12786\ : CascadeMux
    port map (
            O => \N__52750\,
            I => \N__52664\
        );

    \I__12785\ : CascadeMux
    port map (
            O => \N__52749\,
            I => \N__52660\
        );

    \I__12784\ : CascadeMux
    port map (
            O => \N__52748\,
            I => \N__52656\
        );

    \I__12783\ : CascadeMux
    port map (
            O => \N__52747\,
            I => \N__52652\
        );

    \I__12782\ : Span4Mux_v
    port map (
            O => \N__52744\,
            I => \N__52649\
        );

    \I__12781\ : LocalMux
    port map (
            O => \N__52737\,
            I => \N__52644\
        );

    \I__12780\ : LocalMux
    port map (
            O => \N__52728\,
            I => \N__52644\
        );

    \I__12779\ : Span4Mux_v
    port map (
            O => \N__52725\,
            I => \N__52641\
        );

    \I__12778\ : InMux
    port map (
            O => \N__52724\,
            I => \N__52638\
        );

    \I__12777\ : SRMux
    port map (
            O => \N__52723\,
            I => \N__52635\
        );

    \I__12776\ : LocalMux
    port map (
            O => \N__52720\,
            I => \N__52632\
        );

    \I__12775\ : InMux
    port map (
            O => \N__52719\,
            I => \N__52615\
        );

    \I__12774\ : InMux
    port map (
            O => \N__52716\,
            I => \N__52615\
        );

    \I__12773\ : InMux
    port map (
            O => \N__52715\,
            I => \N__52615\
        );

    \I__12772\ : InMux
    port map (
            O => \N__52712\,
            I => \N__52615\
        );

    \I__12771\ : InMux
    port map (
            O => \N__52711\,
            I => \N__52615\
        );

    \I__12770\ : InMux
    port map (
            O => \N__52708\,
            I => \N__52615\
        );

    \I__12769\ : InMux
    port map (
            O => \N__52707\,
            I => \N__52615\
        );

    \I__12768\ : InMux
    port map (
            O => \N__52704\,
            I => \N__52615\
        );

    \I__12767\ : Span4Mux_v
    port map (
            O => \N__52701\,
            I => \N__52610\
        );

    \I__12766\ : LocalMux
    port map (
            O => \N__52686\,
            I => \N__52610\
        );

    \I__12765\ : Span4Mux_h
    port map (
            O => \N__52683\,
            I => \N__52605\
        );

    \I__12764\ : LocalMux
    port map (
            O => \N__52668\,
            I => \N__52605\
        );

    \I__12763\ : InMux
    port map (
            O => \N__52667\,
            I => \N__52588\
        );

    \I__12762\ : InMux
    port map (
            O => \N__52664\,
            I => \N__52588\
        );

    \I__12761\ : InMux
    port map (
            O => \N__52663\,
            I => \N__52588\
        );

    \I__12760\ : InMux
    port map (
            O => \N__52660\,
            I => \N__52588\
        );

    \I__12759\ : InMux
    port map (
            O => \N__52659\,
            I => \N__52588\
        );

    \I__12758\ : InMux
    port map (
            O => \N__52656\,
            I => \N__52588\
        );

    \I__12757\ : InMux
    port map (
            O => \N__52655\,
            I => \N__52588\
        );

    \I__12756\ : InMux
    port map (
            O => \N__52652\,
            I => \N__52588\
        );

    \I__12755\ : Span4Mux_h
    port map (
            O => \N__52649\,
            I => \N__52585\
        );

    \I__12754\ : Span4Mux_v
    port map (
            O => \N__52644\,
            I => \N__52582\
        );

    \I__12753\ : Sp12to4
    port map (
            O => \N__52641\,
            I => \N__52577\
        );

    \I__12752\ : LocalMux
    port map (
            O => \N__52638\,
            I => \N__52577\
        );

    \I__12751\ : LocalMux
    port map (
            O => \N__52635\,
            I => \N__52574\
        );

    \I__12750\ : Span4Mux_v
    port map (
            O => \N__52632\,
            I => \N__52571\
        );

    \I__12749\ : LocalMux
    port map (
            O => \N__52615\,
            I => \N__52568\
        );

    \I__12748\ : Span4Mux_h
    port map (
            O => \N__52610\,
            I => \N__52561\
        );

    \I__12747\ : Span4Mux_h
    port map (
            O => \N__52605\,
            I => \N__52561\
        );

    \I__12746\ : LocalMux
    port map (
            O => \N__52588\,
            I => \N__52561\
        );

    \I__12745\ : Span4Mux_h
    port map (
            O => \N__52585\,
            I => \N__52556\
        );

    \I__12744\ : Span4Mux_v
    port map (
            O => \N__52582\,
            I => \N__52556\
        );

    \I__12743\ : Span12Mux_s10_h
    port map (
            O => \N__52577\,
            I => \N__52551\
        );

    \I__12742\ : Span12Mux_s9_h
    port map (
            O => \N__52574\,
            I => \N__52551\
        );

    \I__12741\ : Span4Mux_h
    port map (
            O => \N__52571\,
            I => \N__52546\
        );

    \I__12740\ : Span4Mux_v
    port map (
            O => \N__52568\,
            I => \N__52546\
        );

    \I__12739\ : Sp12to4
    port map (
            O => \N__52561\,
            I => \N__52543\
        );

    \I__12738\ : Odrv4
    port map (
            O => \N__52556\,
            I => \CONSTANT_ONE_NET\
        );

    \I__12737\ : Odrv12
    port map (
            O => \N__52551\,
            I => \CONSTANT_ONE_NET\
        );

    \I__12736\ : Odrv4
    port map (
            O => \N__52546\,
            I => \CONSTANT_ONE_NET\
        );

    \I__12735\ : Odrv12
    port map (
            O => \N__52543\,
            I => \CONSTANT_ONE_NET\
        );

    \I__12734\ : SRMux
    port map (
            O => \N__52534\,
            I => \N__52531\
        );

    \I__12733\ : LocalMux
    port map (
            O => \N__52531\,
            I => \N__52528\
        );

    \I__12732\ : Sp12to4
    port map (
            O => \N__52528\,
            I => \N__52525\
        );

    \I__12731\ : Odrv12
    port map (
            O => \N__52525\,
            I => \comm_spi.data_tx_7__N_787\
        );

    \I__12730\ : InMux
    port map (
            O => \N__52522\,
            I => \N__52519\
        );

    \I__12729\ : LocalMux
    port map (
            O => \N__52519\,
            I => \N__52515\
        );

    \I__12728\ : InMux
    port map (
            O => \N__52518\,
            I => \N__52512\
        );

    \I__12727\ : Span4Mux_v
    port map (
            O => \N__52515\,
            I => \N__52507\
        );

    \I__12726\ : LocalMux
    port map (
            O => \N__52512\,
            I => \N__52507\
        );

    \I__12725\ : Span4Mux_h
    port map (
            O => \N__52507\,
            I => \N__52504\
        );

    \I__12724\ : Odrv4
    port map (
            O => \N__52504\,
            I => \comm_spi.n14604\
        );

    \I__12723\ : InMux
    port map (
            O => \N__52501\,
            I => \N__52498\
        );

    \I__12722\ : LocalMux
    port map (
            O => \N__52498\,
            I => \N__52494\
        );

    \I__12721\ : InMux
    port map (
            O => \N__52497\,
            I => \N__52491\
        );

    \I__12720\ : Odrv4
    port map (
            O => \N__52494\,
            I => \comm_spi.n14578\
        );

    \I__12719\ : LocalMux
    port map (
            O => \N__52491\,
            I => \comm_spi.n14578\
        );

    \I__12718\ : InMux
    port map (
            O => \N__52486\,
            I => \N__52483\
        );

    \I__12717\ : LocalMux
    port map (
            O => \N__52483\,
            I => \N__52479\
        );

    \I__12716\ : InMux
    port map (
            O => \N__52482\,
            I => \N__52476\
        );

    \I__12715\ : Span4Mux_v
    port map (
            O => \N__52479\,
            I => \N__52471\
        );

    \I__12714\ : LocalMux
    port map (
            O => \N__52476\,
            I => \N__52471\
        );

    \I__12713\ : Odrv4
    port map (
            O => \N__52471\,
            I => \comm_spi.n14577\
        );

    \I__12712\ : InMux
    port map (
            O => \N__52468\,
            I => \N__52465\
        );

    \I__12711\ : LocalMux
    port map (
            O => \N__52465\,
            I => \N__52462\
        );

    \I__12710\ : Span4Mux_h
    port map (
            O => \N__52462\,
            I => \N__52458\
        );

    \I__12709\ : InMux
    port map (
            O => \N__52461\,
            I => \N__52455\
        );

    \I__12708\ : Span4Mux_h
    port map (
            O => \N__52458\,
            I => \N__52452\
        );

    \I__12707\ : LocalMux
    port map (
            O => \N__52455\,
            I => \N__52449\
        );

    \I__12706\ : Odrv4
    port map (
            O => \N__52452\,
            I => \comm_spi.n14603\
        );

    \I__12705\ : Odrv12
    port map (
            O => \N__52449\,
            I => \comm_spi.n14603\
        );

    \I__12704\ : ClkMux
    port map (
            O => \N__52444\,
            I => \N__52438\
        );

    \I__12703\ : ClkMux
    port map (
            O => \N__52443\,
            I => \N__52434\
        );

    \I__12702\ : ClkMux
    port map (
            O => \N__52442\,
            I => \N__52431\
        );

    \I__12701\ : ClkMux
    port map (
            O => \N__52441\,
            I => \N__52427\
        );

    \I__12700\ : LocalMux
    port map (
            O => \N__52438\,
            I => \N__52421\
        );

    \I__12699\ : ClkMux
    port map (
            O => \N__52437\,
            I => \N__52418\
        );

    \I__12698\ : LocalMux
    port map (
            O => \N__52434\,
            I => \N__52408\
        );

    \I__12697\ : LocalMux
    port map (
            O => \N__52431\,
            I => \N__52408\
        );

    \I__12696\ : ClkMux
    port map (
            O => \N__52430\,
            I => \N__52404\
        );

    \I__12695\ : LocalMux
    port map (
            O => \N__52427\,
            I => \N__52401\
        );

    \I__12694\ : ClkMux
    port map (
            O => \N__52426\,
            I => \N__52398\
        );

    \I__12693\ : ClkMux
    port map (
            O => \N__52425\,
            I => \N__52395\
        );

    \I__12692\ : ClkMux
    port map (
            O => \N__52424\,
            I => \N__52392\
        );

    \I__12691\ : Span4Mux_v
    port map (
            O => \N__52421\,
            I => \N__52386\
        );

    \I__12690\ : LocalMux
    port map (
            O => \N__52418\,
            I => \N__52386\
        );

    \I__12689\ : ClkMux
    port map (
            O => \N__52417\,
            I => \N__52383\
        );

    \I__12688\ : ClkMux
    port map (
            O => \N__52416\,
            I => \N__52380\
        );

    \I__12687\ : ClkMux
    port map (
            O => \N__52415\,
            I => \N__52376\
        );

    \I__12686\ : ClkMux
    port map (
            O => \N__52414\,
            I => \N__52372\
        );

    \I__12685\ : ClkMux
    port map (
            O => \N__52413\,
            I => \N__52369\
        );

    \I__12684\ : Span4Mux_v
    port map (
            O => \N__52408\,
            I => \N__52365\
        );

    \I__12683\ : ClkMux
    port map (
            O => \N__52407\,
            I => \N__52361\
        );

    \I__12682\ : LocalMux
    port map (
            O => \N__52404\,
            I => \N__52353\
        );

    \I__12681\ : Span4Mux_h
    port map (
            O => \N__52401\,
            I => \N__52353\
        );

    \I__12680\ : LocalMux
    port map (
            O => \N__52398\,
            I => \N__52353\
        );

    \I__12679\ : LocalMux
    port map (
            O => \N__52395\,
            I => \N__52348\
        );

    \I__12678\ : LocalMux
    port map (
            O => \N__52392\,
            I => \N__52348\
        );

    \I__12677\ : ClkMux
    port map (
            O => \N__52391\,
            I => \N__52345\
        );

    \I__12676\ : Span4Mux_v
    port map (
            O => \N__52386\,
            I => \N__52340\
        );

    \I__12675\ : LocalMux
    port map (
            O => \N__52383\,
            I => \N__52340\
        );

    \I__12674\ : LocalMux
    port map (
            O => \N__52380\,
            I => \N__52337\
        );

    \I__12673\ : ClkMux
    port map (
            O => \N__52379\,
            I => \N__52334\
        );

    \I__12672\ : LocalMux
    port map (
            O => \N__52376\,
            I => \N__52331\
        );

    \I__12671\ : ClkMux
    port map (
            O => \N__52375\,
            I => \N__52328\
        );

    \I__12670\ : LocalMux
    port map (
            O => \N__52372\,
            I => \N__52323\
        );

    \I__12669\ : LocalMux
    port map (
            O => \N__52369\,
            I => \N__52323\
        );

    \I__12668\ : ClkMux
    port map (
            O => \N__52368\,
            I => \N__52320\
        );

    \I__12667\ : Span4Mux_h
    port map (
            O => \N__52365\,
            I => \N__52316\
        );

    \I__12666\ : ClkMux
    port map (
            O => \N__52364\,
            I => \N__52313\
        );

    \I__12665\ : LocalMux
    port map (
            O => \N__52361\,
            I => \N__52310\
        );

    \I__12664\ : ClkMux
    port map (
            O => \N__52360\,
            I => \N__52307\
        );

    \I__12663\ : Span4Mux_v
    port map (
            O => \N__52353\,
            I => \N__52304\
        );

    \I__12662\ : Span4Mux_h
    port map (
            O => \N__52348\,
            I => \N__52293\
        );

    \I__12661\ : LocalMux
    port map (
            O => \N__52345\,
            I => \N__52293\
        );

    \I__12660\ : Span4Mux_h
    port map (
            O => \N__52340\,
            I => \N__52293\
        );

    \I__12659\ : Span4Mux_v
    port map (
            O => \N__52337\,
            I => \N__52293\
        );

    \I__12658\ : LocalMux
    port map (
            O => \N__52334\,
            I => \N__52293\
        );

    \I__12657\ : Span4Mux_v
    port map (
            O => \N__52331\,
            I => \N__52288\
        );

    \I__12656\ : LocalMux
    port map (
            O => \N__52328\,
            I => \N__52288\
        );

    \I__12655\ : Span4Mux_v
    port map (
            O => \N__52323\,
            I => \N__52283\
        );

    \I__12654\ : LocalMux
    port map (
            O => \N__52320\,
            I => \N__52283\
        );

    \I__12653\ : ClkMux
    port map (
            O => \N__52319\,
            I => \N__52280\
        );

    \I__12652\ : Span4Mux_v
    port map (
            O => \N__52316\,
            I => \N__52277\
        );

    \I__12651\ : LocalMux
    port map (
            O => \N__52313\,
            I => \N__52274\
        );

    \I__12650\ : Span4Mux_h
    port map (
            O => \N__52310\,
            I => \N__52267\
        );

    \I__12649\ : LocalMux
    port map (
            O => \N__52307\,
            I => \N__52267\
        );

    \I__12648\ : Span4Mux_h
    port map (
            O => \N__52304\,
            I => \N__52267\
        );

    \I__12647\ : Span4Mux_v
    port map (
            O => \N__52293\,
            I => \N__52264\
        );

    \I__12646\ : Span4Mux_h
    port map (
            O => \N__52288\,
            I => \N__52257\
        );

    \I__12645\ : Span4Mux_h
    port map (
            O => \N__52283\,
            I => \N__52257\
        );

    \I__12644\ : LocalMux
    port map (
            O => \N__52280\,
            I => \N__52257\
        );

    \I__12643\ : Odrv4
    port map (
            O => \N__52277\,
            I => \comm_spi.iclk\
        );

    \I__12642\ : Odrv12
    port map (
            O => \N__52274\,
            I => \comm_spi.iclk\
        );

    \I__12641\ : Odrv4
    port map (
            O => \N__52267\,
            I => \comm_spi.iclk\
        );

    \I__12640\ : Odrv4
    port map (
            O => \N__52264\,
            I => \comm_spi.iclk\
        );

    \I__12639\ : Odrv4
    port map (
            O => \N__52257\,
            I => \comm_spi.iclk\
        );

    \I__12638\ : InMux
    port map (
            O => \N__52246\,
            I => \N__52243\
        );

    \I__12637\ : LocalMux
    port map (
            O => \N__52243\,
            I => \N__52240\
        );

    \I__12636\ : Span4Mux_h
    port map (
            O => \N__52240\,
            I => \N__52237\
        );

    \I__12635\ : Odrv4
    port map (
            O => \N__52237\,
            I => n20863
        );

    \I__12634\ : InMux
    port map (
            O => \N__52234\,
            I => \N__52229\
        );

    \I__12633\ : InMux
    port map (
            O => \N__52233\,
            I => \N__52226\
        );

    \I__12632\ : CascadeMux
    port map (
            O => \N__52232\,
            I => \N__52223\
        );

    \I__12631\ : LocalMux
    port map (
            O => \N__52229\,
            I => \N__52220\
        );

    \I__12630\ : LocalMux
    port map (
            O => \N__52226\,
            I => \N__52217\
        );

    \I__12629\ : InMux
    port map (
            O => \N__52223\,
            I => \N__52214\
        );

    \I__12628\ : Span4Mux_h
    port map (
            O => \N__52220\,
            I => \N__52211\
        );

    \I__12627\ : Span4Mux_h
    port map (
            O => \N__52217\,
            I => \N__52208\
        );

    \I__12626\ : LocalMux
    port map (
            O => \N__52214\,
            I => \N__52205\
        );

    \I__12625\ : Odrv4
    port map (
            O => \N__52211\,
            I => n14514
        );

    \I__12624\ : Odrv4
    port map (
            O => \N__52208\,
            I => n14514
        );

    \I__12623\ : Odrv4
    port map (
            O => \N__52205\,
            I => n14514
        );

    \I__12622\ : CascadeMux
    port map (
            O => \N__52198\,
            I => \n21658_cascade_\
        );

    \I__12621\ : InMux
    port map (
            O => \N__52195\,
            I => \N__52186\
        );

    \I__12620\ : CascadeMux
    port map (
            O => \N__52194\,
            I => \N__52182\
        );

    \I__12619\ : CascadeMux
    port map (
            O => \N__52193\,
            I => \N__52178\
        );

    \I__12618\ : CascadeMux
    port map (
            O => \N__52192\,
            I => \N__52163\
        );

    \I__12617\ : InMux
    port map (
            O => \N__52191\,
            I => \N__52151\
        );

    \I__12616\ : InMux
    port map (
            O => \N__52190\,
            I => \N__52151\
        );

    \I__12615\ : InMux
    port map (
            O => \N__52189\,
            I => \N__52151\
        );

    \I__12614\ : LocalMux
    port map (
            O => \N__52186\,
            I => \N__52148\
        );

    \I__12613\ : InMux
    port map (
            O => \N__52185\,
            I => \N__52140\
        );

    \I__12612\ : InMux
    port map (
            O => \N__52182\,
            I => \N__52140\
        );

    \I__12611\ : InMux
    port map (
            O => \N__52181\,
            I => \N__52140\
        );

    \I__12610\ : InMux
    port map (
            O => \N__52178\,
            I => \N__52135\
        );

    \I__12609\ : InMux
    port map (
            O => \N__52177\,
            I => \N__52135\
        );

    \I__12608\ : InMux
    port map (
            O => \N__52176\,
            I => \N__52132\
        );

    \I__12607\ : InMux
    port map (
            O => \N__52175\,
            I => \N__52125\
        );

    \I__12606\ : InMux
    port map (
            O => \N__52174\,
            I => \N__52125\
        );

    \I__12605\ : InMux
    port map (
            O => \N__52173\,
            I => \N__52125\
        );

    \I__12604\ : CascadeMux
    port map (
            O => \N__52172\,
            I => \N__52120\
        );

    \I__12603\ : CascadeMux
    port map (
            O => \N__52171\,
            I => \N__52117\
        );

    \I__12602\ : CascadeMux
    port map (
            O => \N__52170\,
            I => \N__52114\
        );

    \I__12601\ : InMux
    port map (
            O => \N__52169\,
            I => \N__52105\
        );

    \I__12600\ : InMux
    port map (
            O => \N__52168\,
            I => \N__52102\
        );

    \I__12599\ : CascadeMux
    port map (
            O => \N__52167\,
            I => \N__52099\
        );

    \I__12598\ : CascadeMux
    port map (
            O => \N__52166\,
            I => \N__52096\
        );

    \I__12597\ : InMux
    port map (
            O => \N__52163\,
            I => \N__52093\
        );

    \I__12596\ : InMux
    port map (
            O => \N__52162\,
            I => \N__52088\
        );

    \I__12595\ : CascadeMux
    port map (
            O => \N__52161\,
            I => \N__52084\
        );

    \I__12594\ : CascadeMux
    port map (
            O => \N__52160\,
            I => \N__52081\
        );

    \I__12593\ : CascadeMux
    port map (
            O => \N__52159\,
            I => \N__52078\
        );

    \I__12592\ : CascadeMux
    port map (
            O => \N__52158\,
            I => \N__52074\
        );

    \I__12591\ : LocalMux
    port map (
            O => \N__52151\,
            I => \N__52069\
        );

    \I__12590\ : Span4Mux_v
    port map (
            O => \N__52148\,
            I => \N__52069\
        );

    \I__12589\ : CascadeMux
    port map (
            O => \N__52147\,
            I => \N__52066\
        );

    \I__12588\ : LocalMux
    port map (
            O => \N__52140\,
            I => \N__52050\
        );

    \I__12587\ : LocalMux
    port map (
            O => \N__52135\,
            I => \N__52050\
        );

    \I__12586\ : LocalMux
    port map (
            O => \N__52132\,
            I => \N__52050\
        );

    \I__12585\ : LocalMux
    port map (
            O => \N__52125\,
            I => \N__52050\
        );

    \I__12584\ : CascadeMux
    port map (
            O => \N__52124\,
            I => \N__52047\
        );

    \I__12583\ : CascadeMux
    port map (
            O => \N__52123\,
            I => \N__52044\
        );

    \I__12582\ : InMux
    port map (
            O => \N__52120\,
            I => \N__52037\
        );

    \I__12581\ : InMux
    port map (
            O => \N__52117\,
            I => \N__52037\
        );

    \I__12580\ : InMux
    port map (
            O => \N__52114\,
            I => \N__52034\
        );

    \I__12579\ : CascadeMux
    port map (
            O => \N__52113\,
            I => \N__52030\
        );

    \I__12578\ : InMux
    port map (
            O => \N__52112\,
            I => \N__52027\
        );

    \I__12577\ : InMux
    port map (
            O => \N__52111\,
            I => \N__52024\
        );

    \I__12576\ : InMux
    port map (
            O => \N__52110\,
            I => \N__52017\
        );

    \I__12575\ : InMux
    port map (
            O => \N__52109\,
            I => \N__52017\
        );

    \I__12574\ : InMux
    port map (
            O => \N__52108\,
            I => \N__52017\
        );

    \I__12573\ : LocalMux
    port map (
            O => \N__52105\,
            I => \N__52012\
        );

    \I__12572\ : LocalMux
    port map (
            O => \N__52102\,
            I => \N__52012\
        );

    \I__12571\ : InMux
    port map (
            O => \N__52099\,
            I => \N__52007\
        );

    \I__12570\ : InMux
    port map (
            O => \N__52096\,
            I => \N__52007\
        );

    \I__12569\ : LocalMux
    port map (
            O => \N__52093\,
            I => \N__52004\
        );

    \I__12568\ : CascadeMux
    port map (
            O => \N__52092\,
            I => \N__52001\
        );

    \I__12567\ : CascadeMux
    port map (
            O => \N__52091\,
            I => \N__51998\
        );

    \I__12566\ : LocalMux
    port map (
            O => \N__52088\,
            I => \N__51995\
        );

    \I__12565\ : InMux
    port map (
            O => \N__52087\,
            I => \N__51986\
        );

    \I__12564\ : InMux
    port map (
            O => \N__52084\,
            I => \N__51986\
        );

    \I__12563\ : InMux
    port map (
            O => \N__52081\,
            I => \N__51986\
        );

    \I__12562\ : InMux
    port map (
            O => \N__52078\,
            I => \N__51986\
        );

    \I__12561\ : CascadeMux
    port map (
            O => \N__52077\,
            I => \N__51980\
        );

    \I__12560\ : InMux
    port map (
            O => \N__52074\,
            I => \N__51971\
        );

    \I__12559\ : Span4Mux_h
    port map (
            O => \N__52069\,
            I => \N__51968\
        );

    \I__12558\ : InMux
    port map (
            O => \N__52066\,
            I => \N__51963\
        );

    \I__12557\ : InMux
    port map (
            O => \N__52065\,
            I => \N__51963\
        );

    \I__12556\ : InMux
    port map (
            O => \N__52064\,
            I => \N__51958\
        );

    \I__12555\ : InMux
    port map (
            O => \N__52063\,
            I => \N__51958\
        );

    \I__12554\ : CascadeMux
    port map (
            O => \N__52062\,
            I => \N__51955\
        );

    \I__12553\ : CascadeMux
    port map (
            O => \N__52061\,
            I => \N__51952\
        );

    \I__12552\ : InMux
    port map (
            O => \N__52060\,
            I => \N__51945\
        );

    \I__12551\ : InMux
    port map (
            O => \N__52059\,
            I => \N__51945\
        );

    \I__12550\ : Span4Mux_v
    port map (
            O => \N__52050\,
            I => \N__51942\
        );

    \I__12549\ : InMux
    port map (
            O => \N__52047\,
            I => \N__51937\
        );

    \I__12548\ : InMux
    port map (
            O => \N__52044\,
            I => \N__51937\
        );

    \I__12547\ : CascadeMux
    port map (
            O => \N__52043\,
            I => \N__51934\
        );

    \I__12546\ : CascadeMux
    port map (
            O => \N__52042\,
            I => \N__51931\
        );

    \I__12545\ : LocalMux
    port map (
            O => \N__52037\,
            I => \N__51924\
        );

    \I__12544\ : LocalMux
    port map (
            O => \N__52034\,
            I => \N__51924\
        );

    \I__12543\ : CascadeMux
    port map (
            O => \N__52033\,
            I => \N__51921\
        );

    \I__12542\ : InMux
    port map (
            O => \N__52030\,
            I => \N__51916\
        );

    \I__12541\ : LocalMux
    port map (
            O => \N__52027\,
            I => \N__51907\
        );

    \I__12540\ : LocalMux
    port map (
            O => \N__52024\,
            I => \N__51907\
        );

    \I__12539\ : LocalMux
    port map (
            O => \N__52017\,
            I => \N__51907\
        );

    \I__12538\ : Span4Mux_v
    port map (
            O => \N__52012\,
            I => \N__51900\
        );

    \I__12537\ : LocalMux
    port map (
            O => \N__52007\,
            I => \N__51900\
        );

    \I__12536\ : Span4Mux_v
    port map (
            O => \N__52004\,
            I => \N__51900\
        );

    \I__12535\ : InMux
    port map (
            O => \N__52001\,
            I => \N__51895\
        );

    \I__12534\ : InMux
    port map (
            O => \N__51998\,
            I => \N__51895\
        );

    \I__12533\ : Span4Mux_h
    port map (
            O => \N__51995\,
            I => \N__51888\
        );

    \I__12532\ : LocalMux
    port map (
            O => \N__51986\,
            I => \N__51888\
        );

    \I__12531\ : CascadeMux
    port map (
            O => \N__51985\,
            I => \N__51885\
        );

    \I__12530\ : CascadeMux
    port map (
            O => \N__51984\,
            I => \N__51882\
        );

    \I__12529\ : InMux
    port map (
            O => \N__51983\,
            I => \N__51878\
        );

    \I__12528\ : InMux
    port map (
            O => \N__51980\,
            I => \N__51873\
        );

    \I__12527\ : InMux
    port map (
            O => \N__51979\,
            I => \N__51873\
        );

    \I__12526\ : InMux
    port map (
            O => \N__51978\,
            I => \N__51870\
        );

    \I__12525\ : InMux
    port map (
            O => \N__51977\,
            I => \N__51861\
        );

    \I__12524\ : InMux
    port map (
            O => \N__51976\,
            I => \N__51861\
        );

    \I__12523\ : InMux
    port map (
            O => \N__51975\,
            I => \N__51861\
        );

    \I__12522\ : InMux
    port map (
            O => \N__51974\,
            I => \N__51861\
        );

    \I__12521\ : LocalMux
    port map (
            O => \N__51971\,
            I => \N__51852\
        );

    \I__12520\ : Span4Mux_h
    port map (
            O => \N__51968\,
            I => \N__51852\
        );

    \I__12519\ : LocalMux
    port map (
            O => \N__51963\,
            I => \N__51852\
        );

    \I__12518\ : LocalMux
    port map (
            O => \N__51958\,
            I => \N__51852\
        );

    \I__12517\ : InMux
    port map (
            O => \N__51955\,
            I => \N__51849\
        );

    \I__12516\ : InMux
    port map (
            O => \N__51952\,
            I => \N__51842\
        );

    \I__12515\ : InMux
    port map (
            O => \N__51951\,
            I => \N__51842\
        );

    \I__12514\ : InMux
    port map (
            O => \N__51950\,
            I => \N__51842\
        );

    \I__12513\ : LocalMux
    port map (
            O => \N__51945\,
            I => \N__51835\
        );

    \I__12512\ : Span4Mux_h
    port map (
            O => \N__51942\,
            I => \N__51835\
        );

    \I__12511\ : LocalMux
    port map (
            O => \N__51937\,
            I => \N__51835\
        );

    \I__12510\ : InMux
    port map (
            O => \N__51934\,
            I => \N__51826\
        );

    \I__12509\ : InMux
    port map (
            O => \N__51931\,
            I => \N__51826\
        );

    \I__12508\ : InMux
    port map (
            O => \N__51930\,
            I => \N__51826\
        );

    \I__12507\ : InMux
    port map (
            O => \N__51929\,
            I => \N__51826\
        );

    \I__12506\ : Span4Mux_h
    port map (
            O => \N__51924\,
            I => \N__51823\
        );

    \I__12505\ : InMux
    port map (
            O => \N__51921\,
            I => \N__51818\
        );

    \I__12504\ : InMux
    port map (
            O => \N__51920\,
            I => \N__51818\
        );

    \I__12503\ : InMux
    port map (
            O => \N__51919\,
            I => \N__51815\
        );

    \I__12502\ : LocalMux
    port map (
            O => \N__51916\,
            I => \N__51812\
        );

    \I__12501\ : InMux
    port map (
            O => \N__51915\,
            I => \N__51807\
        );

    \I__12500\ : InMux
    port map (
            O => \N__51914\,
            I => \N__51807\
        );

    \I__12499\ : Span4Mux_v
    port map (
            O => \N__51907\,
            I => \N__51800\
        );

    \I__12498\ : Span4Mux_h
    port map (
            O => \N__51900\,
            I => \N__51800\
        );

    \I__12497\ : LocalMux
    port map (
            O => \N__51895\,
            I => \N__51800\
        );

    \I__12496\ : InMux
    port map (
            O => \N__51894\,
            I => \N__51795\
        );

    \I__12495\ : InMux
    port map (
            O => \N__51893\,
            I => \N__51795\
        );

    \I__12494\ : Span4Mux_v
    port map (
            O => \N__51888\,
            I => \N__51792\
        );

    \I__12493\ : InMux
    port map (
            O => \N__51885\,
            I => \N__51787\
        );

    \I__12492\ : InMux
    port map (
            O => \N__51882\,
            I => \N__51787\
        );

    \I__12491\ : InMux
    port map (
            O => \N__51881\,
            I => \N__51783\
        );

    \I__12490\ : LocalMux
    port map (
            O => \N__51878\,
            I => \N__51763\
        );

    \I__12489\ : LocalMux
    port map (
            O => \N__51873\,
            I => \N__51763\
        );

    \I__12488\ : LocalMux
    port map (
            O => \N__51870\,
            I => \N__51763\
        );

    \I__12487\ : LocalMux
    port map (
            O => \N__51861\,
            I => \N__51763\
        );

    \I__12486\ : Span4Mux_v
    port map (
            O => \N__51852\,
            I => \N__51763\
        );

    \I__12485\ : LocalMux
    port map (
            O => \N__51849\,
            I => \N__51763\
        );

    \I__12484\ : LocalMux
    port map (
            O => \N__51842\,
            I => \N__51763\
        );

    \I__12483\ : Span4Mux_v
    port map (
            O => \N__51835\,
            I => \N__51763\
        );

    \I__12482\ : LocalMux
    port map (
            O => \N__51826\,
            I => \N__51763\
        );

    \I__12481\ : Span4Mux_h
    port map (
            O => \N__51823\,
            I => \N__51758\
        );

    \I__12480\ : LocalMux
    port map (
            O => \N__51818\,
            I => \N__51758\
        );

    \I__12479\ : LocalMux
    port map (
            O => \N__51815\,
            I => \N__51755\
        );

    \I__12478\ : Span4Mux_h
    port map (
            O => \N__51812\,
            I => \N__51752\
        );

    \I__12477\ : LocalMux
    port map (
            O => \N__51807\,
            I => \N__51747\
        );

    \I__12476\ : Span4Mux_h
    port map (
            O => \N__51800\,
            I => \N__51747\
        );

    \I__12475\ : LocalMux
    port map (
            O => \N__51795\,
            I => \N__51740\
        );

    \I__12474\ : Span4Mux_h
    port map (
            O => \N__51792\,
            I => \N__51740\
        );

    \I__12473\ : LocalMux
    port map (
            O => \N__51787\,
            I => \N__51740\
        );

    \I__12472\ : InMux
    port map (
            O => \N__51786\,
            I => \N__51737\
        );

    \I__12471\ : LocalMux
    port map (
            O => \N__51783\,
            I => \N__51734\
        );

    \I__12470\ : InMux
    port map (
            O => \N__51782\,
            I => \N__51731\
        );

    \I__12469\ : Span4Mux_v
    port map (
            O => \N__51763\,
            I => \N__51728\
        );

    \I__12468\ : Span4Mux_h
    port map (
            O => \N__51758\,
            I => \N__51725\
        );

    \I__12467\ : Span4Mux_v
    port map (
            O => \N__51755\,
            I => \N__51716\
        );

    \I__12466\ : Span4Mux_v
    port map (
            O => \N__51752\,
            I => \N__51716\
        );

    \I__12465\ : Span4Mux_h
    port map (
            O => \N__51747\,
            I => \N__51716\
        );

    \I__12464\ : Span4Mux_h
    port map (
            O => \N__51740\,
            I => \N__51716\
        );

    \I__12463\ : LocalMux
    port map (
            O => \N__51737\,
            I => n9273
        );

    \I__12462\ : Odrv4
    port map (
            O => \N__51734\,
            I => n9273
        );

    \I__12461\ : LocalMux
    port map (
            O => \N__51731\,
            I => n9273
        );

    \I__12460\ : Odrv4
    port map (
            O => \N__51728\,
            I => n9273
        );

    \I__12459\ : Odrv4
    port map (
            O => \N__51725\,
            I => n9273
        );

    \I__12458\ : Odrv4
    port map (
            O => \N__51716\,
            I => n9273
        );

    \I__12457\ : CascadeMux
    port map (
            O => \N__51703\,
            I => \n20865_cascade_\
        );

    \I__12456\ : CEMux
    port map (
            O => \N__51700\,
            I => \N__51697\
        );

    \I__12455\ : LocalMux
    port map (
            O => \N__51697\,
            I => \N__51694\
        );

    \I__12454\ : Span4Mux_v
    port map (
            O => \N__51694\,
            I => \N__51691\
        );

    \I__12453\ : Span4Mux_h
    port map (
            O => \N__51691\,
            I => \N__51688\
        );

    \I__12452\ : Odrv4
    port map (
            O => \N__51688\,
            I => n20536
        );

    \I__12451\ : InMux
    port map (
            O => \N__51685\,
            I => \N__51681\
        );

    \I__12450\ : InMux
    port map (
            O => \N__51684\,
            I => \N__51678\
        );

    \I__12449\ : LocalMux
    port map (
            O => \N__51681\,
            I => \N__51674\
        );

    \I__12448\ : LocalMux
    port map (
            O => \N__51678\,
            I => \N__51671\
        );

    \I__12447\ : InMux
    port map (
            O => \N__51677\,
            I => \N__51668\
        );

    \I__12446\ : Span4Mux_v
    port map (
            O => \N__51674\,
            I => \N__51665\
        );

    \I__12445\ : Span4Mux_v
    port map (
            O => \N__51671\,
            I => \N__51660\
        );

    \I__12444\ : LocalMux
    port map (
            O => \N__51668\,
            I => \N__51660\
        );

    \I__12443\ : Sp12to4
    port map (
            O => \N__51665\,
            I => \N__51656\
        );

    \I__12442\ : Span4Mux_h
    port map (
            O => \N__51660\,
            I => \N__51653\
        );

    \I__12441\ : InMux
    port map (
            O => \N__51659\,
            I => \N__51650\
        );

    \I__12440\ : Odrv12
    port map (
            O => \N__51656\,
            I => n10540
        );

    \I__12439\ : Odrv4
    port map (
            O => \N__51653\,
            I => n10540
        );

    \I__12438\ : LocalMux
    port map (
            O => \N__51650\,
            I => n10540
        );

    \I__12437\ : InMux
    port map (
            O => \N__51643\,
            I => \N__51633\
        );

    \I__12436\ : InMux
    port map (
            O => \N__51642\,
            I => \N__51633\
        );

    \I__12435\ : InMux
    port map (
            O => \N__51641\,
            I => \N__51610\
        );

    \I__12434\ : InMux
    port map (
            O => \N__51640\,
            I => \N__51610\
        );

    \I__12433\ : InMux
    port map (
            O => \N__51639\,
            I => \N__51610\
        );

    \I__12432\ : InMux
    port map (
            O => \N__51638\,
            I => \N__51610\
        );

    \I__12431\ : LocalMux
    port map (
            O => \N__51633\,
            I => \N__51607\
        );

    \I__12430\ : InMux
    port map (
            O => \N__51632\,
            I => \N__51601\
        );

    \I__12429\ : InMux
    port map (
            O => \N__51631\,
            I => \N__51592\
        );

    \I__12428\ : InMux
    port map (
            O => \N__51630\,
            I => \N__51592\
        );

    \I__12427\ : InMux
    port map (
            O => \N__51629\,
            I => \N__51592\
        );

    \I__12426\ : InMux
    port map (
            O => \N__51628\,
            I => \N__51592\
        );

    \I__12425\ : InMux
    port map (
            O => \N__51627\,
            I => \N__51583\
        );

    \I__12424\ : InMux
    port map (
            O => \N__51626\,
            I => \N__51583\
        );

    \I__12423\ : InMux
    port map (
            O => \N__51625\,
            I => \N__51583\
        );

    \I__12422\ : InMux
    port map (
            O => \N__51624\,
            I => \N__51583\
        );

    \I__12421\ : InMux
    port map (
            O => \N__51623\,
            I => \N__51580\
        );

    \I__12420\ : InMux
    port map (
            O => \N__51622\,
            I => \N__51570\
        );

    \I__12419\ : InMux
    port map (
            O => \N__51621\,
            I => \N__51570\
        );

    \I__12418\ : InMux
    port map (
            O => \N__51620\,
            I => \N__51570\
        );

    \I__12417\ : CascadeMux
    port map (
            O => \N__51619\,
            I => \N__51567\
        );

    \I__12416\ : LocalMux
    port map (
            O => \N__51610\,
            I => \N__51564\
        );

    \I__12415\ : Span4Mux_v
    port map (
            O => \N__51607\,
            I => \N__51561\
        );

    \I__12414\ : InMux
    port map (
            O => \N__51606\,
            I => \N__51554\
        );

    \I__12413\ : InMux
    port map (
            O => \N__51605\,
            I => \N__51554\
        );

    \I__12412\ : InMux
    port map (
            O => \N__51604\,
            I => \N__51554\
        );

    \I__12411\ : LocalMux
    port map (
            O => \N__51601\,
            I => \N__51551\
        );

    \I__12410\ : LocalMux
    port map (
            O => \N__51592\,
            I => \N__51544\
        );

    \I__12409\ : LocalMux
    port map (
            O => \N__51583\,
            I => \N__51544\
        );

    \I__12408\ : LocalMux
    port map (
            O => \N__51580\,
            I => \N__51544\
        );

    \I__12407\ : InMux
    port map (
            O => \N__51579\,
            I => \N__51541\
        );

    \I__12406\ : InMux
    port map (
            O => \N__51578\,
            I => \N__51538\
        );

    \I__12405\ : CascadeMux
    port map (
            O => \N__51577\,
            I => \N__51534\
        );

    \I__12404\ : LocalMux
    port map (
            O => \N__51570\,
            I => \N__51530\
        );

    \I__12403\ : InMux
    port map (
            O => \N__51567\,
            I => \N__51526\
        );

    \I__12402\ : Span4Mux_v
    port map (
            O => \N__51564\,
            I => \N__51519\
        );

    \I__12401\ : Span4Mux_h
    port map (
            O => \N__51561\,
            I => \N__51519\
        );

    \I__12400\ : LocalMux
    port map (
            O => \N__51554\,
            I => \N__51519\
        );

    \I__12399\ : Span4Mux_v
    port map (
            O => \N__51551\,
            I => \N__51510\
        );

    \I__12398\ : Span4Mux_v
    port map (
            O => \N__51544\,
            I => \N__51510\
        );

    \I__12397\ : LocalMux
    port map (
            O => \N__51541\,
            I => \N__51505\
        );

    \I__12396\ : LocalMux
    port map (
            O => \N__51538\,
            I => \N__51505\
        );

    \I__12395\ : InMux
    port map (
            O => \N__51537\,
            I => \N__51498\
        );

    \I__12394\ : InMux
    port map (
            O => \N__51534\,
            I => \N__51498\
        );

    \I__12393\ : InMux
    port map (
            O => \N__51533\,
            I => \N__51498\
        );

    \I__12392\ : Span12Mux_v
    port map (
            O => \N__51530\,
            I => \N__51495\
        );

    \I__12391\ : InMux
    port map (
            O => \N__51529\,
            I => \N__51492\
        );

    \I__12390\ : LocalMux
    port map (
            O => \N__51526\,
            I => \N__51487\
        );

    \I__12389\ : Span4Mux_h
    port map (
            O => \N__51519\,
            I => \N__51487\
        );

    \I__12388\ : InMux
    port map (
            O => \N__51518\,
            I => \N__51478\
        );

    \I__12387\ : InMux
    port map (
            O => \N__51517\,
            I => \N__51478\
        );

    \I__12386\ : InMux
    port map (
            O => \N__51516\,
            I => \N__51478\
        );

    \I__12385\ : InMux
    port map (
            O => \N__51515\,
            I => \N__51478\
        );

    \I__12384\ : Span4Mux_h
    port map (
            O => \N__51510\,
            I => \N__51473\
        );

    \I__12383\ : Span4Mux_v
    port map (
            O => \N__51505\,
            I => \N__51473\
        );

    \I__12382\ : LocalMux
    port map (
            O => \N__51498\,
            I => comm_index_0
        );

    \I__12381\ : Odrv12
    port map (
            O => \N__51495\,
            I => comm_index_0
        );

    \I__12380\ : LocalMux
    port map (
            O => \N__51492\,
            I => comm_index_0
        );

    \I__12379\ : Odrv4
    port map (
            O => \N__51487\,
            I => comm_index_0
        );

    \I__12378\ : LocalMux
    port map (
            O => \N__51478\,
            I => comm_index_0
        );

    \I__12377\ : Odrv4
    port map (
            O => \N__51473\,
            I => comm_index_0
        );

    \I__12376\ : InMux
    port map (
            O => \N__51460\,
            I => \N__51457\
        );

    \I__12375\ : LocalMux
    port map (
            O => \N__51457\,
            I => n20563
        );

    \I__12374\ : InMux
    port map (
            O => \N__51454\,
            I => \N__51451\
        );

    \I__12373\ : LocalMux
    port map (
            O => \N__51451\,
            I => \N__51448\
        );

    \I__12372\ : Span4Mux_h
    port map (
            O => \N__51448\,
            I => \N__51445\
        );

    \I__12371\ : Odrv4
    port map (
            O => \N__51445\,
            I => n12_adj_1585
        );

    \I__12370\ : InMux
    port map (
            O => \N__51442\,
            I => \N__51439\
        );

    \I__12369\ : LocalMux
    port map (
            O => \N__51439\,
            I => \N__51435\
        );

    \I__12368\ : CascadeMux
    port map (
            O => \N__51438\,
            I => \N__51432\
        );

    \I__12367\ : Span4Mux_v
    port map (
            O => \N__51435\,
            I => \N__51425\
        );

    \I__12366\ : InMux
    port map (
            O => \N__51432\,
            I => \N__51420\
        );

    \I__12365\ : InMux
    port map (
            O => \N__51431\,
            I => \N__51420\
        );

    \I__12364\ : CascadeMux
    port map (
            O => \N__51430\,
            I => \N__51417\
        );

    \I__12363\ : CascadeMux
    port map (
            O => \N__51429\,
            I => \N__51414\
        );

    \I__12362\ : InMux
    port map (
            O => \N__51428\,
            I => \N__51411\
        );

    \I__12361\ : Span4Mux_v
    port map (
            O => \N__51425\,
            I => \N__51406\
        );

    \I__12360\ : LocalMux
    port map (
            O => \N__51420\,
            I => \N__51406\
        );

    \I__12359\ : InMux
    port map (
            O => \N__51417\,
            I => \N__51403\
        );

    \I__12358\ : InMux
    port map (
            O => \N__51414\,
            I => \N__51400\
        );

    \I__12357\ : LocalMux
    port map (
            O => \N__51411\,
            I => \N__51397\
        );

    \I__12356\ : Span4Mux_h
    port map (
            O => \N__51406\,
            I => \N__51394\
        );

    \I__12355\ : LocalMux
    port map (
            O => \N__51403\,
            I => \N__51391\
        );

    \I__12354\ : LocalMux
    port map (
            O => \N__51400\,
            I => \N__51386\
        );

    \I__12353\ : Span4Mux_h
    port map (
            O => \N__51397\,
            I => \N__51386\
        );

    \I__12352\ : Span4Mux_h
    port map (
            O => \N__51394\,
            I => \N__51383\
        );

    \I__12351\ : Odrv12
    port map (
            O => \N__51391\,
            I => comm_buf_1_6
        );

    \I__12350\ : Odrv4
    port map (
            O => \N__51386\,
            I => comm_buf_1_6
        );

    \I__12349\ : Odrv4
    port map (
            O => \N__51383\,
            I => comm_buf_1_6
        );

    \I__12348\ : InMux
    port map (
            O => \N__51376\,
            I => \N__51372\
        );

    \I__12347\ : InMux
    port map (
            O => \N__51375\,
            I => \N__51369\
        );

    \I__12346\ : LocalMux
    port map (
            O => \N__51372\,
            I => \N__51364\
        );

    \I__12345\ : LocalMux
    port map (
            O => \N__51369\,
            I => \N__51364\
        );

    \I__12344\ : Span12Mux_h
    port map (
            O => \N__51364\,
            I => \N__51361\
        );

    \I__12343\ : Odrv12
    port map (
            O => \N__51361\,
            I => n14_adj_1526
        );

    \I__12342\ : InMux
    port map (
            O => \N__51358\,
            I => \N__51355\
        );

    \I__12341\ : LocalMux
    port map (
            O => \N__51355\,
            I => \N__51352\
        );

    \I__12340\ : Span4Mux_v
    port map (
            O => \N__51352\,
            I => \N__51349\
        );

    \I__12339\ : Span4Mux_v
    port map (
            O => \N__51349\,
            I => \N__51346\
        );

    \I__12338\ : Sp12to4
    port map (
            O => \N__51346\,
            I => \N__51343\
        );

    \I__12337\ : Span12Mux_h
    port map (
            O => \N__51343\,
            I => \N__51339\
        );

    \I__12336\ : InMux
    port map (
            O => \N__51342\,
            I => \N__51336\
        );

    \I__12335\ : Odrv12
    port map (
            O => \N__51339\,
            I => buf_adcdata_vdc_4
        );

    \I__12334\ : LocalMux
    port map (
            O => \N__51336\,
            I => buf_adcdata_vdc_4
        );

    \I__12333\ : InMux
    port map (
            O => \N__51331\,
            I => \N__51327\
        );

    \I__12332\ : InMux
    port map (
            O => \N__51330\,
            I => \N__51323\
        );

    \I__12331\ : LocalMux
    port map (
            O => \N__51327\,
            I => \N__51320\
        );

    \I__12330\ : InMux
    port map (
            O => \N__51326\,
            I => \N__51317\
        );

    \I__12329\ : LocalMux
    port map (
            O => \N__51323\,
            I => buf_adcdata_vac_4
        );

    \I__12328\ : Odrv4
    port map (
            O => \N__51320\,
            I => buf_adcdata_vac_4
        );

    \I__12327\ : LocalMux
    port map (
            O => \N__51317\,
            I => buf_adcdata_vac_4
        );

    \I__12326\ : InMux
    port map (
            O => \N__51310\,
            I => \N__51307\
        );

    \I__12325\ : LocalMux
    port map (
            O => \N__51307\,
            I => \N__51304\
        );

    \I__12324\ : Span12Mux_h
    port map (
            O => \N__51304\,
            I => \N__51301\
        );

    \I__12323\ : Odrv12
    port map (
            O => \N__51301\,
            I => n19_adj_1605
        );

    \I__12322\ : InMux
    port map (
            O => \N__51298\,
            I => \N__51294\
        );

    \I__12321\ : CascadeMux
    port map (
            O => \N__51297\,
            I => \N__51290\
        );

    \I__12320\ : LocalMux
    port map (
            O => \N__51294\,
            I => \N__51287\
        );

    \I__12319\ : InMux
    port map (
            O => \N__51293\,
            I => \N__51279\
        );

    \I__12318\ : InMux
    port map (
            O => \N__51290\,
            I => \N__51276\
        );

    \I__12317\ : Span4Mux_v
    port map (
            O => \N__51287\,
            I => \N__51273\
        );

    \I__12316\ : InMux
    port map (
            O => \N__51286\,
            I => \N__51268\
        );

    \I__12315\ : InMux
    port map (
            O => \N__51285\,
            I => \N__51268\
        );

    \I__12314\ : InMux
    port map (
            O => \N__51284\,
            I => \N__51265\
        );

    \I__12313\ : InMux
    port map (
            O => \N__51283\,
            I => \N__51254\
        );

    \I__12312\ : InMux
    port map (
            O => \N__51282\,
            I => \N__51254\
        );

    \I__12311\ : LocalMux
    port map (
            O => \N__51279\,
            I => \N__51251\
        );

    \I__12310\ : LocalMux
    port map (
            O => \N__51276\,
            I => \N__51244\
        );

    \I__12309\ : Span4Mux_h
    port map (
            O => \N__51273\,
            I => \N__51244\
        );

    \I__12308\ : LocalMux
    port map (
            O => \N__51268\,
            I => \N__51244\
        );

    \I__12307\ : LocalMux
    port map (
            O => \N__51265\,
            I => \N__51241\
        );

    \I__12306\ : CascadeMux
    port map (
            O => \N__51264\,
            I => \N__51235\
        );

    \I__12305\ : CascadeMux
    port map (
            O => \N__51263\,
            I => \N__51231\
        );

    \I__12304\ : InMux
    port map (
            O => \N__51262\,
            I => \N__51222\
        );

    \I__12303\ : CascadeMux
    port map (
            O => \N__51261\,
            I => \N__51214\
        );

    \I__12302\ : CascadeMux
    port map (
            O => \N__51260\,
            I => \N__51211\
        );

    \I__12301\ : CascadeMux
    port map (
            O => \N__51259\,
            I => \N__51201\
        );

    \I__12300\ : LocalMux
    port map (
            O => \N__51254\,
            I => \N__51193\
        );

    \I__12299\ : Span4Mux_v
    port map (
            O => \N__51251\,
            I => \N__51186\
        );

    \I__12298\ : Span4Mux_v
    port map (
            O => \N__51244\,
            I => \N__51186\
        );

    \I__12297\ : Span4Mux_h
    port map (
            O => \N__51241\,
            I => \N__51186\
        );

    \I__12296\ : InMux
    port map (
            O => \N__51240\,
            I => \N__51181\
        );

    \I__12295\ : InMux
    port map (
            O => \N__51239\,
            I => \N__51181\
        );

    \I__12294\ : InMux
    port map (
            O => \N__51238\,
            I => \N__51178\
        );

    \I__12293\ : InMux
    port map (
            O => \N__51235\,
            I => \N__51169\
        );

    \I__12292\ : InMux
    port map (
            O => \N__51234\,
            I => \N__51169\
        );

    \I__12291\ : InMux
    port map (
            O => \N__51231\,
            I => \N__51169\
        );

    \I__12290\ : InMux
    port map (
            O => \N__51230\,
            I => \N__51169\
        );

    \I__12289\ : InMux
    port map (
            O => \N__51229\,
            I => \N__51166\
        );

    \I__12288\ : InMux
    port map (
            O => \N__51228\,
            I => \N__51163\
        );

    \I__12287\ : InMux
    port map (
            O => \N__51227\,
            I => \N__51156\
        );

    \I__12286\ : InMux
    port map (
            O => \N__51226\,
            I => \N__51156\
        );

    \I__12285\ : InMux
    port map (
            O => \N__51225\,
            I => \N__51156\
        );

    \I__12284\ : LocalMux
    port map (
            O => \N__51222\,
            I => \N__51153\
        );

    \I__12283\ : InMux
    port map (
            O => \N__51221\,
            I => \N__51150\
        );

    \I__12282\ : InMux
    port map (
            O => \N__51220\,
            I => \N__51143\
        );

    \I__12281\ : InMux
    port map (
            O => \N__51219\,
            I => \N__51143\
        );

    \I__12280\ : InMux
    port map (
            O => \N__51218\,
            I => \N__51143\
        );

    \I__12279\ : InMux
    port map (
            O => \N__51217\,
            I => \N__51134\
        );

    \I__12278\ : InMux
    port map (
            O => \N__51214\,
            I => \N__51134\
        );

    \I__12277\ : InMux
    port map (
            O => \N__51211\,
            I => \N__51134\
        );

    \I__12276\ : InMux
    port map (
            O => \N__51210\,
            I => \N__51134\
        );

    \I__12275\ : InMux
    port map (
            O => \N__51209\,
            I => \N__51129\
        );

    \I__12274\ : InMux
    port map (
            O => \N__51208\,
            I => \N__51129\
        );

    \I__12273\ : InMux
    port map (
            O => \N__51207\,
            I => \N__51126\
        );

    \I__12272\ : InMux
    port map (
            O => \N__51206\,
            I => \N__51123\
        );

    \I__12271\ : InMux
    port map (
            O => \N__51205\,
            I => \N__51118\
        );

    \I__12270\ : InMux
    port map (
            O => \N__51204\,
            I => \N__51118\
        );

    \I__12269\ : InMux
    port map (
            O => \N__51201\,
            I => \N__51115\
        );

    \I__12268\ : InMux
    port map (
            O => \N__51200\,
            I => \N__51112\
        );

    \I__12267\ : CascadeMux
    port map (
            O => \N__51199\,
            I => \N__51107\
        );

    \I__12266\ : InMux
    port map (
            O => \N__51198\,
            I => \N__51101\
        );

    \I__12265\ : InMux
    port map (
            O => \N__51197\,
            I => \N__51096\
        );

    \I__12264\ : InMux
    port map (
            O => \N__51196\,
            I => \N__51096\
        );

    \I__12263\ : Span4Mux_v
    port map (
            O => \N__51193\,
            I => \N__51087\
        );

    \I__12262\ : Span4Mux_h
    port map (
            O => \N__51186\,
            I => \N__51087\
        );

    \I__12261\ : LocalMux
    port map (
            O => \N__51181\,
            I => \N__51087\
        );

    \I__12260\ : LocalMux
    port map (
            O => \N__51178\,
            I => \N__51087\
        );

    \I__12259\ : LocalMux
    port map (
            O => \N__51169\,
            I => \N__51084\
        );

    \I__12258\ : LocalMux
    port map (
            O => \N__51166\,
            I => \N__51075\
        );

    \I__12257\ : LocalMux
    port map (
            O => \N__51163\,
            I => \N__51075\
        );

    \I__12256\ : LocalMux
    port map (
            O => \N__51156\,
            I => \N__51075\
        );

    \I__12255\ : Span4Mux_v
    port map (
            O => \N__51153\,
            I => \N__51075\
        );

    \I__12254\ : LocalMux
    port map (
            O => \N__51150\,
            I => \N__51070\
        );

    \I__12253\ : LocalMux
    port map (
            O => \N__51143\,
            I => \N__51063\
        );

    \I__12252\ : LocalMux
    port map (
            O => \N__51134\,
            I => \N__51063\
        );

    \I__12251\ : LocalMux
    port map (
            O => \N__51129\,
            I => \N__51063\
        );

    \I__12250\ : LocalMux
    port map (
            O => \N__51126\,
            I => \N__51058\
        );

    \I__12249\ : LocalMux
    port map (
            O => \N__51123\,
            I => \N__51049\
        );

    \I__12248\ : LocalMux
    port map (
            O => \N__51118\,
            I => \N__51049\
        );

    \I__12247\ : LocalMux
    port map (
            O => \N__51115\,
            I => \N__51049\
        );

    \I__12246\ : LocalMux
    port map (
            O => \N__51112\,
            I => \N__51049\
        );

    \I__12245\ : InMux
    port map (
            O => \N__51111\,
            I => \N__51044\
        );

    \I__12244\ : InMux
    port map (
            O => \N__51110\,
            I => \N__51044\
        );

    \I__12243\ : InMux
    port map (
            O => \N__51107\,
            I => \N__51041\
        );

    \I__12242\ : InMux
    port map (
            O => \N__51106\,
            I => \N__51038\
        );

    \I__12241\ : InMux
    port map (
            O => \N__51105\,
            I => \N__51033\
        );

    \I__12240\ : InMux
    port map (
            O => \N__51104\,
            I => \N__51033\
        );

    \I__12239\ : LocalMux
    port map (
            O => \N__51101\,
            I => \N__51022\
        );

    \I__12238\ : LocalMux
    port map (
            O => \N__51096\,
            I => \N__51022\
        );

    \I__12237\ : Span4Mux_v
    port map (
            O => \N__51087\,
            I => \N__51022\
        );

    \I__12236\ : Span4Mux_v
    port map (
            O => \N__51084\,
            I => \N__51022\
        );

    \I__12235\ : Span4Mux_v
    port map (
            O => \N__51075\,
            I => \N__51022\
        );

    \I__12234\ : InMux
    port map (
            O => \N__51074\,
            I => \N__51017\
        );

    \I__12233\ : InMux
    port map (
            O => \N__51073\,
            I => \N__51017\
        );

    \I__12232\ : Span4Mux_v
    port map (
            O => \N__51070\,
            I => \N__51014\
        );

    \I__12231\ : Span12Mux_h
    port map (
            O => \N__51063\,
            I => \N__51011\
        );

    \I__12230\ : InMux
    port map (
            O => \N__51062\,
            I => \N__51006\
        );

    \I__12229\ : InMux
    port map (
            O => \N__51061\,
            I => \N__51006\
        );

    \I__12228\ : Span4Mux_h
    port map (
            O => \N__51058\,
            I => \N__51001\
        );

    \I__12227\ : Span4Mux_v
    port map (
            O => \N__51049\,
            I => \N__51001\
        );

    \I__12226\ : LocalMux
    port map (
            O => \N__51044\,
            I => comm_state_2
        );

    \I__12225\ : LocalMux
    port map (
            O => \N__51041\,
            I => comm_state_2
        );

    \I__12224\ : LocalMux
    port map (
            O => \N__51038\,
            I => comm_state_2
        );

    \I__12223\ : LocalMux
    port map (
            O => \N__51033\,
            I => comm_state_2
        );

    \I__12222\ : Odrv4
    port map (
            O => \N__51022\,
            I => comm_state_2
        );

    \I__12221\ : LocalMux
    port map (
            O => \N__51017\,
            I => comm_state_2
        );

    \I__12220\ : Odrv4
    port map (
            O => \N__51014\,
            I => comm_state_2
        );

    \I__12219\ : Odrv12
    port map (
            O => \N__51011\,
            I => comm_state_2
        );

    \I__12218\ : LocalMux
    port map (
            O => \N__51006\,
            I => comm_state_2
        );

    \I__12217\ : Odrv4
    port map (
            O => \N__51001\,
            I => comm_state_2
        );

    \I__12216\ : CascadeMux
    port map (
            O => \N__50980\,
            I => \N__50977\
        );

    \I__12215\ : InMux
    port map (
            O => \N__50977\,
            I => \N__50974\
        );

    \I__12214\ : LocalMux
    port map (
            O => \N__50974\,
            I => \N__50971\
        );

    \I__12213\ : Span4Mux_h
    port map (
            O => \N__50971\,
            I => \N__50968\
        );

    \I__12212\ : Odrv4
    port map (
            O => \N__50968\,
            I => n20734
        );

    \I__12211\ : CascadeMux
    port map (
            O => \N__50965\,
            I => \N__50957\
        );

    \I__12210\ : InMux
    port map (
            O => \N__50964\,
            I => \N__50945\
        );

    \I__12209\ : InMux
    port map (
            O => \N__50963\,
            I => \N__50938\
        );

    \I__12208\ : InMux
    port map (
            O => \N__50962\,
            I => \N__50938\
        );

    \I__12207\ : InMux
    port map (
            O => \N__50961\,
            I => \N__50938\
        );

    \I__12206\ : InMux
    port map (
            O => \N__50960\,
            I => \N__50931\
        );

    \I__12205\ : InMux
    port map (
            O => \N__50957\,
            I => \N__50922\
        );

    \I__12204\ : InMux
    port map (
            O => \N__50956\,
            I => \N__50922\
        );

    \I__12203\ : InMux
    port map (
            O => \N__50955\,
            I => \N__50922\
        );

    \I__12202\ : InMux
    port map (
            O => \N__50954\,
            I => \N__50922\
        );

    \I__12201\ : InMux
    port map (
            O => \N__50953\,
            I => \N__50916\
        );

    \I__12200\ : CascadeMux
    port map (
            O => \N__50952\,
            I => \N__50903\
        );

    \I__12199\ : InMux
    port map (
            O => \N__50951\,
            I => \N__50896\
        );

    \I__12198\ : InMux
    port map (
            O => \N__50950\,
            I => \N__50896\
        );

    \I__12197\ : InMux
    port map (
            O => \N__50949\,
            I => \N__50896\
        );

    \I__12196\ : InMux
    port map (
            O => \N__50948\,
            I => \N__50893\
        );

    \I__12195\ : LocalMux
    port map (
            O => \N__50945\,
            I => \N__50888\
        );

    \I__12194\ : LocalMux
    port map (
            O => \N__50938\,
            I => \N__50888\
        );

    \I__12193\ : CascadeMux
    port map (
            O => \N__50937\,
            I => \N__50885\
        );

    \I__12192\ : InMux
    port map (
            O => \N__50936\,
            I => \N__50877\
        );

    \I__12191\ : InMux
    port map (
            O => \N__50935\,
            I => \N__50872\
        );

    \I__12190\ : InMux
    port map (
            O => \N__50934\,
            I => \N__50872\
        );

    \I__12189\ : LocalMux
    port map (
            O => \N__50931\,
            I => \N__50867\
        );

    \I__12188\ : LocalMux
    port map (
            O => \N__50922\,
            I => \N__50867\
        );

    \I__12187\ : InMux
    port map (
            O => \N__50921\,
            I => \N__50860\
        );

    \I__12186\ : InMux
    port map (
            O => \N__50920\,
            I => \N__50860\
        );

    \I__12185\ : InMux
    port map (
            O => \N__50919\,
            I => \N__50860\
        );

    \I__12184\ : LocalMux
    port map (
            O => \N__50916\,
            I => \N__50857\
        );

    \I__12183\ : InMux
    port map (
            O => \N__50915\,
            I => \N__50852\
        );

    \I__12182\ : InMux
    port map (
            O => \N__50914\,
            I => \N__50849\
        );

    \I__12181\ : InMux
    port map (
            O => \N__50913\,
            I => \N__50844\
        );

    \I__12180\ : InMux
    port map (
            O => \N__50912\,
            I => \N__50844\
        );

    \I__12179\ : InMux
    port map (
            O => \N__50911\,
            I => \N__50841\
        );

    \I__12178\ : CascadeMux
    port map (
            O => \N__50910\,
            I => \N__50838\
        );

    \I__12177\ : CascadeMux
    port map (
            O => \N__50909\,
            I => \N__50831\
        );

    \I__12176\ : InMux
    port map (
            O => \N__50908\,
            I => \N__50825\
        );

    \I__12175\ : InMux
    port map (
            O => \N__50907\,
            I => \N__50825\
        );

    \I__12174\ : InMux
    port map (
            O => \N__50906\,
            I => \N__50822\
        );

    \I__12173\ : InMux
    port map (
            O => \N__50903\,
            I => \N__50818\
        );

    \I__12172\ : LocalMux
    port map (
            O => \N__50896\,
            I => \N__50813\
        );

    \I__12171\ : LocalMux
    port map (
            O => \N__50893\,
            I => \N__50813\
        );

    \I__12170\ : Span4Mux_h
    port map (
            O => \N__50888\,
            I => \N__50810\
        );

    \I__12169\ : InMux
    port map (
            O => \N__50885\,
            I => \N__50805\
        );

    \I__12168\ : InMux
    port map (
            O => \N__50884\,
            I => \N__50805\
        );

    \I__12167\ : InMux
    port map (
            O => \N__50883\,
            I => \N__50802\
        );

    \I__12166\ : InMux
    port map (
            O => \N__50882\,
            I => \N__50798\
        );

    \I__12165\ : InMux
    port map (
            O => \N__50881\,
            I => \N__50793\
        );

    \I__12164\ : InMux
    port map (
            O => \N__50880\,
            I => \N__50793\
        );

    \I__12163\ : LocalMux
    port map (
            O => \N__50877\,
            I => \N__50788\
        );

    \I__12162\ : LocalMux
    port map (
            O => \N__50872\,
            I => \N__50788\
        );

    \I__12161\ : Span4Mux_v
    port map (
            O => \N__50867\,
            I => \N__50781\
        );

    \I__12160\ : LocalMux
    port map (
            O => \N__50860\,
            I => \N__50781\
        );

    \I__12159\ : Span4Mux_v
    port map (
            O => \N__50857\,
            I => \N__50781\
        );

    \I__12158\ : InMux
    port map (
            O => \N__50856\,
            I => \N__50776\
        );

    \I__12157\ : InMux
    port map (
            O => \N__50855\,
            I => \N__50776\
        );

    \I__12156\ : LocalMux
    port map (
            O => \N__50852\,
            I => \N__50771\
        );

    \I__12155\ : LocalMux
    port map (
            O => \N__50849\,
            I => \N__50771\
        );

    \I__12154\ : LocalMux
    port map (
            O => \N__50844\,
            I => \N__50766\
        );

    \I__12153\ : LocalMux
    port map (
            O => \N__50841\,
            I => \N__50766\
        );

    \I__12152\ : InMux
    port map (
            O => \N__50838\,
            I => \N__50763\
        );

    \I__12151\ : CascadeMux
    port map (
            O => \N__50837\,
            I => \N__50760\
        );

    \I__12150\ : CascadeMux
    port map (
            O => \N__50836\,
            I => \N__50756\
        );

    \I__12149\ : CascadeMux
    port map (
            O => \N__50835\,
            I => \N__50753\
        );

    \I__12148\ : CascadeMux
    port map (
            O => \N__50834\,
            I => \N__50750\
        );

    \I__12147\ : InMux
    port map (
            O => \N__50831\,
            I => \N__50741\
        );

    \I__12146\ : InMux
    port map (
            O => \N__50830\,
            I => \N__50741\
        );

    \I__12145\ : LocalMux
    port map (
            O => \N__50825\,
            I => \N__50736\
        );

    \I__12144\ : LocalMux
    port map (
            O => \N__50822\,
            I => \N__50736\
        );

    \I__12143\ : InMux
    port map (
            O => \N__50821\,
            I => \N__50733\
        );

    \I__12142\ : LocalMux
    port map (
            O => \N__50818\,
            I => \N__50730\
        );

    \I__12141\ : Span4Mux_h
    port map (
            O => \N__50813\,
            I => \N__50725\
        );

    \I__12140\ : Span4Mux_v
    port map (
            O => \N__50810\,
            I => \N__50725\
        );

    \I__12139\ : LocalMux
    port map (
            O => \N__50805\,
            I => \N__50718\
        );

    \I__12138\ : LocalMux
    port map (
            O => \N__50802\,
            I => \N__50718\
        );

    \I__12137\ : InMux
    port map (
            O => \N__50801\,
            I => \N__50707\
        );

    \I__12136\ : LocalMux
    port map (
            O => \N__50798\,
            I => \N__50704\
        );

    \I__12135\ : LocalMux
    port map (
            O => \N__50793\,
            I => \N__50695\
        );

    \I__12134\ : Span4Mux_v
    port map (
            O => \N__50788\,
            I => \N__50695\
        );

    \I__12133\ : Span4Mux_h
    port map (
            O => \N__50781\,
            I => \N__50695\
        );

    \I__12132\ : LocalMux
    port map (
            O => \N__50776\,
            I => \N__50695\
        );

    \I__12131\ : Span4Mux_v
    port map (
            O => \N__50771\,
            I => \N__50692\
        );

    \I__12130\ : Sp12to4
    port map (
            O => \N__50766\,
            I => \N__50689\
        );

    \I__12129\ : LocalMux
    port map (
            O => \N__50763\,
            I => \N__50686\
        );

    \I__12128\ : InMux
    port map (
            O => \N__50760\,
            I => \N__50681\
        );

    \I__12127\ : InMux
    port map (
            O => \N__50759\,
            I => \N__50681\
        );

    \I__12126\ : InMux
    port map (
            O => \N__50756\,
            I => \N__50666\
        );

    \I__12125\ : InMux
    port map (
            O => \N__50753\,
            I => \N__50666\
        );

    \I__12124\ : InMux
    port map (
            O => \N__50750\,
            I => \N__50666\
        );

    \I__12123\ : InMux
    port map (
            O => \N__50749\,
            I => \N__50666\
        );

    \I__12122\ : InMux
    port map (
            O => \N__50748\,
            I => \N__50666\
        );

    \I__12121\ : InMux
    port map (
            O => \N__50747\,
            I => \N__50666\
        );

    \I__12120\ : InMux
    port map (
            O => \N__50746\,
            I => \N__50666\
        );

    \I__12119\ : LocalMux
    port map (
            O => \N__50741\,
            I => \N__50663\
        );

    \I__12118\ : Span4Mux_h
    port map (
            O => \N__50736\,
            I => \N__50660\
        );

    \I__12117\ : LocalMux
    port map (
            O => \N__50733\,
            I => \N__50657\
        );

    \I__12116\ : Span4Mux_v
    port map (
            O => \N__50730\,
            I => \N__50652\
        );

    \I__12115\ : Span4Mux_h
    port map (
            O => \N__50725\,
            I => \N__50652\
        );

    \I__12114\ : InMux
    port map (
            O => \N__50724\,
            I => \N__50642\
        );

    \I__12113\ : InMux
    port map (
            O => \N__50723\,
            I => \N__50639\
        );

    \I__12112\ : Span4Mux_h
    port map (
            O => \N__50718\,
            I => \N__50636\
        );

    \I__12111\ : InMux
    port map (
            O => \N__50717\,
            I => \N__50619\
        );

    \I__12110\ : InMux
    port map (
            O => \N__50716\,
            I => \N__50619\
        );

    \I__12109\ : InMux
    port map (
            O => \N__50715\,
            I => \N__50619\
        );

    \I__12108\ : InMux
    port map (
            O => \N__50714\,
            I => \N__50619\
        );

    \I__12107\ : InMux
    port map (
            O => \N__50713\,
            I => \N__50619\
        );

    \I__12106\ : InMux
    port map (
            O => \N__50712\,
            I => \N__50619\
        );

    \I__12105\ : InMux
    port map (
            O => \N__50711\,
            I => \N__50619\
        );

    \I__12104\ : InMux
    port map (
            O => \N__50710\,
            I => \N__50619\
        );

    \I__12103\ : LocalMux
    port map (
            O => \N__50707\,
            I => \N__50614\
        );

    \I__12102\ : Span4Mux_v
    port map (
            O => \N__50704\,
            I => \N__50614\
        );

    \I__12101\ : Span4Mux_v
    port map (
            O => \N__50695\,
            I => \N__50611\
        );

    \I__12100\ : Sp12to4
    port map (
            O => \N__50692\,
            I => \N__50606\
        );

    \I__12099\ : Span12Mux_v
    port map (
            O => \N__50689\,
            I => \N__50606\
        );

    \I__12098\ : Span12Mux_s11_h
    port map (
            O => \N__50686\,
            I => \N__50603\
        );

    \I__12097\ : LocalMux
    port map (
            O => \N__50681\,
            I => \N__50594\
        );

    \I__12096\ : LocalMux
    port map (
            O => \N__50666\,
            I => \N__50594\
        );

    \I__12095\ : Span4Mux_h
    port map (
            O => \N__50663\,
            I => \N__50594\
        );

    \I__12094\ : Span4Mux_v
    port map (
            O => \N__50660\,
            I => \N__50594\
        );

    \I__12093\ : Span4Mux_h
    port map (
            O => \N__50657\,
            I => \N__50589\
        );

    \I__12092\ : Span4Mux_h
    port map (
            O => \N__50652\,
            I => \N__50589\
        );

    \I__12091\ : InMux
    port map (
            O => \N__50651\,
            I => \N__50582\
        );

    \I__12090\ : InMux
    port map (
            O => \N__50650\,
            I => \N__50582\
        );

    \I__12089\ : InMux
    port map (
            O => \N__50649\,
            I => \N__50582\
        );

    \I__12088\ : InMux
    port map (
            O => \N__50648\,
            I => \N__50573\
        );

    \I__12087\ : InMux
    port map (
            O => \N__50647\,
            I => \N__50573\
        );

    \I__12086\ : InMux
    port map (
            O => \N__50646\,
            I => \N__50573\
        );

    \I__12085\ : InMux
    port map (
            O => \N__50645\,
            I => \N__50573\
        );

    \I__12084\ : LocalMux
    port map (
            O => \N__50642\,
            I => adc_state_0
        );

    \I__12083\ : LocalMux
    port map (
            O => \N__50639\,
            I => adc_state_0
        );

    \I__12082\ : Odrv4
    port map (
            O => \N__50636\,
            I => adc_state_0
        );

    \I__12081\ : LocalMux
    port map (
            O => \N__50619\,
            I => adc_state_0
        );

    \I__12080\ : Odrv4
    port map (
            O => \N__50614\,
            I => adc_state_0
        );

    \I__12079\ : Odrv4
    port map (
            O => \N__50611\,
            I => adc_state_0
        );

    \I__12078\ : Odrv12
    port map (
            O => \N__50606\,
            I => adc_state_0
        );

    \I__12077\ : Odrv12
    port map (
            O => \N__50603\,
            I => adc_state_0
        );

    \I__12076\ : Odrv4
    port map (
            O => \N__50594\,
            I => adc_state_0
        );

    \I__12075\ : Odrv4
    port map (
            O => \N__50589\,
            I => adc_state_0
        );

    \I__12074\ : LocalMux
    port map (
            O => \N__50582\,
            I => adc_state_0
        );

    \I__12073\ : LocalMux
    port map (
            O => \N__50573\,
            I => adc_state_0
        );

    \I__12072\ : CascadeMux
    port map (
            O => \N__50548\,
            I => \N__50544\
        );

    \I__12071\ : CascadeMux
    port map (
            O => \N__50547\,
            I => \N__50541\
        );

    \I__12070\ : InMux
    port map (
            O => \N__50544\,
            I => \N__50537\
        );

    \I__12069\ : InMux
    port map (
            O => \N__50541\,
            I => \N__50532\
        );

    \I__12068\ : InMux
    port map (
            O => \N__50540\,
            I => \N__50532\
        );

    \I__12067\ : LocalMux
    port map (
            O => \N__50537\,
            I => cmd_rdadctmp_12
        );

    \I__12066\ : LocalMux
    port map (
            O => \N__50532\,
            I => cmd_rdadctmp_12
        );

    \I__12065\ : InMux
    port map (
            O => \N__50527\,
            I => \N__50523\
        );

    \I__12064\ : InMux
    port map (
            O => \N__50526\,
            I => \N__50520\
        );

    \I__12063\ : LocalMux
    port map (
            O => \N__50523\,
            I => \N__50507\
        );

    \I__12062\ : LocalMux
    port map (
            O => \N__50520\,
            I => \N__50507\
        );

    \I__12061\ : InMux
    port map (
            O => \N__50519\,
            I => \N__50502\
        );

    \I__12060\ : InMux
    port map (
            O => \N__50518\,
            I => \N__50502\
        );

    \I__12059\ : InMux
    port map (
            O => \N__50517\,
            I => \N__50497\
        );

    \I__12058\ : InMux
    port map (
            O => \N__50516\,
            I => \N__50486\
        );

    \I__12057\ : InMux
    port map (
            O => \N__50515\,
            I => \N__50486\
        );

    \I__12056\ : InMux
    port map (
            O => \N__50514\,
            I => \N__50483\
        );

    \I__12055\ : InMux
    port map (
            O => \N__50513\,
            I => \N__50480\
        );

    \I__12054\ : InMux
    port map (
            O => \N__50512\,
            I => \N__50476\
        );

    \I__12053\ : Span4Mux_v
    port map (
            O => \N__50507\,
            I => \N__50471\
        );

    \I__12052\ : LocalMux
    port map (
            O => \N__50502\,
            I => \N__50471\
        );

    \I__12051\ : InMux
    port map (
            O => \N__50501\,
            I => \N__50466\
        );

    \I__12050\ : InMux
    port map (
            O => \N__50500\,
            I => \N__50463\
        );

    \I__12049\ : LocalMux
    port map (
            O => \N__50497\,
            I => \N__50460\
        );

    \I__12048\ : InMux
    port map (
            O => \N__50496\,
            I => \N__50448\
        );

    \I__12047\ : InMux
    port map (
            O => \N__50495\,
            I => \N__50448\
        );

    \I__12046\ : InMux
    port map (
            O => \N__50494\,
            I => \N__50443\
        );

    \I__12045\ : InMux
    port map (
            O => \N__50493\,
            I => \N__50443\
        );

    \I__12044\ : InMux
    port map (
            O => \N__50492\,
            I => \N__50438\
        );

    \I__12043\ : InMux
    port map (
            O => \N__50491\,
            I => \N__50438\
        );

    \I__12042\ : LocalMux
    port map (
            O => \N__50486\,
            I => \N__50431\
        );

    \I__12041\ : LocalMux
    port map (
            O => \N__50483\,
            I => \N__50431\
        );

    \I__12040\ : LocalMux
    port map (
            O => \N__50480\,
            I => \N__50431\
        );

    \I__12039\ : InMux
    port map (
            O => \N__50479\,
            I => \N__50428\
        );

    \I__12038\ : LocalMux
    port map (
            O => \N__50476\,
            I => \N__50425\
        );

    \I__12037\ : Span4Mux_h
    port map (
            O => \N__50471\,
            I => \N__50422\
        );

    \I__12036\ : CascadeMux
    port map (
            O => \N__50470\,
            I => \N__50419\
        );

    \I__12035\ : InMux
    port map (
            O => \N__50469\,
            I => \N__50412\
        );

    \I__12034\ : LocalMux
    port map (
            O => \N__50466\,
            I => \N__50409\
        );

    \I__12033\ : LocalMux
    port map (
            O => \N__50463\,
            I => \N__50406\
        );

    \I__12032\ : Span12Mux_v
    port map (
            O => \N__50460\,
            I => \N__50403\
        );

    \I__12031\ : InMux
    port map (
            O => \N__50459\,
            I => \N__50390\
        );

    \I__12030\ : InMux
    port map (
            O => \N__50458\,
            I => \N__50390\
        );

    \I__12029\ : InMux
    port map (
            O => \N__50457\,
            I => \N__50390\
        );

    \I__12028\ : InMux
    port map (
            O => \N__50456\,
            I => \N__50390\
        );

    \I__12027\ : InMux
    port map (
            O => \N__50455\,
            I => \N__50390\
        );

    \I__12026\ : InMux
    port map (
            O => \N__50454\,
            I => \N__50390\
        );

    \I__12025\ : InMux
    port map (
            O => \N__50453\,
            I => \N__50387\
        );

    \I__12024\ : LocalMux
    port map (
            O => \N__50448\,
            I => \N__50378\
        );

    \I__12023\ : LocalMux
    port map (
            O => \N__50443\,
            I => \N__50378\
        );

    \I__12022\ : LocalMux
    port map (
            O => \N__50438\,
            I => \N__50378\
        );

    \I__12021\ : Span4Mux_v
    port map (
            O => \N__50431\,
            I => \N__50378\
        );

    \I__12020\ : LocalMux
    port map (
            O => \N__50428\,
            I => \N__50373\
        );

    \I__12019\ : Span4Mux_v
    port map (
            O => \N__50425\,
            I => \N__50373\
        );

    \I__12018\ : Span4Mux_h
    port map (
            O => \N__50422\,
            I => \N__50370\
        );

    \I__12017\ : InMux
    port map (
            O => \N__50419\,
            I => \N__50367\
        );

    \I__12016\ : InMux
    port map (
            O => \N__50418\,
            I => \N__50358\
        );

    \I__12015\ : InMux
    port map (
            O => \N__50417\,
            I => \N__50358\
        );

    \I__12014\ : InMux
    port map (
            O => \N__50416\,
            I => \N__50358\
        );

    \I__12013\ : InMux
    port map (
            O => \N__50415\,
            I => \N__50358\
        );

    \I__12012\ : LocalMux
    port map (
            O => \N__50412\,
            I => \N__50353\
        );

    \I__12011\ : Span4Mux_v
    port map (
            O => \N__50409\,
            I => \N__50353\
        );

    \I__12010\ : Span4Mux_h
    port map (
            O => \N__50406\,
            I => \N__50350\
        );

    \I__12009\ : Span12Mux_h
    port map (
            O => \N__50403\,
            I => \N__50347\
        );

    \I__12008\ : LocalMux
    port map (
            O => \N__50390\,
            I => \N__50336\
        );

    \I__12007\ : LocalMux
    port map (
            O => \N__50387\,
            I => \N__50336\
        );

    \I__12006\ : Span4Mux_v
    port map (
            O => \N__50378\,
            I => \N__50336\
        );

    \I__12005\ : Span4Mux_v
    port map (
            O => \N__50373\,
            I => \N__50336\
        );

    \I__12004\ : Span4Mux_v
    port map (
            O => \N__50370\,
            I => \N__50336\
        );

    \I__12003\ : LocalMux
    port map (
            O => \N__50367\,
            I => n12542
        );

    \I__12002\ : LocalMux
    port map (
            O => \N__50358\,
            I => n12542
        );

    \I__12001\ : Odrv4
    port map (
            O => \N__50353\,
            I => n12542
        );

    \I__12000\ : Odrv4
    port map (
            O => \N__50350\,
            I => n12542
        );

    \I__11999\ : Odrv12
    port map (
            O => \N__50347\,
            I => n12542
        );

    \I__11998\ : Odrv4
    port map (
            O => \N__50336\,
            I => n12542
        );

    \I__11997\ : CascadeMux
    port map (
            O => \N__50323\,
            I => \N__50319\
        );

    \I__11996\ : CascadeMux
    port map (
            O => \N__50322\,
            I => \N__50316\
        );

    \I__11995\ : InMux
    port map (
            O => \N__50319\,
            I => \N__50312\
        );

    \I__11994\ : InMux
    port map (
            O => \N__50316\,
            I => \N__50309\
        );

    \I__11993\ : InMux
    port map (
            O => \N__50315\,
            I => \N__50306\
        );

    \I__11992\ : LocalMux
    port map (
            O => \N__50312\,
            I => cmd_rdadctmp_13
        );

    \I__11991\ : LocalMux
    port map (
            O => \N__50309\,
            I => cmd_rdadctmp_13
        );

    \I__11990\ : LocalMux
    port map (
            O => \N__50306\,
            I => cmd_rdadctmp_13
        );

    \I__11989\ : InMux
    port map (
            O => \N__50299\,
            I => \N__50296\
        );

    \I__11988\ : LocalMux
    port map (
            O => \N__50296\,
            I => \N__50293\
        );

    \I__11987\ : Span4Mux_h
    port map (
            O => \N__50293\,
            I => \N__50289\
        );

    \I__11986\ : InMux
    port map (
            O => \N__50292\,
            I => \N__50286\
        );

    \I__11985\ : Span4Mux_h
    port map (
            O => \N__50289\,
            I => \N__50282\
        );

    \I__11984\ : LocalMux
    port map (
            O => \N__50286\,
            I => \N__50279\
        );

    \I__11983\ : InMux
    port map (
            O => \N__50285\,
            I => \N__50276\
        );

    \I__11982\ : Span4Mux_v
    port map (
            O => \N__50282\,
            I => \N__50273\
        );

    \I__11981\ : Odrv12
    port map (
            O => \N__50279\,
            I => buf_control_0
        );

    \I__11980\ : LocalMux
    port map (
            O => \N__50276\,
            I => buf_control_0
        );

    \I__11979\ : Odrv4
    port map (
            O => \N__50273\,
            I => buf_control_0
        );

    \I__11978\ : InMux
    port map (
            O => \N__50266\,
            I => \N__50263\
        );

    \I__11977\ : LocalMux
    port map (
            O => \N__50263\,
            I => \N__50260\
        );

    \I__11976\ : Sp12to4
    port map (
            O => \N__50260\,
            I => \N__50257\
        );

    \I__11975\ : Span12Mux_v
    port map (
            O => \N__50257\,
            I => \N__50252\
        );

    \I__11974\ : InMux
    port map (
            O => \N__50256\,
            I => \N__50249\
        );

    \I__11973\ : InMux
    port map (
            O => \N__50255\,
            I => \N__50246\
        );

    \I__11972\ : Odrv12
    port map (
            O => \N__50252\,
            I => wdtick_flag
        );

    \I__11971\ : LocalMux
    port map (
            O => \N__50249\,
            I => wdtick_flag
        );

    \I__11970\ : LocalMux
    port map (
            O => \N__50246\,
            I => wdtick_flag
        );

    \I__11969\ : IoInMux
    port map (
            O => \N__50239\,
            I => \N__50236\
        );

    \I__11968\ : LocalMux
    port map (
            O => \N__50236\,
            I => \N__50233\
        );

    \I__11967\ : Span4Mux_s1_v
    port map (
            O => \N__50233\,
            I => \N__50230\
        );

    \I__11966\ : Span4Mux_v
    port map (
            O => \N__50230\,
            I => \N__50227\
        );

    \I__11965\ : Span4Mux_v
    port map (
            O => \N__50227\,
            I => \N__50224\
        );

    \I__11964\ : Odrv4
    port map (
            O => \N__50224\,
            I => \CONT_SD\
        );

    \I__11963\ : InMux
    port map (
            O => \N__50221\,
            I => \N__50217\
        );

    \I__11962\ : InMux
    port map (
            O => \N__50220\,
            I => \N__50214\
        );

    \I__11961\ : LocalMux
    port map (
            O => \N__50217\,
            I => \N__50211\
        );

    \I__11960\ : LocalMux
    port map (
            O => \N__50214\,
            I => \N__50206\
        );

    \I__11959\ : Span4Mux_v
    port map (
            O => \N__50211\,
            I => \N__50206\
        );

    \I__11958\ : Span4Mux_h
    port map (
            O => \N__50206\,
            I => \N__50202\
        );

    \I__11957\ : InMux
    port map (
            O => \N__50205\,
            I => \N__50199\
        );

    \I__11956\ : Odrv4
    port map (
            O => \N__50202\,
            I => \comm_spi.n22647\
        );

    \I__11955\ : LocalMux
    port map (
            O => \N__50199\,
            I => \comm_spi.n22647\
        );

    \I__11954\ : InMux
    port map (
            O => \N__50194\,
            I => \N__50191\
        );

    \I__11953\ : LocalMux
    port map (
            O => \N__50191\,
            I => \N__50187\
        );

    \I__11952\ : CascadeMux
    port map (
            O => \N__50190\,
            I => \N__50184\
        );

    \I__11951\ : Span4Mux_v
    port map (
            O => \N__50187\,
            I => \N__50178\
        );

    \I__11950\ : InMux
    port map (
            O => \N__50184\,
            I => \N__50175\
        );

    \I__11949\ : InMux
    port map (
            O => \N__50183\,
            I => \N__50172\
        );

    \I__11948\ : InMux
    port map (
            O => \N__50182\,
            I => \N__50169\
        );

    \I__11947\ : InMux
    port map (
            O => \N__50181\,
            I => \N__50166\
        );

    \I__11946\ : Span4Mux_v
    port map (
            O => \N__50178\,
            I => \N__50163\
        );

    \I__11945\ : LocalMux
    port map (
            O => \N__50175\,
            I => \N__50158\
        );

    \I__11944\ : LocalMux
    port map (
            O => \N__50172\,
            I => \N__50158\
        );

    \I__11943\ : LocalMux
    port map (
            O => \N__50169\,
            I => \N__50155\
        );

    \I__11942\ : LocalMux
    port map (
            O => \N__50166\,
            I => \N__50148\
        );

    \I__11941\ : Span4Mux_h
    port map (
            O => \N__50163\,
            I => \N__50148\
        );

    \I__11940\ : Span4Mux_v
    port map (
            O => \N__50158\,
            I => \N__50148\
        );

    \I__11939\ : Span4Mux_h
    port map (
            O => \N__50155\,
            I => \N__50145\
        );

    \I__11938\ : Span4Mux_h
    port map (
            O => \N__50148\,
            I => \N__50142\
        );

    \I__11937\ : Odrv4
    port map (
            O => \N__50145\,
            I => comm_buf_1_5
        );

    \I__11936\ : Odrv4
    port map (
            O => \N__50142\,
            I => comm_buf_1_5
        );

    \I__11935\ : CascadeMux
    port map (
            O => \N__50137\,
            I => \N__50133\
        );

    \I__11934\ : InMux
    port map (
            O => \N__50136\,
            I => \N__50129\
        );

    \I__11933\ : InMux
    port map (
            O => \N__50133\,
            I => \N__50126\
        );

    \I__11932\ : InMux
    port map (
            O => \N__50132\,
            I => \N__50123\
        );

    \I__11931\ : LocalMux
    port map (
            O => \N__50129\,
            I => \N__50120\
        );

    \I__11930\ : LocalMux
    port map (
            O => \N__50126\,
            I => \N__50115\
        );

    \I__11929\ : LocalMux
    port map (
            O => \N__50123\,
            I => \N__50115\
        );

    \I__11928\ : Span4Mux_v
    port map (
            O => \N__50120\,
            I => \N__50110\
        );

    \I__11927\ : Span4Mux_h
    port map (
            O => \N__50115\,
            I => \N__50110\
        );

    \I__11926\ : Span4Mux_h
    port map (
            O => \N__50110\,
            I => \N__50107\
        );

    \I__11925\ : Span4Mux_h
    port map (
            O => \N__50107\,
            I => \N__50104\
        );

    \I__11924\ : Odrv4
    port map (
            O => \N__50104\,
            I => n14_adj_1557
        );

    \I__11923\ : InMux
    port map (
            O => \N__50101\,
            I => \N__50089\
        );

    \I__11922\ : InMux
    port map (
            O => \N__50100\,
            I => \N__50089\
        );

    \I__11921\ : InMux
    port map (
            O => \N__50099\,
            I => \N__50082\
        );

    \I__11920\ : InMux
    port map (
            O => \N__50098\,
            I => \N__50082\
        );

    \I__11919\ : InMux
    port map (
            O => \N__50097\,
            I => \N__50079\
        );

    \I__11918\ : InMux
    port map (
            O => \N__50096\,
            I => \N__50070\
        );

    \I__11917\ : InMux
    port map (
            O => \N__50095\,
            I => \N__50070\
        );

    \I__11916\ : CascadeMux
    port map (
            O => \N__50094\,
            I => \N__50064\
        );

    \I__11915\ : LocalMux
    port map (
            O => \N__50089\,
            I => \N__50061\
        );

    \I__11914\ : InMux
    port map (
            O => \N__50088\,
            I => \N__50058\
        );

    \I__11913\ : InMux
    port map (
            O => \N__50087\,
            I => \N__50055\
        );

    \I__11912\ : LocalMux
    port map (
            O => \N__50082\,
            I => \N__50050\
        );

    \I__11911\ : LocalMux
    port map (
            O => \N__50079\,
            I => \N__50050\
        );

    \I__11910\ : InMux
    port map (
            O => \N__50078\,
            I => \N__50047\
        );

    \I__11909\ : InMux
    port map (
            O => \N__50077\,
            I => \N__50040\
        );

    \I__11908\ : InMux
    port map (
            O => \N__50076\,
            I => \N__50040\
        );

    \I__11907\ : InMux
    port map (
            O => \N__50075\,
            I => \N__50040\
        );

    \I__11906\ : LocalMux
    port map (
            O => \N__50070\,
            I => \N__50037\
        );

    \I__11905\ : InMux
    port map (
            O => \N__50069\,
            I => \N__50030\
        );

    \I__11904\ : InMux
    port map (
            O => \N__50068\,
            I => \N__50030\
        );

    \I__11903\ : InMux
    port map (
            O => \N__50067\,
            I => \N__50030\
        );

    \I__11902\ : InMux
    port map (
            O => \N__50064\,
            I => \N__50027\
        );

    \I__11901\ : Span4Mux_v
    port map (
            O => \N__50061\,
            I => \N__50016\
        );

    \I__11900\ : LocalMux
    port map (
            O => \N__50058\,
            I => \N__50016\
        );

    \I__11899\ : LocalMux
    port map (
            O => \N__50055\,
            I => \N__50016\
        );

    \I__11898\ : Span4Mux_h
    port map (
            O => \N__50050\,
            I => \N__50016\
        );

    \I__11897\ : LocalMux
    port map (
            O => \N__50047\,
            I => \N__50016\
        );

    \I__11896\ : LocalMux
    port map (
            O => \N__50040\,
            I => \N__50011\
        );

    \I__11895\ : Span4Mux_v
    port map (
            O => \N__50037\,
            I => \N__50011\
        );

    \I__11894\ : LocalMux
    port map (
            O => \N__50030\,
            I => \N__50003\
        );

    \I__11893\ : LocalMux
    port map (
            O => \N__50027\,
            I => \N__49999\
        );

    \I__11892\ : Span4Mux_v
    port map (
            O => \N__50016\,
            I => \N__49994\
        );

    \I__11891\ : Span4Mux_h
    port map (
            O => \N__50011\,
            I => \N__49994\
        );

    \I__11890\ : InMux
    port map (
            O => \N__50010\,
            I => \N__49989\
        );

    \I__11889\ : InMux
    port map (
            O => \N__50009\,
            I => \N__49989\
        );

    \I__11888\ : InMux
    port map (
            O => \N__50008\,
            I => \N__49986\
        );

    \I__11887\ : InMux
    port map (
            O => \N__50007\,
            I => \N__49981\
        );

    \I__11886\ : InMux
    port map (
            O => \N__50006\,
            I => \N__49981\
        );

    \I__11885\ : Span12Mux_v
    port map (
            O => \N__50003\,
            I => \N__49978\
        );

    \I__11884\ : InMux
    port map (
            O => \N__50002\,
            I => \N__49975\
        );

    \I__11883\ : Span4Mux_h
    port map (
            O => \N__49999\,
            I => \N__49968\
        );

    \I__11882\ : Span4Mux_h
    port map (
            O => \N__49994\,
            I => \N__49968\
        );

    \I__11881\ : LocalMux
    port map (
            O => \N__49989\,
            I => \N__49968\
        );

    \I__11880\ : LocalMux
    port map (
            O => \N__49986\,
            I => comm_index_2
        );

    \I__11879\ : LocalMux
    port map (
            O => \N__49981\,
            I => comm_index_2
        );

    \I__11878\ : Odrv12
    port map (
            O => \N__49978\,
            I => comm_index_2
        );

    \I__11877\ : LocalMux
    port map (
            O => \N__49975\,
            I => comm_index_2
        );

    \I__11876\ : Odrv4
    port map (
            O => \N__49968\,
            I => comm_index_2
        );

    \I__11875\ : CascadeMux
    port map (
            O => \N__49957\,
            I => \N__49954\
        );

    \I__11874\ : InMux
    port map (
            O => \N__49954\,
            I => \N__49951\
        );

    \I__11873\ : LocalMux
    port map (
            O => \N__49951\,
            I => \N__49948\
        );

    \I__11872\ : Span4Mux_h
    port map (
            O => \N__49948\,
            I => \N__49944\
        );

    \I__11871\ : InMux
    port map (
            O => \N__49947\,
            I => \N__49941\
        );

    \I__11870\ : Span4Mux_h
    port map (
            O => \N__49944\,
            I => \N__49936\
        );

    \I__11869\ : LocalMux
    port map (
            O => \N__49941\,
            I => \N__49933\
        );

    \I__11868\ : InMux
    port map (
            O => \N__49940\,
            I => \N__49930\
        );

    \I__11867\ : InMux
    port map (
            O => \N__49939\,
            I => \N__49927\
        );

    \I__11866\ : Odrv4
    port map (
            O => \N__49936\,
            I => n18824
        );

    \I__11865\ : Odrv12
    port map (
            O => \N__49933\,
            I => n18824
        );

    \I__11864\ : LocalMux
    port map (
            O => \N__49930\,
            I => n18824
        );

    \I__11863\ : LocalMux
    port map (
            O => \N__49927\,
            I => n18824
        );

    \I__11862\ : CascadeMux
    port map (
            O => \N__49918\,
            I => \n20563_cascade_\
        );

    \I__11861\ : InMux
    port map (
            O => \N__49915\,
            I => \N__49911\
        );

    \I__11860\ : InMux
    port map (
            O => \N__49914\,
            I => \N__49905\
        );

    \I__11859\ : LocalMux
    port map (
            O => \N__49911\,
            I => \N__49902\
        );

    \I__11858\ : InMux
    port map (
            O => \N__49910\,
            I => \N__49897\
        );

    \I__11857\ : InMux
    port map (
            O => \N__49909\,
            I => \N__49897\
        );

    \I__11856\ : InMux
    port map (
            O => \N__49908\,
            I => \N__49894\
        );

    \I__11855\ : LocalMux
    port map (
            O => \N__49905\,
            I => \N__49891\
        );

    \I__11854\ : Span4Mux_h
    port map (
            O => \N__49902\,
            I => \N__49888\
        );

    \I__11853\ : LocalMux
    port map (
            O => \N__49897\,
            I => \N__49883\
        );

    \I__11852\ : LocalMux
    port map (
            O => \N__49894\,
            I => \N__49883\
        );

    \I__11851\ : Span4Mux_h
    port map (
            O => \N__49891\,
            I => \N__49876\
        );

    \I__11850\ : Span4Mux_h
    port map (
            O => \N__49888\,
            I => \N__49876\
        );

    \I__11849\ : Span4Mux_v
    port map (
            O => \N__49883\,
            I => \N__49876\
        );

    \I__11848\ : Odrv4
    port map (
            O => \N__49876\,
            I => n20627
        );

    \I__11847\ : CascadeMux
    port map (
            O => \N__49873\,
            I => \n12_adj_1539_cascade_\
        );

    \I__11846\ : InMux
    port map (
            O => \N__49870\,
            I => \N__49864\
        );

    \I__11845\ : InMux
    port map (
            O => \N__49869\,
            I => \N__49864\
        );

    \I__11844\ : LocalMux
    port map (
            O => \N__49864\,
            I => \N__49861\
        );

    \I__11843\ : Span4Mux_h
    port map (
            O => \N__49861\,
            I => \N__49855\
        );

    \I__11842\ : InMux
    port map (
            O => \N__49860\,
            I => \N__49850\
        );

    \I__11841\ : InMux
    port map (
            O => \N__49859\,
            I => \N__49850\
        );

    \I__11840\ : InMux
    port map (
            O => \N__49858\,
            I => \N__49847\
        );

    \I__11839\ : Span4Mux_h
    port map (
            O => \N__49855\,
            I => \N__49839\
        );

    \I__11838\ : LocalMux
    port map (
            O => \N__49850\,
            I => \N__49839\
        );

    \I__11837\ : LocalMux
    port map (
            O => \N__49847\,
            I => \N__49839\
        );

    \I__11836\ : InMux
    port map (
            O => \N__49846\,
            I => \N__49836\
        );

    \I__11835\ : Span4Mux_v
    port map (
            O => \N__49839\,
            I => \N__49831\
        );

    \I__11834\ : LocalMux
    port map (
            O => \N__49836\,
            I => \N__49831\
        );

    \I__11833\ : Span4Mux_h
    port map (
            O => \N__49831\,
            I => \N__49828\
        );

    \I__11832\ : Odrv4
    port map (
            O => \N__49828\,
            I => n20556
        );

    \I__11831\ : CEMux
    port map (
            O => \N__49825\,
            I => \N__49822\
        );

    \I__11830\ : LocalMux
    port map (
            O => \N__49822\,
            I => \N__49818\
        );

    \I__11829\ : InMux
    port map (
            O => \N__49821\,
            I => \N__49815\
        );

    \I__11828\ : Span4Mux_v
    port map (
            O => \N__49818\,
            I => \N__49812\
        );

    \I__11827\ : LocalMux
    port map (
            O => \N__49815\,
            I => \N__49809\
        );

    \I__11826\ : Span4Mux_h
    port map (
            O => \N__49812\,
            I => \N__49804\
        );

    \I__11825\ : Span4Mux_h
    port map (
            O => \N__49809\,
            I => \N__49804\
        );

    \I__11824\ : Odrv4
    port map (
            O => \N__49804\,
            I => n12164
        );

    \I__11823\ : InMux
    port map (
            O => \N__49801\,
            I => \N__49792\
        );

    \I__11822\ : InMux
    port map (
            O => \N__49800\,
            I => \N__49783\
        );

    \I__11821\ : InMux
    port map (
            O => \N__49799\,
            I => \N__49783\
        );

    \I__11820\ : InMux
    port map (
            O => \N__49798\,
            I => \N__49783\
        );

    \I__11819\ : CascadeMux
    port map (
            O => \N__49797\,
            I => \N__49778\
        );

    \I__11818\ : CascadeMux
    port map (
            O => \N__49796\,
            I => \N__49775\
        );

    \I__11817\ : CascadeMux
    port map (
            O => \N__49795\,
            I => \N__49771\
        );

    \I__11816\ : LocalMux
    port map (
            O => \N__49792\,
            I => \N__49764\
        );

    \I__11815\ : InMux
    port map (
            O => \N__49791\,
            I => \N__49759\
        );

    \I__11814\ : InMux
    port map (
            O => \N__49790\,
            I => \N__49759\
        );

    \I__11813\ : LocalMux
    port map (
            O => \N__49783\,
            I => \N__49756\
        );

    \I__11812\ : CascadeMux
    port map (
            O => \N__49782\,
            I => \N__49752\
        );

    \I__11811\ : InMux
    port map (
            O => \N__49781\,
            I => \N__49747\
        );

    \I__11810\ : InMux
    port map (
            O => \N__49778\,
            I => \N__49744\
        );

    \I__11809\ : InMux
    port map (
            O => \N__49775\,
            I => \N__49735\
        );

    \I__11808\ : InMux
    port map (
            O => \N__49774\,
            I => \N__49735\
        );

    \I__11807\ : InMux
    port map (
            O => \N__49771\,
            I => \N__49735\
        );

    \I__11806\ : InMux
    port map (
            O => \N__49770\,
            I => \N__49735\
        );

    \I__11805\ : InMux
    port map (
            O => \N__49769\,
            I => \N__49730\
        );

    \I__11804\ : InMux
    port map (
            O => \N__49768\,
            I => \N__49730\
        );

    \I__11803\ : InMux
    port map (
            O => \N__49767\,
            I => \N__49727\
        );

    \I__11802\ : Span4Mux_v
    port map (
            O => \N__49764\,
            I => \N__49722\
        );

    \I__11801\ : LocalMux
    port map (
            O => \N__49759\,
            I => \N__49722\
        );

    \I__11800\ : Span4Mux_v
    port map (
            O => \N__49756\,
            I => \N__49719\
        );

    \I__11799\ : InMux
    port map (
            O => \N__49755\,
            I => \N__49712\
        );

    \I__11798\ : InMux
    port map (
            O => \N__49752\,
            I => \N__49712\
        );

    \I__11797\ : InMux
    port map (
            O => \N__49751\,
            I => \N__49712\
        );

    \I__11796\ : InMux
    port map (
            O => \N__49750\,
            I => \N__49709\
        );

    \I__11795\ : LocalMux
    port map (
            O => \N__49747\,
            I => \N__49700\
        );

    \I__11794\ : LocalMux
    port map (
            O => \N__49744\,
            I => \N__49700\
        );

    \I__11793\ : LocalMux
    port map (
            O => \N__49735\,
            I => \N__49700\
        );

    \I__11792\ : LocalMux
    port map (
            O => \N__49730\,
            I => \N__49700\
        );

    \I__11791\ : LocalMux
    port map (
            O => \N__49727\,
            I => \N__49696\
        );

    \I__11790\ : Span4Mux_v
    port map (
            O => \N__49722\,
            I => \N__49693\
        );

    \I__11789\ : Span4Mux_h
    port map (
            O => \N__49719\,
            I => \N__49690\
        );

    \I__11788\ : LocalMux
    port map (
            O => \N__49712\,
            I => \N__49683\
        );

    \I__11787\ : LocalMux
    port map (
            O => \N__49709\,
            I => \N__49683\
        );

    \I__11786\ : Span4Mux_v
    port map (
            O => \N__49700\,
            I => \N__49683\
        );

    \I__11785\ : InMux
    port map (
            O => \N__49699\,
            I => \N__49680\
        );

    \I__11784\ : Sp12to4
    port map (
            O => \N__49696\,
            I => \N__49677\
        );

    \I__11783\ : Sp12to4
    port map (
            O => \N__49693\,
            I => \N__49674\
        );

    \I__11782\ : Span4Mux_h
    port map (
            O => \N__49690\,
            I => \N__49671\
        );

    \I__11781\ : Sp12to4
    port map (
            O => \N__49683\,
            I => \N__49666\
        );

    \I__11780\ : LocalMux
    port map (
            O => \N__49680\,
            I => \N__49666\
        );

    \I__11779\ : Span12Mux_v
    port map (
            O => \N__49677\,
            I => \N__49661\
        );

    \I__11778\ : Span12Mux_s10_h
    port map (
            O => \N__49674\,
            I => \N__49661\
        );

    \I__11777\ : Sp12to4
    port map (
            O => \N__49671\,
            I => \N__49656\
        );

    \I__11776\ : Span12Mux_h
    port map (
            O => \N__49666\,
            I => \N__49656\
        );

    \I__11775\ : Span12Mux_v
    port map (
            O => \N__49661\,
            I => \N__49653\
        );

    \I__11774\ : Span12Mux_v
    port map (
            O => \N__49656\,
            I => \N__49650\
        );

    \I__11773\ : Odrv12
    port map (
            O => \N__49653\,
            I => \ICE_SPI_CE0\
        );

    \I__11772\ : Odrv12
    port map (
            O => \N__49650\,
            I => \ICE_SPI_CE0\
        );

    \I__11771\ : InMux
    port map (
            O => \N__49645\,
            I => \N__49642\
        );

    \I__11770\ : LocalMux
    port map (
            O => \N__49642\,
            I => \N__49636\
        );

    \I__11769\ : InMux
    port map (
            O => \N__49641\,
            I => \N__49629\
        );

    \I__11768\ : InMux
    port map (
            O => \N__49640\,
            I => \N__49619\
        );

    \I__11767\ : InMux
    port map (
            O => \N__49639\,
            I => \N__49619\
        );

    \I__11766\ : Span4Mux_v
    port map (
            O => \N__49636\,
            I => \N__49616\
        );

    \I__11765\ : InMux
    port map (
            O => \N__49635\,
            I => \N__49613\
        );

    \I__11764\ : InMux
    port map (
            O => \N__49634\,
            I => \N__49610\
        );

    \I__11763\ : InMux
    port map (
            O => \N__49633\,
            I => \N__49605\
        );

    \I__11762\ : InMux
    port map (
            O => \N__49632\,
            I => \N__49605\
        );

    \I__11761\ : LocalMux
    port map (
            O => \N__49629\,
            I => \N__49602\
        );

    \I__11760\ : InMux
    port map (
            O => \N__49628\,
            I => \N__49593\
        );

    \I__11759\ : InMux
    port map (
            O => \N__49627\,
            I => \N__49593\
        );

    \I__11758\ : InMux
    port map (
            O => \N__49626\,
            I => \N__49593\
        );

    \I__11757\ : InMux
    port map (
            O => \N__49625\,
            I => \N__49593\
        );

    \I__11756\ : InMux
    port map (
            O => \N__49624\,
            I => \N__49590\
        );

    \I__11755\ : LocalMux
    port map (
            O => \N__49619\,
            I => comm_data_vld
        );

    \I__11754\ : Odrv4
    port map (
            O => \N__49616\,
            I => comm_data_vld
        );

    \I__11753\ : LocalMux
    port map (
            O => \N__49613\,
            I => comm_data_vld
        );

    \I__11752\ : LocalMux
    port map (
            O => \N__49610\,
            I => comm_data_vld
        );

    \I__11751\ : LocalMux
    port map (
            O => \N__49605\,
            I => comm_data_vld
        );

    \I__11750\ : Odrv4
    port map (
            O => \N__49602\,
            I => comm_data_vld
        );

    \I__11749\ : LocalMux
    port map (
            O => \N__49593\,
            I => comm_data_vld
        );

    \I__11748\ : LocalMux
    port map (
            O => \N__49590\,
            I => comm_data_vld
        );

    \I__11747\ : InMux
    port map (
            O => \N__49573\,
            I => \N__49570\
        );

    \I__11746\ : LocalMux
    port map (
            O => \N__49570\,
            I => \N__49567\
        );

    \I__11745\ : Span4Mux_h
    port map (
            O => \N__49567\,
            I => \N__49564\
        );

    \I__11744\ : Span4Mux_v
    port map (
            O => \N__49564\,
            I => \N__49561\
        );

    \I__11743\ : Odrv4
    port map (
            O => \N__49561\,
            I => n23_adj_1574
        );

    \I__11742\ : CascadeMux
    port map (
            O => \N__49558\,
            I => \n21_adj_1573_cascade_\
        );

    \I__11741\ : CEMux
    port map (
            O => \N__49555\,
            I => \N__49552\
        );

    \I__11740\ : LocalMux
    port map (
            O => \N__49552\,
            I => \N__49549\
        );

    \I__11739\ : Span4Mux_h
    port map (
            O => \N__49549\,
            I => \N__49546\
        );

    \I__11738\ : Odrv4
    port map (
            O => \N__49546\,
            I => n18
        );

    \I__11737\ : CascadeMux
    port map (
            O => \N__49543\,
            I => \N__49540\
        );

    \I__11736\ : InMux
    port map (
            O => \N__49540\,
            I => \N__49526\
        );

    \I__11735\ : InMux
    port map (
            O => \N__49539\,
            I => \N__49515\
        );

    \I__11734\ : InMux
    port map (
            O => \N__49538\,
            I => \N__49515\
        );

    \I__11733\ : InMux
    port map (
            O => \N__49537\,
            I => \N__49506\
        );

    \I__11732\ : InMux
    port map (
            O => \N__49536\,
            I => \N__49506\
        );

    \I__11731\ : InMux
    port map (
            O => \N__49535\,
            I => \N__49506\
        );

    \I__11730\ : InMux
    port map (
            O => \N__49534\,
            I => \N__49503\
        );

    \I__11729\ : InMux
    port map (
            O => \N__49533\,
            I => \N__49500\
        );

    \I__11728\ : InMux
    port map (
            O => \N__49532\,
            I => \N__49493\
        );

    \I__11727\ : InMux
    port map (
            O => \N__49531\,
            I => \N__49493\
        );

    \I__11726\ : InMux
    port map (
            O => \N__49530\,
            I => \N__49493\
        );

    \I__11725\ : InMux
    port map (
            O => \N__49529\,
            I => \N__49489\
        );

    \I__11724\ : LocalMux
    port map (
            O => \N__49526\,
            I => \N__49486\
        );

    \I__11723\ : InMux
    port map (
            O => \N__49525\,
            I => \N__49481\
        );

    \I__11722\ : InMux
    port map (
            O => \N__49524\,
            I => \N__49481\
        );

    \I__11721\ : InMux
    port map (
            O => \N__49523\,
            I => \N__49476\
        );

    \I__11720\ : InMux
    port map (
            O => \N__49522\,
            I => \N__49476\
        );

    \I__11719\ : InMux
    port map (
            O => \N__49521\,
            I => \N__49471\
        );

    \I__11718\ : InMux
    port map (
            O => \N__49520\,
            I => \N__49471\
        );

    \I__11717\ : LocalMux
    port map (
            O => \N__49515\,
            I => \N__49468\
        );

    \I__11716\ : CascadeMux
    port map (
            O => \N__49514\,
            I => \N__49464\
        );

    \I__11715\ : CascadeMux
    port map (
            O => \N__49513\,
            I => \N__49459\
        );

    \I__11714\ : LocalMux
    port map (
            O => \N__49506\,
            I => \N__49456\
        );

    \I__11713\ : LocalMux
    port map (
            O => \N__49503\,
            I => \N__49451\
        );

    \I__11712\ : LocalMux
    port map (
            O => \N__49500\,
            I => \N__49451\
        );

    \I__11711\ : LocalMux
    port map (
            O => \N__49493\,
            I => \N__49448\
        );

    \I__11710\ : InMux
    port map (
            O => \N__49492\,
            I => \N__49445\
        );

    \I__11709\ : LocalMux
    port map (
            O => \N__49489\,
            I => \N__49442\
        );

    \I__11708\ : Span4Mux_v
    port map (
            O => \N__49486\,
            I => \N__49435\
        );

    \I__11707\ : LocalMux
    port map (
            O => \N__49481\,
            I => \N__49435\
        );

    \I__11706\ : LocalMux
    port map (
            O => \N__49476\,
            I => \N__49435\
        );

    \I__11705\ : LocalMux
    port map (
            O => \N__49471\,
            I => \N__49430\
        );

    \I__11704\ : Span4Mux_h
    port map (
            O => \N__49468\,
            I => \N__49430\
        );

    \I__11703\ : InMux
    port map (
            O => \N__49467\,
            I => \N__49426\
        );

    \I__11702\ : InMux
    port map (
            O => \N__49464\,
            I => \N__49423\
        );

    \I__11701\ : InMux
    port map (
            O => \N__49463\,
            I => \N__49420\
        );

    \I__11700\ : InMux
    port map (
            O => \N__49462\,
            I => \N__49417\
        );

    \I__11699\ : InMux
    port map (
            O => \N__49459\,
            I => \N__49414\
        );

    \I__11698\ : Span4Mux_v
    port map (
            O => \N__49456\,
            I => \N__49407\
        );

    \I__11697\ : Span4Mux_v
    port map (
            O => \N__49451\,
            I => \N__49407\
        );

    \I__11696\ : Span4Mux_v
    port map (
            O => \N__49448\,
            I => \N__49407\
        );

    \I__11695\ : LocalMux
    port map (
            O => \N__49445\,
            I => \N__49404\
        );

    \I__11694\ : Span4Mux_v
    port map (
            O => \N__49442\,
            I => \N__49397\
        );

    \I__11693\ : Span4Mux_v
    port map (
            O => \N__49435\,
            I => \N__49397\
        );

    \I__11692\ : Span4Mux_h
    port map (
            O => \N__49430\,
            I => \N__49397\
        );

    \I__11691\ : CascadeMux
    port map (
            O => \N__49429\,
            I => \N__49392\
        );

    \I__11690\ : LocalMux
    port map (
            O => \N__49426\,
            I => \N__49387\
        );

    \I__11689\ : LocalMux
    port map (
            O => \N__49423\,
            I => \N__49387\
        );

    \I__11688\ : LocalMux
    port map (
            O => \N__49420\,
            I => \N__49384\
        );

    \I__11687\ : LocalMux
    port map (
            O => \N__49417\,
            I => \N__49375\
        );

    \I__11686\ : LocalMux
    port map (
            O => \N__49414\,
            I => \N__49375\
        );

    \I__11685\ : Span4Mux_h
    port map (
            O => \N__49407\,
            I => \N__49375\
        );

    \I__11684\ : Span4Mux_v
    port map (
            O => \N__49404\,
            I => \N__49375\
        );

    \I__11683\ : Span4Mux_h
    port map (
            O => \N__49397\,
            I => \N__49372\
        );

    \I__11682\ : InMux
    port map (
            O => \N__49396\,
            I => \N__49367\
        );

    \I__11681\ : InMux
    port map (
            O => \N__49395\,
            I => \N__49367\
        );

    \I__11680\ : InMux
    port map (
            O => \N__49392\,
            I => \N__49364\
        );

    \I__11679\ : Span4Mux_h
    port map (
            O => \N__49387\,
            I => \N__49361\
        );

    \I__11678\ : Odrv4
    port map (
            O => \N__49384\,
            I => comm_index_1
        );

    \I__11677\ : Odrv4
    port map (
            O => \N__49375\,
            I => comm_index_1
        );

    \I__11676\ : Odrv4
    port map (
            O => \N__49372\,
            I => comm_index_1
        );

    \I__11675\ : LocalMux
    port map (
            O => \N__49367\,
            I => comm_index_1
        );

    \I__11674\ : LocalMux
    port map (
            O => \N__49364\,
            I => comm_index_1
        );

    \I__11673\ : Odrv4
    port map (
            O => \N__49361\,
            I => comm_index_1
        );

    \I__11672\ : CascadeMux
    port map (
            O => \N__49348\,
            I => \N__49345\
        );

    \I__11671\ : InMux
    port map (
            O => \N__49345\,
            I => \N__49341\
        );

    \I__11670\ : InMux
    port map (
            O => \N__49344\,
            I => \N__49338\
        );

    \I__11669\ : LocalMux
    port map (
            O => \N__49341\,
            I => \N__49335\
        );

    \I__11668\ : LocalMux
    port map (
            O => \N__49338\,
            I => \N__49332\
        );

    \I__11667\ : Span4Mux_v
    port map (
            O => \N__49335\,
            I => \N__49327\
        );

    \I__11666\ : Span4Mux_h
    port map (
            O => \N__49332\,
            I => \N__49327\
        );

    \I__11665\ : Odrv4
    port map (
            O => \N__49327\,
            I => comm_length_1
        );

    \I__11664\ : InMux
    port map (
            O => \N__49324\,
            I => \N__49320\
        );

    \I__11663\ : InMux
    port map (
            O => \N__49323\,
            I => \N__49317\
        );

    \I__11662\ : LocalMux
    port map (
            O => \N__49320\,
            I => \N__49314\
        );

    \I__11661\ : LocalMux
    port map (
            O => \N__49317\,
            I => \N__49311\
        );

    \I__11660\ : Span4Mux_v
    port map (
            O => \N__49314\,
            I => \N__49306\
        );

    \I__11659\ : Span4Mux_h
    port map (
            O => \N__49311\,
            I => \N__49306\
        );

    \I__11658\ : Odrv4
    port map (
            O => \N__49306\,
            I => n4_adj_1576
        );

    \I__11657\ : InMux
    port map (
            O => \N__49303\,
            I => \N__49299\
        );

    \I__11656\ : InMux
    port map (
            O => \N__49302\,
            I => \N__49295\
        );

    \I__11655\ : LocalMux
    port map (
            O => \N__49299\,
            I => \N__49292\
        );

    \I__11654\ : InMux
    port map (
            O => \N__49298\,
            I => \N__49289\
        );

    \I__11653\ : LocalMux
    port map (
            O => \N__49295\,
            I => \N__49281\
        );

    \I__11652\ : Span4Mux_v
    port map (
            O => \N__49292\,
            I => \N__49281\
        );

    \I__11651\ : LocalMux
    port map (
            O => \N__49289\,
            I => \N__49281\
        );

    \I__11650\ : InMux
    port map (
            O => \N__49288\,
            I => \N__49278\
        );

    \I__11649\ : Span4Mux_h
    port map (
            O => \N__49281\,
            I => \N__49275\
        );

    \I__11648\ : LocalMux
    port map (
            O => \N__49278\,
            I => comm_cmd_7
        );

    \I__11647\ : Odrv4
    port map (
            O => \N__49275\,
            I => comm_cmd_7
        );

    \I__11646\ : CascadeMux
    port map (
            O => \N__49270\,
            I => \n5_cascade_\
        );

    \I__11645\ : IoInMux
    port map (
            O => \N__49267\,
            I => \N__49264\
        );

    \I__11644\ : LocalMux
    port map (
            O => \N__49264\,
            I => \N__49261\
        );

    \I__11643\ : Span4Mux_s1_h
    port map (
            O => \N__49261\,
            I => \N__49258\
        );

    \I__11642\ : Sp12to4
    port map (
            O => \N__49258\,
            I => \N__49255\
        );

    \I__11641\ : Span12Mux_v
    port map (
            O => \N__49255\,
            I => \N__49252\
        );

    \I__11640\ : Odrv12
    port map (
            O => \N__49252\,
            I => \ICE_GPMI_0\
        );

    \I__11639\ : CEMux
    port map (
            O => \N__49249\,
            I => \N__49246\
        );

    \I__11638\ : LocalMux
    port map (
            O => \N__49246\,
            I => \N__49243\
        );

    \I__11637\ : Odrv4
    port map (
            O => \N__49243\,
            I => n11406
        );

    \I__11636\ : InMux
    port map (
            O => \N__49240\,
            I => \N__49232\
        );

    \I__11635\ : InMux
    port map (
            O => \N__49239\,
            I => \N__49229\
        );

    \I__11634\ : InMux
    port map (
            O => \N__49238\,
            I => \N__49226\
        );

    \I__11633\ : InMux
    port map (
            O => \N__49237\,
            I => \N__49223\
        );

    \I__11632\ : InMux
    port map (
            O => \N__49236\,
            I => \N__49220\
        );

    \I__11631\ : CascadeMux
    port map (
            O => \N__49235\,
            I => \N__49217\
        );

    \I__11630\ : LocalMux
    port map (
            O => \N__49232\,
            I => \N__49212\
        );

    \I__11629\ : LocalMux
    port map (
            O => \N__49229\,
            I => \N__49207\
        );

    \I__11628\ : LocalMux
    port map (
            O => \N__49226\,
            I => \N__49200\
        );

    \I__11627\ : LocalMux
    port map (
            O => \N__49223\,
            I => \N__49200\
        );

    \I__11626\ : LocalMux
    port map (
            O => \N__49220\,
            I => \N__49200\
        );

    \I__11625\ : InMux
    port map (
            O => \N__49217\,
            I => \N__49193\
        );

    \I__11624\ : InMux
    port map (
            O => \N__49216\,
            I => \N__49193\
        );

    \I__11623\ : InMux
    port map (
            O => \N__49215\,
            I => \N__49193\
        );

    \I__11622\ : Span4Mux_h
    port map (
            O => \N__49212\,
            I => \N__49190\
        );

    \I__11621\ : InMux
    port map (
            O => \N__49211\,
            I => \N__49187\
        );

    \I__11620\ : InMux
    port map (
            O => \N__49210\,
            I => \N__49182\
        );

    \I__11619\ : Sp12to4
    port map (
            O => \N__49207\,
            I => \N__49179\
        );

    \I__11618\ : Span4Mux_v
    port map (
            O => \N__49200\,
            I => \N__49176\
        );

    \I__11617\ : LocalMux
    port map (
            O => \N__49193\,
            I => \N__49169\
        );

    \I__11616\ : Span4Mux_v
    port map (
            O => \N__49190\,
            I => \N__49169\
        );

    \I__11615\ : LocalMux
    port map (
            O => \N__49187\,
            I => \N__49169\
        );

    \I__11614\ : InMux
    port map (
            O => \N__49186\,
            I => \N__49164\
        );

    \I__11613\ : InMux
    port map (
            O => \N__49185\,
            I => \N__49164\
        );

    \I__11612\ : LocalMux
    port map (
            O => \N__49182\,
            I => \N__49159\
        );

    \I__11611\ : Span12Mux_v
    port map (
            O => \N__49179\,
            I => \N__49159\
        );

    \I__11610\ : Span4Mux_h
    port map (
            O => \N__49176\,
            I => \N__49154\
        );

    \I__11609\ : Span4Mux_v
    port map (
            O => \N__49169\,
            I => \N__49154\
        );

    \I__11608\ : LocalMux
    port map (
            O => \N__49164\,
            I => n12220
        );

    \I__11607\ : Odrv12
    port map (
            O => \N__49159\,
            I => n12220
        );

    \I__11606\ : Odrv4
    port map (
            O => \N__49154\,
            I => n12220
        );

    \I__11605\ : CascadeMux
    port map (
            O => \N__49147\,
            I => \n10_adj_1572_cascade_\
        );

    \I__11604\ : CascadeMux
    port map (
            O => \N__49144\,
            I => \N__49141\
        );

    \I__11603\ : InMux
    port map (
            O => \N__49141\,
            I => \N__49135\
        );

    \I__11602\ : InMux
    port map (
            O => \N__49140\,
            I => \N__49135\
        );

    \I__11601\ : LocalMux
    port map (
            O => \N__49135\,
            I => \N__49132\
        );

    \I__11600\ : Span4Mux_h
    port map (
            O => \N__49132\,
            I => \N__49129\
        );

    \I__11599\ : Odrv4
    port map (
            O => \N__49129\,
            I => n20643
        );

    \I__11598\ : InMux
    port map (
            O => \N__49126\,
            I => \N__49123\
        );

    \I__11597\ : LocalMux
    port map (
            O => \N__49123\,
            I => n4_adj_1596
        );

    \I__11596\ : InMux
    port map (
            O => \N__49120\,
            I => \N__49117\
        );

    \I__11595\ : LocalMux
    port map (
            O => \N__49117\,
            I => \N__49114\
        );

    \I__11594\ : Span4Mux_h
    port map (
            O => \N__49114\,
            I => \N__49110\
        );

    \I__11593\ : InMux
    port map (
            O => \N__49113\,
            I => \N__49107\
        );

    \I__11592\ : Odrv4
    port map (
            O => \N__49110\,
            I => n2342
        );

    \I__11591\ : LocalMux
    port map (
            O => \N__49107\,
            I => n2342
        );

    \I__11590\ : CEMux
    port map (
            O => \N__49102\,
            I => \N__49099\
        );

    \I__11589\ : LocalMux
    port map (
            O => \N__49099\,
            I => \N__49096\
        );

    \I__11588\ : Odrv12
    port map (
            O => \N__49096\,
            I => n11836
        );

    \I__11587\ : SRMux
    port map (
            O => \N__49093\,
            I => \N__49090\
        );

    \I__11586\ : LocalMux
    port map (
            O => \N__49090\,
            I => \N__49087\
        );

    \I__11585\ : Span4Mux_h
    port map (
            O => \N__49087\,
            I => \N__49084\
        );

    \I__11584\ : Span4Mux_h
    port map (
            O => \N__49084\,
            I => \N__49081\
        );

    \I__11583\ : Odrv4
    port map (
            O => \N__49081\,
            I => n14722
        );

    \I__11582\ : InMux
    port map (
            O => \N__49078\,
            I => \N__49074\
        );

    \I__11581\ : InMux
    port map (
            O => \N__49077\,
            I => \N__49071\
        );

    \I__11580\ : LocalMux
    port map (
            O => \N__49074\,
            I => \N__49067\
        );

    \I__11579\ : LocalMux
    port map (
            O => \N__49071\,
            I => \N__49064\
        );

    \I__11578\ : InMux
    port map (
            O => \N__49070\,
            I => \N__49061\
        );

    \I__11577\ : Span4Mux_h
    port map (
            O => \N__49067\,
            I => \N__49058\
        );

    \I__11576\ : Span4Mux_h
    port map (
            O => \N__49064\,
            I => \N__49055\
        );

    \I__11575\ : LocalMux
    port map (
            O => \N__49061\,
            I => buf_adcdata_iac_5
        );

    \I__11574\ : Odrv4
    port map (
            O => \N__49058\,
            I => buf_adcdata_iac_5
        );

    \I__11573\ : Odrv4
    port map (
            O => \N__49055\,
            I => buf_adcdata_iac_5
        );

    \I__11572\ : CascadeMux
    port map (
            O => \N__49048\,
            I => \N__49045\
        );

    \I__11571\ : InMux
    port map (
            O => \N__49045\,
            I => \N__49042\
        );

    \I__11570\ : LocalMux
    port map (
            O => \N__49042\,
            I => \N__49038\
        );

    \I__11569\ : CascadeMux
    port map (
            O => \N__49041\,
            I => \N__49035\
        );

    \I__11568\ : Span4Mux_v
    port map (
            O => \N__49038\,
            I => \N__49032\
        );

    \I__11567\ : InMux
    port map (
            O => \N__49035\,
            I => \N__49029\
        );

    \I__11566\ : Sp12to4
    port map (
            O => \N__49032\,
            I => \N__49026\
        );

    \I__11565\ : LocalMux
    port map (
            O => \N__49029\,
            I => \N__49022\
        );

    \I__11564\ : Span12Mux_h
    port map (
            O => \N__49026\,
            I => \N__49019\
        );

    \I__11563\ : InMux
    port map (
            O => \N__49025\,
            I => \N__49016\
        );

    \I__11562\ : Odrv4
    port map (
            O => \N__49022\,
            I => cmd_rdadctmp_11
        );

    \I__11561\ : Odrv12
    port map (
            O => \N__49019\,
            I => cmd_rdadctmp_11
        );

    \I__11560\ : LocalMux
    port map (
            O => \N__49016\,
            I => cmd_rdadctmp_11
        );

    \I__11559\ : InMux
    port map (
            O => \N__49009\,
            I => \N__49005\
        );

    \I__11558\ : InMux
    port map (
            O => \N__49008\,
            I => \N__49001\
        );

    \I__11557\ : LocalMux
    port map (
            O => \N__49005\,
            I => \N__48994\
        );

    \I__11556\ : InMux
    port map (
            O => \N__49004\,
            I => \N__48991\
        );

    \I__11555\ : LocalMux
    port map (
            O => \N__49001\,
            I => \N__48987\
        );

    \I__11554\ : InMux
    port map (
            O => \N__49000\,
            I => \N__48984\
        );

    \I__11553\ : InMux
    port map (
            O => \N__48999\,
            I => \N__48979\
        );

    \I__11552\ : InMux
    port map (
            O => \N__48998\,
            I => \N__48979\
        );

    \I__11551\ : InMux
    port map (
            O => \N__48997\,
            I => \N__48976\
        );

    \I__11550\ : Span4Mux_v
    port map (
            O => \N__48994\,
            I => \N__48970\
        );

    \I__11549\ : LocalMux
    port map (
            O => \N__48991\,
            I => \N__48970\
        );

    \I__11548\ : InMux
    port map (
            O => \N__48990\,
            I => \N__48963\
        );

    \I__11547\ : Span4Mux_h
    port map (
            O => \N__48987\,
            I => \N__48954\
        );

    \I__11546\ : LocalMux
    port map (
            O => \N__48984\,
            I => \N__48954\
        );

    \I__11545\ : LocalMux
    port map (
            O => \N__48979\,
            I => \N__48948\
        );

    \I__11544\ : LocalMux
    port map (
            O => \N__48976\,
            I => \N__48948\
        );

    \I__11543\ : InMux
    port map (
            O => \N__48975\,
            I => \N__48945\
        );

    \I__11542\ : Span4Mux_h
    port map (
            O => \N__48970\,
            I => \N__48942\
        );

    \I__11541\ : InMux
    port map (
            O => \N__48969\,
            I => \N__48939\
        );

    \I__11540\ : InMux
    port map (
            O => \N__48968\,
            I => \N__48936\
        );

    \I__11539\ : InMux
    port map (
            O => \N__48967\,
            I => \N__48931\
        );

    \I__11538\ : InMux
    port map (
            O => \N__48966\,
            I => \N__48931\
        );

    \I__11537\ : LocalMux
    port map (
            O => \N__48963\,
            I => \N__48928\
        );

    \I__11536\ : InMux
    port map (
            O => \N__48962\,
            I => \N__48923\
        );

    \I__11535\ : InMux
    port map (
            O => \N__48961\,
            I => \N__48923\
        );

    \I__11534\ : InMux
    port map (
            O => \N__48960\,
            I => \N__48918\
        );

    \I__11533\ : InMux
    port map (
            O => \N__48959\,
            I => \N__48918\
        );

    \I__11532\ : Span4Mux_v
    port map (
            O => \N__48954\,
            I => \N__48915\
        );

    \I__11531\ : InMux
    port map (
            O => \N__48953\,
            I => \N__48912\
        );

    \I__11530\ : Span4Mux_h
    port map (
            O => \N__48948\,
            I => \N__48905\
        );

    \I__11529\ : LocalMux
    port map (
            O => \N__48945\,
            I => \N__48905\
        );

    \I__11528\ : Span4Mux_h
    port map (
            O => \N__48942\,
            I => \N__48898\
        );

    \I__11527\ : LocalMux
    port map (
            O => \N__48939\,
            I => \N__48898\
        );

    \I__11526\ : LocalMux
    port map (
            O => \N__48936\,
            I => \N__48898\
        );

    \I__11525\ : LocalMux
    port map (
            O => \N__48931\,
            I => \N__48895\
        );

    \I__11524\ : Span4Mux_v
    port map (
            O => \N__48928\,
            I => \N__48887\
        );

    \I__11523\ : LocalMux
    port map (
            O => \N__48923\,
            I => \N__48887\
        );

    \I__11522\ : LocalMux
    port map (
            O => \N__48918\,
            I => \N__48884\
        );

    \I__11521\ : Span4Mux_h
    port map (
            O => \N__48915\,
            I => \N__48879\
        );

    \I__11520\ : LocalMux
    port map (
            O => \N__48912\,
            I => \N__48879\
        );

    \I__11519\ : InMux
    port map (
            O => \N__48911\,
            I => \N__48874\
        );

    \I__11518\ : InMux
    port map (
            O => \N__48910\,
            I => \N__48874\
        );

    \I__11517\ : Span4Mux_v
    port map (
            O => \N__48905\,
            I => \N__48870\
        );

    \I__11516\ : Span4Mux_h
    port map (
            O => \N__48898\,
            I => \N__48867\
        );

    \I__11515\ : Span4Mux_h
    port map (
            O => \N__48895\,
            I => \N__48864\
        );

    \I__11514\ : InMux
    port map (
            O => \N__48894\,
            I => \N__48859\
        );

    \I__11513\ : InMux
    port map (
            O => \N__48893\,
            I => \N__48859\
        );

    \I__11512\ : InMux
    port map (
            O => \N__48892\,
            I => \N__48856\
        );

    \I__11511\ : Span4Mux_v
    port map (
            O => \N__48887\,
            I => \N__48847\
        );

    \I__11510\ : Span4Mux_v
    port map (
            O => \N__48884\,
            I => \N__48847\
        );

    \I__11509\ : Span4Mux_h
    port map (
            O => \N__48879\,
            I => \N__48847\
        );

    \I__11508\ : LocalMux
    port map (
            O => \N__48874\,
            I => \N__48847\
        );

    \I__11507\ : InMux
    port map (
            O => \N__48873\,
            I => \N__48844\
        );

    \I__11506\ : Odrv4
    port map (
            O => \N__48870\,
            I => n20543
        );

    \I__11505\ : Odrv4
    port map (
            O => \N__48867\,
            I => n20543
        );

    \I__11504\ : Odrv4
    port map (
            O => \N__48864\,
            I => n20543
        );

    \I__11503\ : LocalMux
    port map (
            O => \N__48859\,
            I => n20543
        );

    \I__11502\ : LocalMux
    port map (
            O => \N__48856\,
            I => n20543
        );

    \I__11501\ : Odrv4
    port map (
            O => \N__48847\,
            I => n20543
        );

    \I__11500\ : LocalMux
    port map (
            O => \N__48844\,
            I => n20543
        );

    \I__11499\ : InMux
    port map (
            O => \N__48829\,
            I => \N__48825\
        );

    \I__11498\ : InMux
    port map (
            O => \N__48828\,
            I => \N__48822\
        );

    \I__11497\ : LocalMux
    port map (
            O => \N__48825\,
            I => \N__48818\
        );

    \I__11496\ : LocalMux
    port map (
            O => \N__48822\,
            I => \N__48815\
        );

    \I__11495\ : InMux
    port map (
            O => \N__48821\,
            I => \N__48812\
        );

    \I__11494\ : Span4Mux_h
    port map (
            O => \N__48818\,
            I => \N__48809\
        );

    \I__11493\ : Span4Mux_h
    port map (
            O => \N__48815\,
            I => \N__48806\
        );

    \I__11492\ : LocalMux
    port map (
            O => \N__48812\,
            I => buf_adcdata_iac_4
        );

    \I__11491\ : Odrv4
    port map (
            O => \N__48809\,
            I => buf_adcdata_iac_4
        );

    \I__11490\ : Odrv4
    port map (
            O => \N__48806\,
            I => buf_adcdata_iac_4
        );

    \I__11489\ : CascadeMux
    port map (
            O => \N__48799\,
            I => \N__48795\
        );

    \I__11488\ : InMux
    port map (
            O => \N__48798\,
            I => \N__48792\
        );

    \I__11487\ : InMux
    port map (
            O => \N__48795\,
            I => \N__48789\
        );

    \I__11486\ : LocalMux
    port map (
            O => \N__48792\,
            I => \N__48786\
        );

    \I__11485\ : LocalMux
    port map (
            O => \N__48789\,
            I => \N__48782\
        );

    \I__11484\ : Span4Mux_v
    port map (
            O => \N__48786\,
            I => \N__48779\
        );

    \I__11483\ : InMux
    port map (
            O => \N__48785\,
            I => \N__48776\
        );

    \I__11482\ : Odrv12
    port map (
            O => \N__48782\,
            I => cmd_rdadctmp_14
        );

    \I__11481\ : Odrv4
    port map (
            O => \N__48779\,
            I => cmd_rdadctmp_14
        );

    \I__11480\ : LocalMux
    port map (
            O => \N__48776\,
            I => cmd_rdadctmp_14
        );

    \I__11479\ : InMux
    port map (
            O => \N__48769\,
            I => \N__48766\
        );

    \I__11478\ : LocalMux
    port map (
            O => \N__48766\,
            I => \N__48763\
        );

    \I__11477\ : Odrv4
    port map (
            O => \N__48763\,
            I => \comm_spi.n14581\
        );

    \I__11476\ : SRMux
    port map (
            O => \N__48760\,
            I => \N__48757\
        );

    \I__11475\ : LocalMux
    port map (
            O => \N__48757\,
            I => \N__48754\
        );

    \I__11474\ : Span4Mux_h
    port map (
            O => \N__48754\,
            I => \N__48751\
        );

    \I__11473\ : Odrv4
    port map (
            O => \N__48751\,
            I => \comm_spi.iclk_N_754\
        );

    \I__11472\ : InMux
    port map (
            O => \N__48748\,
            I => \N__48745\
        );

    \I__11471\ : LocalMux
    port map (
            O => \N__48745\,
            I => \N__48741\
        );

    \I__11470\ : InMux
    port map (
            O => \N__48744\,
            I => \N__48738\
        );

    \I__11469\ : Span4Mux_v
    port map (
            O => \N__48741\,
            I => \N__48734\
        );

    \I__11468\ : LocalMux
    port map (
            O => \N__48738\,
            I => \N__48731\
        );

    \I__11467\ : InMux
    port map (
            O => \N__48737\,
            I => \N__48728\
        );

    \I__11466\ : Sp12to4
    port map (
            O => \N__48734\,
            I => \N__48725\
        );

    \I__11465\ : Span4Mux_h
    port map (
            O => \N__48731\,
            I => \N__48720\
        );

    \I__11464\ : LocalMux
    port map (
            O => \N__48728\,
            I => \N__48720\
        );

    \I__11463\ : Span12Mux_h
    port map (
            O => \N__48725\,
            I => \N__48717\
        );

    \I__11462\ : Span4Mux_v
    port map (
            O => \N__48720\,
            I => \N__48714\
        );

    \I__11461\ : Odrv12
    port map (
            O => \N__48717\,
            I => comm_tx_buf_5
        );

    \I__11460\ : Odrv4
    port map (
            O => \N__48714\,
            I => comm_tx_buf_5
        );

    \I__11459\ : SRMux
    port map (
            O => \N__48709\,
            I => \N__48706\
        );

    \I__11458\ : LocalMux
    port map (
            O => \N__48706\,
            I => \N__48703\
        );

    \I__11457\ : Odrv12
    port map (
            O => \N__48703\,
            I => \comm_spi.data_tx_7__N_760\
        );

    \I__11456\ : InMux
    port map (
            O => \N__48700\,
            I => \N__48696\
        );

    \I__11455\ : InMux
    port map (
            O => \N__48699\,
            I => \N__48693\
        );

    \I__11454\ : LocalMux
    port map (
            O => \N__48696\,
            I => data_cntvec_14
        );

    \I__11453\ : LocalMux
    port map (
            O => \N__48693\,
            I => data_cntvec_14
        );

    \I__11452\ : InMux
    port map (
            O => \N__48688\,
            I => n19309
        );

    \I__11451\ : InMux
    port map (
            O => \N__48685\,
            I => n19310
        );

    \I__11450\ : InMux
    port map (
            O => \N__48682\,
            I => \N__48678\
        );

    \I__11449\ : InMux
    port map (
            O => \N__48681\,
            I => \N__48675\
        );

    \I__11448\ : LocalMux
    port map (
            O => \N__48678\,
            I => \N__48672\
        );

    \I__11447\ : LocalMux
    port map (
            O => \N__48675\,
            I => data_cntvec_15
        );

    \I__11446\ : Odrv4
    port map (
            O => \N__48672\,
            I => data_cntvec_15
        );

    \I__11445\ : CEMux
    port map (
            O => \N__48667\,
            I => \N__48664\
        );

    \I__11444\ : LocalMux
    port map (
            O => \N__48664\,
            I => \N__48659\
        );

    \I__11443\ : CEMux
    port map (
            O => \N__48663\,
            I => \N__48656\
        );

    \I__11442\ : CEMux
    port map (
            O => \N__48662\,
            I => \N__48652\
        );

    \I__11441\ : Span4Mux_h
    port map (
            O => \N__48659\,
            I => \N__48649\
        );

    \I__11440\ : LocalMux
    port map (
            O => \N__48656\,
            I => \N__48646\
        );

    \I__11439\ : CEMux
    port map (
            O => \N__48655\,
            I => \N__48643\
        );

    \I__11438\ : LocalMux
    port map (
            O => \N__48652\,
            I => \N__48640\
        );

    \I__11437\ : Span4Mux_v
    port map (
            O => \N__48649\,
            I => \N__48635\
        );

    \I__11436\ : Span4Mux_v
    port map (
            O => \N__48646\,
            I => \N__48635\
        );

    \I__11435\ : LocalMux
    port map (
            O => \N__48643\,
            I => \N__48632\
        );

    \I__11434\ : Span4Mux_h
    port map (
            O => \N__48640\,
            I => \N__48628\
        );

    \I__11433\ : Span4Mux_h
    port map (
            O => \N__48635\,
            I => \N__48623\
        );

    \I__11432\ : Span4Mux_h
    port map (
            O => \N__48632\,
            I => \N__48623\
        );

    \I__11431\ : InMux
    port map (
            O => \N__48631\,
            I => \N__48620\
        );

    \I__11430\ : Span4Mux_h
    port map (
            O => \N__48628\,
            I => \N__48617\
        );

    \I__11429\ : Span4Mux_h
    port map (
            O => \N__48623\,
            I => \N__48614\
        );

    \I__11428\ : LocalMux
    port map (
            O => \N__48620\,
            I => \N__48611\
        );

    \I__11427\ : Odrv4
    port map (
            O => \N__48617\,
            I => n13443
        );

    \I__11426\ : Odrv4
    port map (
            O => \N__48614\,
            I => n13443
        );

    \I__11425\ : Odrv12
    port map (
            O => \N__48611\,
            I => n13443
        );

    \I__11424\ : SRMux
    port map (
            O => \N__48604\,
            I => \N__48600\
        );

    \I__11423\ : SRMux
    port map (
            O => \N__48603\,
            I => \N__48597\
        );

    \I__11422\ : LocalMux
    port map (
            O => \N__48600\,
            I => \N__48593\
        );

    \I__11421\ : LocalMux
    port map (
            O => \N__48597\,
            I => \N__48590\
        );

    \I__11420\ : SRMux
    port map (
            O => \N__48596\,
            I => \N__48587\
        );

    \I__11419\ : Span4Mux_h
    port map (
            O => \N__48593\,
            I => \N__48583\
        );

    \I__11418\ : Span4Mux_v
    port map (
            O => \N__48590\,
            I => \N__48580\
        );

    \I__11417\ : LocalMux
    port map (
            O => \N__48587\,
            I => \N__48577\
        );

    \I__11416\ : SRMux
    port map (
            O => \N__48586\,
            I => \N__48574\
        );

    \I__11415\ : Odrv4
    port map (
            O => \N__48583\,
            I => n14632
        );

    \I__11414\ : Odrv4
    port map (
            O => \N__48580\,
            I => n14632
        );

    \I__11413\ : Odrv12
    port map (
            O => \N__48577\,
            I => n14632
        );

    \I__11412\ : LocalMux
    port map (
            O => \N__48574\,
            I => n14632
        );

    \I__11411\ : InMux
    port map (
            O => \N__48565\,
            I => \N__48561\
        );

    \I__11410\ : InMux
    port map (
            O => \N__48564\,
            I => \N__48558\
        );

    \I__11409\ : LocalMux
    port map (
            O => \N__48561\,
            I => \N__48554\
        );

    \I__11408\ : LocalMux
    port map (
            O => \N__48558\,
            I => \N__48551\
        );

    \I__11407\ : InMux
    port map (
            O => \N__48557\,
            I => \N__48548\
        );

    \I__11406\ : Span4Mux_v
    port map (
            O => \N__48554\,
            I => \N__48545\
        );

    \I__11405\ : Span4Mux_h
    port map (
            O => \N__48551\,
            I => \N__48542\
        );

    \I__11404\ : LocalMux
    port map (
            O => \N__48548\,
            I => buf_adcdata_iac_6
        );

    \I__11403\ : Odrv4
    port map (
            O => \N__48545\,
            I => buf_adcdata_iac_6
        );

    \I__11402\ : Odrv4
    port map (
            O => \N__48542\,
            I => buf_adcdata_iac_6
        );

    \I__11401\ : InMux
    port map (
            O => \N__48535\,
            I => \N__48530\
        );

    \I__11400\ : InMux
    port map (
            O => \N__48534\,
            I => \N__48527\
        );

    \I__11399\ : CascadeMux
    port map (
            O => \N__48533\,
            I => \N__48521\
        );

    \I__11398\ : LocalMux
    port map (
            O => \N__48530\,
            I => \N__48518\
        );

    \I__11397\ : LocalMux
    port map (
            O => \N__48527\,
            I => \N__48515\
        );

    \I__11396\ : InMux
    port map (
            O => \N__48526\,
            I => \N__48512\
        );

    \I__11395\ : InMux
    port map (
            O => \N__48525\,
            I => \N__48499\
        );

    \I__11394\ : InMux
    port map (
            O => \N__48524\,
            I => \N__48499\
        );

    \I__11393\ : InMux
    port map (
            O => \N__48521\,
            I => \N__48496\
        );

    \I__11392\ : Span4Mux_h
    port map (
            O => \N__48518\,
            I => \N__48489\
        );

    \I__11391\ : Span4Mux_h
    port map (
            O => \N__48515\,
            I => \N__48484\
        );

    \I__11390\ : LocalMux
    port map (
            O => \N__48512\,
            I => \N__48484\
        );

    \I__11389\ : CascadeMux
    port map (
            O => \N__48511\,
            I => \N__48481\
        );

    \I__11388\ : InMux
    port map (
            O => \N__48510\,
            I => \N__48469\
        );

    \I__11387\ : InMux
    port map (
            O => \N__48509\,
            I => \N__48469\
        );

    \I__11386\ : InMux
    port map (
            O => \N__48508\,
            I => \N__48469\
        );

    \I__11385\ : InMux
    port map (
            O => \N__48507\,
            I => \N__48469\
        );

    \I__11384\ : InMux
    port map (
            O => \N__48506\,
            I => \N__48464\
        );

    \I__11383\ : InMux
    port map (
            O => \N__48505\,
            I => \N__48464\
        );

    \I__11382\ : InMux
    port map (
            O => \N__48504\,
            I => \N__48461\
        );

    \I__11381\ : LocalMux
    port map (
            O => \N__48499\,
            I => \N__48456\
        );

    \I__11380\ : LocalMux
    port map (
            O => \N__48496\,
            I => \N__48456\
        );

    \I__11379\ : InMux
    port map (
            O => \N__48495\,
            I => \N__48453\
        );

    \I__11378\ : InMux
    port map (
            O => \N__48494\,
            I => \N__48448\
        );

    \I__11377\ : InMux
    port map (
            O => \N__48493\,
            I => \N__48448\
        );

    \I__11376\ : InMux
    port map (
            O => \N__48492\,
            I => \N__48445\
        );

    \I__11375\ : Span4Mux_h
    port map (
            O => \N__48489\,
            I => \N__48440\
        );

    \I__11374\ : Span4Mux_h
    port map (
            O => \N__48484\,
            I => \N__48440\
        );

    \I__11373\ : InMux
    port map (
            O => \N__48481\,
            I => \N__48432\
        );

    \I__11372\ : InMux
    port map (
            O => \N__48480\,
            I => \N__48432\
        );

    \I__11371\ : InMux
    port map (
            O => \N__48479\,
            I => \N__48427\
        );

    \I__11370\ : InMux
    port map (
            O => \N__48478\,
            I => \N__48427\
        );

    \I__11369\ : LocalMux
    port map (
            O => \N__48469\,
            I => \N__48422\
        );

    \I__11368\ : LocalMux
    port map (
            O => \N__48464\,
            I => \N__48422\
        );

    \I__11367\ : LocalMux
    port map (
            O => \N__48461\,
            I => \N__48419\
        );

    \I__11366\ : Span4Mux_h
    port map (
            O => \N__48456\,
            I => \N__48416\
        );

    \I__11365\ : LocalMux
    port map (
            O => \N__48453\,
            I => \N__48413\
        );

    \I__11364\ : LocalMux
    port map (
            O => \N__48448\,
            I => \N__48408\
        );

    \I__11363\ : LocalMux
    port map (
            O => \N__48445\,
            I => \N__48408\
        );

    \I__11362\ : Span4Mux_h
    port map (
            O => \N__48440\,
            I => \N__48405\
        );

    \I__11361\ : InMux
    port map (
            O => \N__48439\,
            I => \N__48402\
        );

    \I__11360\ : InMux
    port map (
            O => \N__48438\,
            I => \N__48399\
        );

    \I__11359\ : InMux
    port map (
            O => \N__48437\,
            I => \N__48396\
        );

    \I__11358\ : LocalMux
    port map (
            O => \N__48432\,
            I => \N__48389\
        );

    \I__11357\ : LocalMux
    port map (
            O => \N__48427\,
            I => \N__48389\
        );

    \I__11356\ : Span4Mux_h
    port map (
            O => \N__48422\,
            I => \N__48389\
        );

    \I__11355\ : Span12Mux_h
    port map (
            O => \N__48419\,
            I => \N__48386\
        );

    \I__11354\ : Span4Mux_v
    port map (
            O => \N__48416\,
            I => \N__48383\
        );

    \I__11353\ : Span4Mux_v
    port map (
            O => \N__48413\,
            I => \N__48378\
        );

    \I__11352\ : Span4Mux_h
    port map (
            O => \N__48408\,
            I => \N__48378\
        );

    \I__11351\ : Span4Mux_h
    port map (
            O => \N__48405\,
            I => \N__48375\
        );

    \I__11350\ : LocalMux
    port map (
            O => \N__48402\,
            I => n20540
        );

    \I__11349\ : LocalMux
    port map (
            O => \N__48399\,
            I => n20540
        );

    \I__11348\ : LocalMux
    port map (
            O => \N__48396\,
            I => n20540
        );

    \I__11347\ : Odrv4
    port map (
            O => \N__48389\,
            I => n20540
        );

    \I__11346\ : Odrv12
    port map (
            O => \N__48386\,
            I => n20540
        );

    \I__11345\ : Odrv4
    port map (
            O => \N__48383\,
            I => n20540
        );

    \I__11344\ : Odrv4
    port map (
            O => \N__48378\,
            I => n20540
        );

    \I__11343\ : Odrv4
    port map (
            O => \N__48375\,
            I => n20540
        );

    \I__11342\ : CascadeMux
    port map (
            O => \N__48358\,
            I => \N__48355\
        );

    \I__11341\ : InMux
    port map (
            O => \N__48355\,
            I => \N__48352\
        );

    \I__11340\ : LocalMux
    port map (
            O => \N__48352\,
            I => \N__48343\
        );

    \I__11339\ : InMux
    port map (
            O => \N__48351\,
            I => \N__48336\
        );

    \I__11338\ : InMux
    port map (
            O => \N__48350\,
            I => \N__48336\
        );

    \I__11337\ : InMux
    port map (
            O => \N__48349\,
            I => \N__48336\
        );

    \I__11336\ : InMux
    port map (
            O => \N__48348\,
            I => \N__48332\
        );

    \I__11335\ : InMux
    port map (
            O => \N__48347\,
            I => \N__48329\
        );

    \I__11334\ : CascadeMux
    port map (
            O => \N__48346\,
            I => \N__48326\
        );

    \I__11333\ : Span4Mux_h
    port map (
            O => \N__48343\,
            I => \N__48316\
        );

    \I__11332\ : LocalMux
    port map (
            O => \N__48336\,
            I => \N__48311\
        );

    \I__11331\ : CascadeMux
    port map (
            O => \N__48335\,
            I => \N__48308\
        );

    \I__11330\ : LocalMux
    port map (
            O => \N__48332\,
            I => \N__48305\
        );

    \I__11329\ : LocalMux
    port map (
            O => \N__48329\,
            I => \N__48302\
        );

    \I__11328\ : InMux
    port map (
            O => \N__48326\,
            I => \N__48293\
        );

    \I__11327\ : InMux
    port map (
            O => \N__48325\,
            I => \N__48293\
        );

    \I__11326\ : InMux
    port map (
            O => \N__48324\,
            I => \N__48293\
        );

    \I__11325\ : InMux
    port map (
            O => \N__48323\,
            I => \N__48293\
        );

    \I__11324\ : InMux
    port map (
            O => \N__48322\,
            I => \N__48288\
        );

    \I__11323\ : InMux
    port map (
            O => \N__48321\,
            I => \N__48288\
        );

    \I__11322\ : InMux
    port map (
            O => \N__48320\,
            I => \N__48275\
        );

    \I__11321\ : InMux
    port map (
            O => \N__48319\,
            I => \N__48275\
        );

    \I__11320\ : Span4Mux_h
    port map (
            O => \N__48316\,
            I => \N__48272\
        );

    \I__11319\ : InMux
    port map (
            O => \N__48315\,
            I => \N__48269\
        );

    \I__11318\ : InMux
    port map (
            O => \N__48314\,
            I => \N__48266\
        );

    \I__11317\ : Span4Mux_v
    port map (
            O => \N__48311\,
            I => \N__48259\
        );

    \I__11316\ : InMux
    port map (
            O => \N__48308\,
            I => \N__48256\
        );

    \I__11315\ : Span4Mux_v
    port map (
            O => \N__48305\,
            I => \N__48251\
        );

    \I__11314\ : Span4Mux_v
    port map (
            O => \N__48302\,
            I => \N__48251\
        );

    \I__11313\ : LocalMux
    port map (
            O => \N__48293\,
            I => \N__48248\
        );

    \I__11312\ : LocalMux
    port map (
            O => \N__48288\,
            I => \N__48245\
        );

    \I__11311\ : InMux
    port map (
            O => \N__48287\,
            I => \N__48242\
        );

    \I__11310\ : InMux
    port map (
            O => \N__48286\,
            I => \N__48235\
        );

    \I__11309\ : InMux
    port map (
            O => \N__48285\,
            I => \N__48235\
        );

    \I__11308\ : InMux
    port map (
            O => \N__48284\,
            I => \N__48235\
        );

    \I__11307\ : CascadeMux
    port map (
            O => \N__48283\,
            I => \N__48232\
        );

    \I__11306\ : CascadeMux
    port map (
            O => \N__48282\,
            I => \N__48229\
        );

    \I__11305\ : CascadeMux
    port map (
            O => \N__48281\,
            I => \N__48226\
        );

    \I__11304\ : CascadeMux
    port map (
            O => \N__48280\,
            I => \N__48220\
        );

    \I__11303\ : LocalMux
    port map (
            O => \N__48275\,
            I => \N__48209\
        );

    \I__11302\ : Span4Mux_v
    port map (
            O => \N__48272\,
            I => \N__48209\
        );

    \I__11301\ : LocalMux
    port map (
            O => \N__48269\,
            I => \N__48209\
        );

    \I__11300\ : LocalMux
    port map (
            O => \N__48266\,
            I => \N__48206\
        );

    \I__11299\ : CascadeMux
    port map (
            O => \N__48265\,
            I => \N__48199\
        );

    \I__11298\ : CascadeMux
    port map (
            O => \N__48264\,
            I => \N__48191\
        );

    \I__11297\ : CascadeMux
    port map (
            O => \N__48263\,
            I => \N__48188\
        );

    \I__11296\ : CascadeMux
    port map (
            O => \N__48262\,
            I => \N__48185\
        );

    \I__11295\ : Span4Mux_h
    port map (
            O => \N__48259\,
            I => \N__48166\
        );

    \I__11294\ : LocalMux
    port map (
            O => \N__48256\,
            I => \N__48166\
        );

    \I__11293\ : Span4Mux_h
    port map (
            O => \N__48251\,
            I => \N__48166\
        );

    \I__11292\ : Span4Mux_h
    port map (
            O => \N__48248\,
            I => \N__48157\
        );

    \I__11291\ : Span4Mux_h
    port map (
            O => \N__48245\,
            I => \N__48157\
        );

    \I__11290\ : LocalMux
    port map (
            O => \N__48242\,
            I => \N__48157\
        );

    \I__11289\ : LocalMux
    port map (
            O => \N__48235\,
            I => \N__48157\
        );

    \I__11288\ : InMux
    port map (
            O => \N__48232\,
            I => \N__48144\
        );

    \I__11287\ : InMux
    port map (
            O => \N__48229\,
            I => \N__48144\
        );

    \I__11286\ : InMux
    port map (
            O => \N__48226\,
            I => \N__48144\
        );

    \I__11285\ : InMux
    port map (
            O => \N__48225\,
            I => \N__48144\
        );

    \I__11284\ : InMux
    port map (
            O => \N__48224\,
            I => \N__48144\
        );

    \I__11283\ : InMux
    port map (
            O => \N__48223\,
            I => \N__48144\
        );

    \I__11282\ : InMux
    port map (
            O => \N__48220\,
            I => \N__48139\
        );

    \I__11281\ : InMux
    port map (
            O => \N__48219\,
            I => \N__48139\
        );

    \I__11280\ : InMux
    port map (
            O => \N__48218\,
            I => \N__48136\
        );

    \I__11279\ : InMux
    port map (
            O => \N__48217\,
            I => \N__48131\
        );

    \I__11278\ : InMux
    port map (
            O => \N__48216\,
            I => \N__48131\
        );

    \I__11277\ : Span4Mux_h
    port map (
            O => \N__48209\,
            I => \N__48128\
        );

    \I__11276\ : Span4Mux_h
    port map (
            O => \N__48206\,
            I => \N__48125\
        );

    \I__11275\ : InMux
    port map (
            O => \N__48205\,
            I => \N__48118\
        );

    \I__11274\ : InMux
    port map (
            O => \N__48204\,
            I => \N__48118\
        );

    \I__11273\ : InMux
    port map (
            O => \N__48203\,
            I => \N__48118\
        );

    \I__11272\ : CascadeMux
    port map (
            O => \N__48202\,
            I => \N__48114\
        );

    \I__11271\ : InMux
    port map (
            O => \N__48199\,
            I => \N__48109\
        );

    \I__11270\ : InMux
    port map (
            O => \N__48198\,
            I => \N__48098\
        );

    \I__11269\ : InMux
    port map (
            O => \N__48197\,
            I => \N__48098\
        );

    \I__11268\ : InMux
    port map (
            O => \N__48196\,
            I => \N__48098\
        );

    \I__11267\ : InMux
    port map (
            O => \N__48195\,
            I => \N__48098\
        );

    \I__11266\ : InMux
    port map (
            O => \N__48194\,
            I => \N__48098\
        );

    \I__11265\ : InMux
    port map (
            O => \N__48191\,
            I => \N__48081\
        );

    \I__11264\ : InMux
    port map (
            O => \N__48188\,
            I => \N__48081\
        );

    \I__11263\ : InMux
    port map (
            O => \N__48185\,
            I => \N__48081\
        );

    \I__11262\ : InMux
    port map (
            O => \N__48184\,
            I => \N__48081\
        );

    \I__11261\ : InMux
    port map (
            O => \N__48183\,
            I => \N__48081\
        );

    \I__11260\ : InMux
    port map (
            O => \N__48182\,
            I => \N__48081\
        );

    \I__11259\ : InMux
    port map (
            O => \N__48181\,
            I => \N__48081\
        );

    \I__11258\ : InMux
    port map (
            O => \N__48180\,
            I => \N__48081\
        );

    \I__11257\ : InMux
    port map (
            O => \N__48179\,
            I => \N__48076\
        );

    \I__11256\ : InMux
    port map (
            O => \N__48178\,
            I => \N__48076\
        );

    \I__11255\ : InMux
    port map (
            O => \N__48177\,
            I => \N__48065\
        );

    \I__11254\ : InMux
    port map (
            O => \N__48176\,
            I => \N__48065\
        );

    \I__11253\ : InMux
    port map (
            O => \N__48175\,
            I => \N__48065\
        );

    \I__11252\ : InMux
    port map (
            O => \N__48174\,
            I => \N__48065\
        );

    \I__11251\ : InMux
    port map (
            O => \N__48173\,
            I => \N__48065\
        );

    \I__11250\ : Span4Mux_h
    port map (
            O => \N__48166\,
            I => \N__48060\
        );

    \I__11249\ : Span4Mux_v
    port map (
            O => \N__48157\,
            I => \N__48060\
        );

    \I__11248\ : LocalMux
    port map (
            O => \N__48144\,
            I => \N__48051\
        );

    \I__11247\ : LocalMux
    port map (
            O => \N__48139\,
            I => \N__48051\
        );

    \I__11246\ : LocalMux
    port map (
            O => \N__48136\,
            I => \N__48051\
        );

    \I__11245\ : LocalMux
    port map (
            O => \N__48131\,
            I => \N__48051\
        );

    \I__11244\ : Span4Mux_v
    port map (
            O => \N__48128\,
            I => \N__48048\
        );

    \I__11243\ : Span4Mux_h
    port map (
            O => \N__48125\,
            I => \N__48043\
        );

    \I__11242\ : LocalMux
    port map (
            O => \N__48118\,
            I => \N__48043\
        );

    \I__11241\ : InMux
    port map (
            O => \N__48117\,
            I => \N__48032\
        );

    \I__11240\ : InMux
    port map (
            O => \N__48114\,
            I => \N__48025\
        );

    \I__11239\ : InMux
    port map (
            O => \N__48113\,
            I => \N__48025\
        );

    \I__11238\ : InMux
    port map (
            O => \N__48112\,
            I => \N__48025\
        );

    \I__11237\ : LocalMux
    port map (
            O => \N__48109\,
            I => \N__48018\
        );

    \I__11236\ : LocalMux
    port map (
            O => \N__48098\,
            I => \N__48018\
        );

    \I__11235\ : LocalMux
    port map (
            O => \N__48081\,
            I => \N__48018\
        );

    \I__11234\ : LocalMux
    port map (
            O => \N__48076\,
            I => \N__48013\
        );

    \I__11233\ : LocalMux
    port map (
            O => \N__48065\,
            I => \N__48013\
        );

    \I__11232\ : Sp12to4
    port map (
            O => \N__48060\,
            I => \N__48010\
        );

    \I__11231\ : Span4Mux_v
    port map (
            O => \N__48051\,
            I => \N__48003\
        );

    \I__11230\ : Span4Mux_h
    port map (
            O => \N__48048\,
            I => \N__48003\
        );

    \I__11229\ : Span4Mux_h
    port map (
            O => \N__48043\,
            I => \N__48003\
        );

    \I__11228\ : InMux
    port map (
            O => \N__48042\,
            I => \N__47994\
        );

    \I__11227\ : InMux
    port map (
            O => \N__48041\,
            I => \N__47994\
        );

    \I__11226\ : InMux
    port map (
            O => \N__48040\,
            I => \N__47994\
        );

    \I__11225\ : InMux
    port map (
            O => \N__48039\,
            I => \N__47994\
        );

    \I__11224\ : InMux
    port map (
            O => \N__48038\,
            I => \N__47985\
        );

    \I__11223\ : InMux
    port map (
            O => \N__48037\,
            I => \N__47985\
        );

    \I__11222\ : InMux
    port map (
            O => \N__48036\,
            I => \N__47985\
        );

    \I__11221\ : InMux
    port map (
            O => \N__48035\,
            I => \N__47985\
        );

    \I__11220\ : LocalMux
    port map (
            O => \N__48032\,
            I => adc_state_0_adj_1411
        );

    \I__11219\ : LocalMux
    port map (
            O => \N__48025\,
            I => adc_state_0_adj_1411
        );

    \I__11218\ : Odrv4
    port map (
            O => \N__48018\,
            I => adc_state_0_adj_1411
        );

    \I__11217\ : Odrv12
    port map (
            O => \N__48013\,
            I => adc_state_0_adj_1411
        );

    \I__11216\ : Odrv12
    port map (
            O => \N__48010\,
            I => adc_state_0_adj_1411
        );

    \I__11215\ : Odrv4
    port map (
            O => \N__48003\,
            I => adc_state_0_adj_1411
        );

    \I__11214\ : LocalMux
    port map (
            O => \N__47994\,
            I => adc_state_0_adj_1411
        );

    \I__11213\ : LocalMux
    port map (
            O => \N__47985\,
            I => adc_state_0_adj_1411
        );

    \I__11212\ : CascadeMux
    port map (
            O => \N__47968\,
            I => \N__47964\
        );

    \I__11211\ : InMux
    port map (
            O => \N__47967\,
            I => \N__47961\
        );

    \I__11210\ : InMux
    port map (
            O => \N__47964\,
            I => \N__47958\
        );

    \I__11209\ : LocalMux
    port map (
            O => \N__47961\,
            I => \N__47955\
        );

    \I__11208\ : LocalMux
    port map (
            O => \N__47958\,
            I => \N__47952\
        );

    \I__11207\ : Span4Mux_v
    port map (
            O => \N__47955\,
            I => \N__47949\
        );

    \I__11206\ : Span12Mux_v
    port map (
            O => \N__47952\,
            I => \N__47945\
        );

    \I__11205\ : Span4Mux_h
    port map (
            O => \N__47949\,
            I => \N__47942\
        );

    \I__11204\ : InMux
    port map (
            O => \N__47948\,
            I => \N__47939\
        );

    \I__11203\ : Odrv12
    port map (
            O => \N__47945\,
            I => cmd_rdadctmp_12_adj_1431
        );

    \I__11202\ : Odrv4
    port map (
            O => \N__47942\,
            I => cmd_rdadctmp_12_adj_1431
        );

    \I__11201\ : LocalMux
    port map (
            O => \N__47939\,
            I => cmd_rdadctmp_12_adj_1431
        );

    \I__11200\ : InMux
    port map (
            O => \N__47932\,
            I => \N__47929\
        );

    \I__11199\ : LocalMux
    port map (
            O => \N__47929\,
            I => \N__47925\
        );

    \I__11198\ : InMux
    port map (
            O => \N__47928\,
            I => \N__47921\
        );

    \I__11197\ : Span4Mux_v
    port map (
            O => \N__47925\,
            I => \N__47918\
        );

    \I__11196\ : InMux
    port map (
            O => \N__47924\,
            I => \N__47915\
        );

    \I__11195\ : LocalMux
    port map (
            O => \N__47921\,
            I => buf_adcdata_vac_7
        );

    \I__11194\ : Odrv4
    port map (
            O => \N__47918\,
            I => buf_adcdata_vac_7
        );

    \I__11193\ : LocalMux
    port map (
            O => \N__47915\,
            I => buf_adcdata_vac_7
        );

    \I__11192\ : InMux
    port map (
            O => \N__47908\,
            I => \N__47905\
        );

    \I__11191\ : LocalMux
    port map (
            O => \N__47905\,
            I => \N__47902\
        );

    \I__11190\ : Span4Mux_v
    port map (
            O => \N__47902\,
            I => \N__47899\
        );

    \I__11189\ : Span4Mux_v
    port map (
            O => \N__47899\,
            I => \N__47895\
        );

    \I__11188\ : CascadeMux
    port map (
            O => \N__47898\,
            I => \N__47892\
        );

    \I__11187\ : Sp12to4
    port map (
            O => \N__47895\,
            I => \N__47889\
        );

    \I__11186\ : InMux
    port map (
            O => \N__47892\,
            I => \N__47886\
        );

    \I__11185\ : Odrv12
    port map (
            O => \N__47889\,
            I => buf_adcdata_vdc_7
        );

    \I__11184\ : LocalMux
    port map (
            O => \N__47886\,
            I => buf_adcdata_vdc_7
        );

    \I__11183\ : InMux
    port map (
            O => \N__47881\,
            I => \N__47877\
        );

    \I__11182\ : CascadeMux
    port map (
            O => \N__47880\,
            I => \N__47874\
        );

    \I__11181\ : LocalMux
    port map (
            O => \N__47877\,
            I => \N__47870\
        );

    \I__11180\ : InMux
    port map (
            O => \N__47874\,
            I => \N__47867\
        );

    \I__11179\ : InMux
    port map (
            O => \N__47873\,
            I => \N__47864\
        );

    \I__11178\ : Span4Mux_h
    port map (
            O => \N__47870\,
            I => \N__47861\
        );

    \I__11177\ : LocalMux
    port map (
            O => \N__47867\,
            I => buf_adcdata_iac_7
        );

    \I__11176\ : LocalMux
    port map (
            O => \N__47864\,
            I => buf_adcdata_iac_7
        );

    \I__11175\ : Odrv4
    port map (
            O => \N__47861\,
            I => buf_adcdata_iac_7
        );

    \I__11174\ : CascadeMux
    port map (
            O => \N__47854\,
            I => \n19_adj_1589_cascade_\
        );

    \I__11173\ : InMux
    port map (
            O => \N__47851\,
            I => \N__47840\
        );

    \I__11172\ : InMux
    port map (
            O => \N__47850\,
            I => \N__47837\
        );

    \I__11171\ : CascadeMux
    port map (
            O => \N__47849\,
            I => \N__47826\
        );

    \I__11170\ : InMux
    port map (
            O => \N__47848\,
            I => \N__47817\
        );

    \I__11169\ : InMux
    port map (
            O => \N__47847\,
            I => \N__47814\
        );

    \I__11168\ : InMux
    port map (
            O => \N__47846\,
            I => \N__47811\
        );

    \I__11167\ : InMux
    port map (
            O => \N__47845\,
            I => \N__47806\
        );

    \I__11166\ : InMux
    port map (
            O => \N__47844\,
            I => \N__47806\
        );

    \I__11165\ : InMux
    port map (
            O => \N__47843\,
            I => \N__47803\
        );

    \I__11164\ : LocalMux
    port map (
            O => \N__47840\,
            I => \N__47800\
        );

    \I__11163\ : LocalMux
    port map (
            O => \N__47837\,
            I => \N__47797\
        );

    \I__11162\ : InMux
    port map (
            O => \N__47836\,
            I => \N__47794\
        );

    \I__11161\ : InMux
    port map (
            O => \N__47835\,
            I => \N__47791\
        );

    \I__11160\ : InMux
    port map (
            O => \N__47834\,
            I => \N__47775\
        );

    \I__11159\ : InMux
    port map (
            O => \N__47833\,
            I => \N__47771\
        );

    \I__11158\ : InMux
    port map (
            O => \N__47832\,
            I => \N__47768\
        );

    \I__11157\ : InMux
    port map (
            O => \N__47831\,
            I => \N__47763\
        );

    \I__11156\ : InMux
    port map (
            O => \N__47830\,
            I => \N__47763\
        );

    \I__11155\ : InMux
    port map (
            O => \N__47829\,
            I => \N__47758\
        );

    \I__11154\ : InMux
    port map (
            O => \N__47826\,
            I => \N__47758\
        );

    \I__11153\ : InMux
    port map (
            O => \N__47825\,
            I => \N__47755\
        );

    \I__11152\ : InMux
    port map (
            O => \N__47824\,
            I => \N__47749\
        );

    \I__11151\ : InMux
    port map (
            O => \N__47823\,
            I => \N__47738\
        );

    \I__11150\ : InMux
    port map (
            O => \N__47822\,
            I => \N__47734\
        );

    \I__11149\ : InMux
    port map (
            O => \N__47821\,
            I => \N__47731\
        );

    \I__11148\ : InMux
    port map (
            O => \N__47820\,
            I => \N__47728\
        );

    \I__11147\ : LocalMux
    port map (
            O => \N__47817\,
            I => \N__47721\
        );

    \I__11146\ : LocalMux
    port map (
            O => \N__47814\,
            I => \N__47721\
        );

    \I__11145\ : LocalMux
    port map (
            O => \N__47811\,
            I => \N__47718\
        );

    \I__11144\ : LocalMux
    port map (
            O => \N__47806\,
            I => \N__47705\
        );

    \I__11143\ : LocalMux
    port map (
            O => \N__47803\,
            I => \N__47705\
        );

    \I__11142\ : Span4Mux_v
    port map (
            O => \N__47800\,
            I => \N__47705\
        );

    \I__11141\ : Span4Mux_h
    port map (
            O => \N__47797\,
            I => \N__47705\
        );

    \I__11140\ : LocalMux
    port map (
            O => \N__47794\,
            I => \N__47705\
        );

    \I__11139\ : LocalMux
    port map (
            O => \N__47791\,
            I => \N__47705\
        );

    \I__11138\ : InMux
    port map (
            O => \N__47790\,
            I => \N__47702\
        );

    \I__11137\ : InMux
    port map (
            O => \N__47789\,
            I => \N__47691\
        );

    \I__11136\ : InMux
    port map (
            O => \N__47788\,
            I => \N__47688\
        );

    \I__11135\ : InMux
    port map (
            O => \N__47787\,
            I => \N__47683\
        );

    \I__11134\ : InMux
    port map (
            O => \N__47786\,
            I => \N__47683\
        );

    \I__11133\ : InMux
    port map (
            O => \N__47785\,
            I => \N__47674\
        );

    \I__11132\ : InMux
    port map (
            O => \N__47784\,
            I => \N__47674\
        );

    \I__11131\ : InMux
    port map (
            O => \N__47783\,
            I => \N__47674\
        );

    \I__11130\ : InMux
    port map (
            O => \N__47782\,
            I => \N__47674\
        );

    \I__11129\ : InMux
    port map (
            O => \N__47781\,
            I => \N__47665\
        );

    \I__11128\ : InMux
    port map (
            O => \N__47780\,
            I => \N__47665\
        );

    \I__11127\ : InMux
    port map (
            O => \N__47779\,
            I => \N__47665\
        );

    \I__11126\ : InMux
    port map (
            O => \N__47778\,
            I => \N__47665\
        );

    \I__11125\ : LocalMux
    port map (
            O => \N__47775\,
            I => \N__47662\
        );

    \I__11124\ : InMux
    port map (
            O => \N__47774\,
            I => \N__47659\
        );

    \I__11123\ : LocalMux
    port map (
            O => \N__47771\,
            I => \N__47654\
        );

    \I__11122\ : LocalMux
    port map (
            O => \N__47768\,
            I => \N__47654\
        );

    \I__11121\ : LocalMux
    port map (
            O => \N__47763\,
            I => \N__47649\
        );

    \I__11120\ : LocalMux
    port map (
            O => \N__47758\,
            I => \N__47649\
        );

    \I__11119\ : LocalMux
    port map (
            O => \N__47755\,
            I => \N__47646\
        );

    \I__11118\ : InMux
    port map (
            O => \N__47754\,
            I => \N__47643\
        );

    \I__11117\ : InMux
    port map (
            O => \N__47753\,
            I => \N__47640\
        );

    \I__11116\ : InMux
    port map (
            O => \N__47752\,
            I => \N__47637\
        );

    \I__11115\ : LocalMux
    port map (
            O => \N__47749\,
            I => \N__47634\
        );

    \I__11114\ : InMux
    port map (
            O => \N__47748\,
            I => \N__47631\
        );

    \I__11113\ : InMux
    port map (
            O => \N__47747\,
            I => \N__47628\
        );

    \I__11112\ : InMux
    port map (
            O => \N__47746\,
            I => \N__47623\
        );

    \I__11111\ : InMux
    port map (
            O => \N__47745\,
            I => \N__47623\
        );

    \I__11110\ : InMux
    port map (
            O => \N__47744\,
            I => \N__47618\
        );

    \I__11109\ : InMux
    port map (
            O => \N__47743\,
            I => \N__47618\
        );

    \I__11108\ : InMux
    port map (
            O => \N__47742\,
            I => \N__47615\
        );

    \I__11107\ : InMux
    port map (
            O => \N__47741\,
            I => \N__47612\
        );

    \I__11106\ : LocalMux
    port map (
            O => \N__47738\,
            I => \N__47609\
        );

    \I__11105\ : InMux
    port map (
            O => \N__47737\,
            I => \N__47606\
        );

    \I__11104\ : LocalMux
    port map (
            O => \N__47734\,
            I => \N__47601\
        );

    \I__11103\ : LocalMux
    port map (
            O => \N__47731\,
            I => \N__47601\
        );

    \I__11102\ : LocalMux
    port map (
            O => \N__47728\,
            I => \N__47598\
        );

    \I__11101\ : InMux
    port map (
            O => \N__47727\,
            I => \N__47593\
        );

    \I__11100\ : InMux
    port map (
            O => \N__47726\,
            I => \N__47593\
        );

    \I__11099\ : Span4Mux_v
    port map (
            O => \N__47721\,
            I => \N__47584\
        );

    \I__11098\ : Span4Mux_v
    port map (
            O => \N__47718\,
            I => \N__47584\
        );

    \I__11097\ : Span4Mux_v
    port map (
            O => \N__47705\,
            I => \N__47584\
        );

    \I__11096\ : LocalMux
    port map (
            O => \N__47702\,
            I => \N__47584\
        );

    \I__11095\ : CascadeMux
    port map (
            O => \N__47701\,
            I => \N__47581\
        );

    \I__11094\ : InMux
    port map (
            O => \N__47700\,
            I => \N__47573\
        );

    \I__11093\ : InMux
    port map (
            O => \N__47699\,
            I => \N__47573\
        );

    \I__11092\ : InMux
    port map (
            O => \N__47698\,
            I => \N__47568\
        );

    \I__11091\ : InMux
    port map (
            O => \N__47697\,
            I => \N__47568\
        );

    \I__11090\ : InMux
    port map (
            O => \N__47696\,
            I => \N__47565\
        );

    \I__11089\ : InMux
    port map (
            O => \N__47695\,
            I => \N__47562\
        );

    \I__11088\ : InMux
    port map (
            O => \N__47694\,
            I => \N__47559\
        );

    \I__11087\ : LocalMux
    port map (
            O => \N__47691\,
            I => \N__47556\
        );

    \I__11086\ : LocalMux
    port map (
            O => \N__47688\,
            I => \N__47545\
        );

    \I__11085\ : LocalMux
    port map (
            O => \N__47683\,
            I => \N__47545\
        );

    \I__11084\ : LocalMux
    port map (
            O => \N__47674\,
            I => \N__47545\
        );

    \I__11083\ : LocalMux
    port map (
            O => \N__47665\,
            I => \N__47545\
        );

    \I__11082\ : Span4Mux_v
    port map (
            O => \N__47662\,
            I => \N__47545\
        );

    \I__11081\ : LocalMux
    port map (
            O => \N__47659\,
            I => \N__47542\
        );

    \I__11080\ : Span4Mux_v
    port map (
            O => \N__47654\,
            I => \N__47533\
        );

    \I__11079\ : Span4Mux_v
    port map (
            O => \N__47649\,
            I => \N__47533\
        );

    \I__11078\ : Span4Mux_v
    port map (
            O => \N__47646\,
            I => \N__47533\
        );

    \I__11077\ : LocalMux
    port map (
            O => \N__47643\,
            I => \N__47533\
        );

    \I__11076\ : LocalMux
    port map (
            O => \N__47640\,
            I => \N__47520\
        );

    \I__11075\ : LocalMux
    port map (
            O => \N__47637\,
            I => \N__47520\
        );

    \I__11074\ : Span4Mux_v
    port map (
            O => \N__47634\,
            I => \N__47520\
        );

    \I__11073\ : LocalMux
    port map (
            O => \N__47631\,
            I => \N__47520\
        );

    \I__11072\ : LocalMux
    port map (
            O => \N__47628\,
            I => \N__47520\
        );

    \I__11071\ : LocalMux
    port map (
            O => \N__47623\,
            I => \N__47520\
        );

    \I__11070\ : LocalMux
    port map (
            O => \N__47618\,
            I => \N__47509\
        );

    \I__11069\ : LocalMux
    port map (
            O => \N__47615\,
            I => \N__47509\
        );

    \I__11068\ : LocalMux
    port map (
            O => \N__47612\,
            I => \N__47509\
        );

    \I__11067\ : Span4Mux_v
    port map (
            O => \N__47609\,
            I => \N__47509\
        );

    \I__11066\ : LocalMux
    port map (
            O => \N__47606\,
            I => \N__47509\
        );

    \I__11065\ : Span4Mux_v
    port map (
            O => \N__47601\,
            I => \N__47503\
        );

    \I__11064\ : Span4Mux_v
    port map (
            O => \N__47598\,
            I => \N__47503\
        );

    \I__11063\ : LocalMux
    port map (
            O => \N__47593\,
            I => \N__47498\
        );

    \I__11062\ : Span4Mux_h
    port map (
            O => \N__47584\,
            I => \N__47498\
        );

    \I__11061\ : InMux
    port map (
            O => \N__47581\,
            I => \N__47495\
        );

    \I__11060\ : InMux
    port map (
            O => \N__47580\,
            I => \N__47488\
        );

    \I__11059\ : InMux
    port map (
            O => \N__47579\,
            I => \N__47488\
        );

    \I__11058\ : InMux
    port map (
            O => \N__47578\,
            I => \N__47488\
        );

    \I__11057\ : LocalMux
    port map (
            O => \N__47573\,
            I => \N__47479\
        );

    \I__11056\ : LocalMux
    port map (
            O => \N__47568\,
            I => \N__47479\
        );

    \I__11055\ : LocalMux
    port map (
            O => \N__47565\,
            I => \N__47479\
        );

    \I__11054\ : LocalMux
    port map (
            O => \N__47562\,
            I => \N__47479\
        );

    \I__11053\ : LocalMux
    port map (
            O => \N__47559\,
            I => \N__47464\
        );

    \I__11052\ : Span4Mux_v
    port map (
            O => \N__47556\,
            I => \N__47464\
        );

    \I__11051\ : Span4Mux_v
    port map (
            O => \N__47545\,
            I => \N__47464\
        );

    \I__11050\ : Span4Mux_v
    port map (
            O => \N__47542\,
            I => \N__47464\
        );

    \I__11049\ : Span4Mux_h
    port map (
            O => \N__47533\,
            I => \N__47464\
        );

    \I__11048\ : Span4Mux_v
    port map (
            O => \N__47520\,
            I => \N__47464\
        );

    \I__11047\ : Span4Mux_h
    port map (
            O => \N__47509\,
            I => \N__47464\
        );

    \I__11046\ : InMux
    port map (
            O => \N__47508\,
            I => \N__47461\
        );

    \I__11045\ : Span4Mux_h
    port map (
            O => \N__47503\,
            I => \N__47456\
        );

    \I__11044\ : Span4Mux_h
    port map (
            O => \N__47498\,
            I => \N__47456\
        );

    \I__11043\ : LocalMux
    port map (
            O => \N__47495\,
            I => comm_cmd_2
        );

    \I__11042\ : LocalMux
    port map (
            O => \N__47488\,
            I => comm_cmd_2
        );

    \I__11041\ : Odrv12
    port map (
            O => \N__47479\,
            I => comm_cmd_2
        );

    \I__11040\ : Odrv4
    port map (
            O => \N__47464\,
            I => comm_cmd_2
        );

    \I__11039\ : LocalMux
    port map (
            O => \N__47461\,
            I => comm_cmd_2
        );

    \I__11038\ : Odrv4
    port map (
            O => \N__47456\,
            I => comm_cmd_2
        );

    \I__11037\ : InMux
    port map (
            O => \N__47443\,
            I => \N__47440\
        );

    \I__11036\ : LocalMux
    port map (
            O => \N__47440\,
            I => \N__47437\
        );

    \I__11035\ : Span4Mux_h
    port map (
            O => \N__47437\,
            I => \N__47434\
        );

    \I__11034\ : Odrv4
    port map (
            O => \N__47434\,
            I => buf_data_iac_7
        );

    \I__11033\ : CascadeMux
    port map (
            O => \N__47431\,
            I => \n22_adj_1590_cascade_\
        );

    \I__11032\ : InMux
    port map (
            O => \N__47428\,
            I => \N__47425\
        );

    \I__11031\ : LocalMux
    port map (
            O => \N__47425\,
            I => \N__47422\
        );

    \I__11030\ : Span4Mux_v
    port map (
            O => \N__47422\,
            I => \N__47419\
        );

    \I__11029\ : Span4Mux_h
    port map (
            O => \N__47419\,
            I => \N__47416\
        );

    \I__11028\ : Odrv4
    port map (
            O => \N__47416\,
            I => n30_adj_1591
        );

    \I__11027\ : InMux
    port map (
            O => \N__47413\,
            I => \N__47409\
        );

    \I__11026\ : InMux
    port map (
            O => \N__47412\,
            I => \N__47406\
        );

    \I__11025\ : LocalMux
    port map (
            O => \N__47409\,
            I => \N__47403\
        );

    \I__11024\ : LocalMux
    port map (
            O => \N__47406\,
            I => \N__47399\
        );

    \I__11023\ : Span4Mux_h
    port map (
            O => \N__47403\,
            I => \N__47396\
        );

    \I__11022\ : InMux
    port map (
            O => \N__47402\,
            I => \N__47393\
        );

    \I__11021\ : Span4Mux_h
    port map (
            O => \N__47399\,
            I => \N__47390\
        );

    \I__11020\ : Span4Mux_h
    port map (
            O => \N__47396\,
            I => \N__47387\
        );

    \I__11019\ : LocalMux
    port map (
            O => \N__47393\,
            I => data_cntvec_6
        );

    \I__11018\ : Odrv4
    port map (
            O => \N__47390\,
            I => data_cntvec_6
        );

    \I__11017\ : Odrv4
    port map (
            O => \N__47387\,
            I => data_cntvec_6
        );

    \I__11016\ : InMux
    port map (
            O => \N__47380\,
            I => n19301
        );

    \I__11015\ : InMux
    port map (
            O => \N__47377\,
            I => \N__47373\
        );

    \I__11014\ : InMux
    port map (
            O => \N__47376\,
            I => \N__47370\
        );

    \I__11013\ : LocalMux
    port map (
            O => \N__47373\,
            I => \N__47366\
        );

    \I__11012\ : LocalMux
    port map (
            O => \N__47370\,
            I => \N__47363\
        );

    \I__11011\ : InMux
    port map (
            O => \N__47369\,
            I => \N__47360\
        );

    \I__11010\ : Span4Mux_h
    port map (
            O => \N__47366\,
            I => \N__47357\
        );

    \I__11009\ : Span4Mux_v
    port map (
            O => \N__47363\,
            I => \N__47354\
        );

    \I__11008\ : LocalMux
    port map (
            O => \N__47360\,
            I => data_cntvec_7
        );

    \I__11007\ : Odrv4
    port map (
            O => \N__47357\,
            I => data_cntvec_7
        );

    \I__11006\ : Odrv4
    port map (
            O => \N__47354\,
            I => data_cntvec_7
        );

    \I__11005\ : InMux
    port map (
            O => \N__47347\,
            I => n19302
        );

    \I__11004\ : InMux
    port map (
            O => \N__47344\,
            I => \N__47340\
        );

    \I__11003\ : InMux
    port map (
            O => \N__47343\,
            I => \N__47337\
        );

    \I__11002\ : LocalMux
    port map (
            O => \N__47340\,
            I => \N__47333\
        );

    \I__11001\ : LocalMux
    port map (
            O => \N__47337\,
            I => \N__47330\
        );

    \I__11000\ : InMux
    port map (
            O => \N__47336\,
            I => \N__47327\
        );

    \I__10999\ : Span4Mux_h
    port map (
            O => \N__47333\,
            I => \N__47324\
        );

    \I__10998\ : Span4Mux_h
    port map (
            O => \N__47330\,
            I => \N__47321\
        );

    \I__10997\ : LocalMux
    port map (
            O => \N__47327\,
            I => data_cntvec_8
        );

    \I__10996\ : Odrv4
    port map (
            O => \N__47324\,
            I => data_cntvec_8
        );

    \I__10995\ : Odrv4
    port map (
            O => \N__47321\,
            I => data_cntvec_8
        );

    \I__10994\ : InMux
    port map (
            O => \N__47314\,
            I => \bfn_18_13_0_\
        );

    \I__10993\ : InMux
    port map (
            O => \N__47311\,
            I => \N__47308\
        );

    \I__10992\ : LocalMux
    port map (
            O => \N__47308\,
            I => \N__47304\
        );

    \I__10991\ : InMux
    port map (
            O => \N__47307\,
            I => \N__47301\
        );

    \I__10990\ : Span4Mux_v
    port map (
            O => \N__47304\,
            I => \N__47298\
        );

    \I__10989\ : LocalMux
    port map (
            O => \N__47301\,
            I => \N__47292\
        );

    \I__10988\ : Span4Mux_h
    port map (
            O => \N__47298\,
            I => \N__47292\
        );

    \I__10987\ : InMux
    port map (
            O => \N__47297\,
            I => \N__47289\
        );

    \I__10986\ : Span4Mux_h
    port map (
            O => \N__47292\,
            I => \N__47286\
        );

    \I__10985\ : LocalMux
    port map (
            O => \N__47289\,
            I => data_cntvec_9
        );

    \I__10984\ : Odrv4
    port map (
            O => \N__47286\,
            I => data_cntvec_9
        );

    \I__10983\ : InMux
    port map (
            O => \N__47281\,
            I => n19304
        );

    \I__10982\ : CascadeMux
    port map (
            O => \N__47278\,
            I => \N__47275\
        );

    \I__10981\ : InMux
    port map (
            O => \N__47275\,
            I => \N__47271\
        );

    \I__10980\ : InMux
    port map (
            O => \N__47274\,
            I => \N__47268\
        );

    \I__10979\ : LocalMux
    port map (
            O => \N__47271\,
            I => \N__47264\
        );

    \I__10978\ : LocalMux
    port map (
            O => \N__47268\,
            I => \N__47261\
        );

    \I__10977\ : InMux
    port map (
            O => \N__47267\,
            I => \N__47258\
        );

    \I__10976\ : Span4Mux_v
    port map (
            O => \N__47264\,
            I => \N__47255\
        );

    \I__10975\ : Span12Mux_h
    port map (
            O => \N__47261\,
            I => \N__47252\
        );

    \I__10974\ : LocalMux
    port map (
            O => \N__47258\,
            I => data_cntvec_10
        );

    \I__10973\ : Odrv4
    port map (
            O => \N__47255\,
            I => data_cntvec_10
        );

    \I__10972\ : Odrv12
    port map (
            O => \N__47252\,
            I => data_cntvec_10
        );

    \I__10971\ : InMux
    port map (
            O => \N__47245\,
            I => n19305
        );

    \I__10970\ : InMux
    port map (
            O => \N__47242\,
            I => \N__47237\
        );

    \I__10969\ : InMux
    port map (
            O => \N__47241\,
            I => \N__47234\
        );

    \I__10968\ : InMux
    port map (
            O => \N__47240\,
            I => \N__47231\
        );

    \I__10967\ : LocalMux
    port map (
            O => \N__47237\,
            I => data_cntvec_11
        );

    \I__10966\ : LocalMux
    port map (
            O => \N__47234\,
            I => data_cntvec_11
        );

    \I__10965\ : LocalMux
    port map (
            O => \N__47231\,
            I => data_cntvec_11
        );

    \I__10964\ : InMux
    port map (
            O => \N__47224\,
            I => n19306
        );

    \I__10963\ : InMux
    port map (
            O => \N__47221\,
            I => \N__47218\
        );

    \I__10962\ : LocalMux
    port map (
            O => \N__47218\,
            I => \N__47214\
        );

    \I__10961\ : InMux
    port map (
            O => \N__47217\,
            I => \N__47211\
        );

    \I__10960\ : Span4Mux_v
    port map (
            O => \N__47214\,
            I => \N__47208\
        );

    \I__10959\ : LocalMux
    port map (
            O => \N__47211\,
            I => data_cntvec_12
        );

    \I__10958\ : Odrv4
    port map (
            O => \N__47208\,
            I => data_cntvec_12
        );

    \I__10957\ : InMux
    port map (
            O => \N__47203\,
            I => n19307
        );

    \I__10956\ : InMux
    port map (
            O => \N__47200\,
            I => \N__47197\
        );

    \I__10955\ : LocalMux
    port map (
            O => \N__47197\,
            I => \N__47193\
        );

    \I__10954\ : InMux
    port map (
            O => \N__47196\,
            I => \N__47190\
        );

    \I__10953\ : Span4Mux_v
    port map (
            O => \N__47193\,
            I => \N__47187\
        );

    \I__10952\ : LocalMux
    port map (
            O => \N__47190\,
            I => data_cntvec_13
        );

    \I__10951\ : Odrv4
    port map (
            O => \N__47187\,
            I => data_cntvec_13
        );

    \I__10950\ : InMux
    port map (
            O => \N__47182\,
            I => n19308
        );

    \I__10949\ : CascadeMux
    port map (
            O => \N__47179\,
            I => \n4_adj_1569_cascade_\
        );

    \I__10948\ : InMux
    port map (
            O => \N__47176\,
            I => \N__47173\
        );

    \I__10947\ : LocalMux
    port map (
            O => \N__47173\,
            I => \N__47169\
        );

    \I__10946\ : InMux
    port map (
            O => \N__47172\,
            I => \N__47166\
        );

    \I__10945\ : Sp12to4
    port map (
            O => \N__47169\,
            I => \N__47163\
        );

    \I__10944\ : LocalMux
    port map (
            O => \N__47166\,
            I => comm_buf_6_1
        );

    \I__10943\ : Odrv12
    port map (
            O => \N__47163\,
            I => comm_buf_6_1
        );

    \I__10942\ : CascadeMux
    port map (
            O => \N__47158\,
            I => \n20792_cascade_\
        );

    \I__10941\ : InMux
    port map (
            O => \N__47155\,
            I => \N__47152\
        );

    \I__10940\ : LocalMux
    port map (
            O => \N__47152\,
            I => \N__47149\
        );

    \I__10939\ : Span4Mux_v
    port map (
            O => \N__47149\,
            I => \N__47146\
        );

    \I__10938\ : Span4Mux_h
    port map (
            O => \N__47146\,
            I => \N__47143\
        );

    \I__10937\ : Odrv4
    port map (
            O => \N__47143\,
            I => n21994
        );

    \I__10936\ : CEMux
    port map (
            O => \N__47140\,
            I => \N__47137\
        );

    \I__10935\ : LocalMux
    port map (
            O => \N__47137\,
            I => \N__47132\
        );

    \I__10934\ : CEMux
    port map (
            O => \N__47136\,
            I => \N__47129\
        );

    \I__10933\ : CEMux
    port map (
            O => \N__47135\,
            I => \N__47125\
        );

    \I__10932\ : Span4Mux_v
    port map (
            O => \N__47132\,
            I => \N__47119\
        );

    \I__10931\ : LocalMux
    port map (
            O => \N__47129\,
            I => \N__47119\
        );

    \I__10930\ : CEMux
    port map (
            O => \N__47128\,
            I => \N__47116\
        );

    \I__10929\ : LocalMux
    port map (
            O => \N__47125\,
            I => \N__47113\
        );

    \I__10928\ : CEMux
    port map (
            O => \N__47124\,
            I => \N__47110\
        );

    \I__10927\ : Span4Mux_v
    port map (
            O => \N__47119\,
            I => \N__47105\
        );

    \I__10926\ : LocalMux
    port map (
            O => \N__47116\,
            I => \N__47105\
        );

    \I__10925\ : Span4Mux_v
    port map (
            O => \N__47113\,
            I => \N__47101\
        );

    \I__10924\ : LocalMux
    port map (
            O => \N__47110\,
            I => \N__47098\
        );

    \I__10923\ : Span4Mux_v
    port map (
            O => \N__47105\,
            I => \N__47095\
        );

    \I__10922\ : CEMux
    port map (
            O => \N__47104\,
            I => \N__47092\
        );

    \I__10921\ : Span4Mux_h
    port map (
            O => \N__47101\,
            I => \N__47085\
        );

    \I__10920\ : Span4Mux_v
    port map (
            O => \N__47098\,
            I => \N__47085\
        );

    \I__10919\ : Span4Mux_h
    port map (
            O => \N__47095\,
            I => \N__47085\
        );

    \I__10918\ : LocalMux
    port map (
            O => \N__47092\,
            I => \N__47082\
        );

    \I__10917\ : Sp12to4
    port map (
            O => \N__47085\,
            I => \N__47078\
        );

    \I__10916\ : Span4Mux_h
    port map (
            O => \N__47082\,
            I => \N__47075\
        );

    \I__10915\ : InMux
    port map (
            O => \N__47081\,
            I => \N__47072\
        );

    \I__10914\ : Odrv12
    port map (
            O => \N__47078\,
            I => n12322
        );

    \I__10913\ : Odrv4
    port map (
            O => \N__47075\,
            I => n12322
        );

    \I__10912\ : LocalMux
    port map (
            O => \N__47072\,
            I => n12322
        );

    \I__10911\ : SRMux
    port map (
            O => \N__47065\,
            I => \N__47062\
        );

    \I__10910\ : LocalMux
    port map (
            O => \N__47062\,
            I => \N__47058\
        );

    \I__10909\ : SRMux
    port map (
            O => \N__47061\,
            I => \N__47053\
        );

    \I__10908\ : Span4Mux_v
    port map (
            O => \N__47058\,
            I => \N__47049\
        );

    \I__10907\ : SRMux
    port map (
            O => \N__47057\,
            I => \N__47045\
        );

    \I__10906\ : SRMux
    port map (
            O => \N__47056\,
            I => \N__47042\
        );

    \I__10905\ : LocalMux
    port map (
            O => \N__47053\,
            I => \N__47039\
        );

    \I__10904\ : SRMux
    port map (
            O => \N__47052\,
            I => \N__47036\
        );

    \I__10903\ : Span4Mux_h
    port map (
            O => \N__47049\,
            I => \N__47033\
        );

    \I__10902\ : SRMux
    port map (
            O => \N__47048\,
            I => \N__47030\
        );

    \I__10901\ : LocalMux
    port map (
            O => \N__47045\,
            I => \N__47027\
        );

    \I__10900\ : LocalMux
    port map (
            O => \N__47042\,
            I => \N__47024\
        );

    \I__10899\ : Span4Mux_h
    port map (
            O => \N__47039\,
            I => \N__47019\
        );

    \I__10898\ : LocalMux
    port map (
            O => \N__47036\,
            I => \N__47019\
        );

    \I__10897\ : Span4Mux_v
    port map (
            O => \N__47033\,
            I => \N__47014\
        );

    \I__10896\ : LocalMux
    port map (
            O => \N__47030\,
            I => \N__47014\
        );

    \I__10895\ : Span4Mux_v
    port map (
            O => \N__47027\,
            I => \N__47011\
        );

    \I__10894\ : Span4Mux_h
    port map (
            O => \N__47024\,
            I => \N__47006\
        );

    \I__10893\ : Span4Mux_h
    port map (
            O => \N__47019\,
            I => \N__47006\
        );

    \I__10892\ : Span4Mux_h
    port map (
            O => \N__47014\,
            I => \N__47003\
        );

    \I__10891\ : Odrv4
    port map (
            O => \N__47011\,
            I => n14784
        );

    \I__10890\ : Odrv4
    port map (
            O => \N__47006\,
            I => n14784
        );

    \I__10889\ : Odrv4
    port map (
            O => \N__47003\,
            I => n14784
        );

    \I__10888\ : InMux
    port map (
            O => \N__46996\,
            I => \N__46993\
        );

    \I__10887\ : LocalMux
    port map (
            O => \N__46993\,
            I => \N__46990\
        );

    \I__10886\ : Odrv4
    port map (
            O => \N__46990\,
            I => n21069
        );

    \I__10885\ : CascadeMux
    port map (
            O => \N__46987\,
            I => \N__46983\
        );

    \I__10884\ : InMux
    port map (
            O => \N__46986\,
            I => \N__46980\
        );

    \I__10883\ : InMux
    port map (
            O => \N__46983\,
            I => \N__46977\
        );

    \I__10882\ : LocalMux
    port map (
            O => \N__46980\,
            I => \N__46972\
        );

    \I__10881\ : LocalMux
    port map (
            O => \N__46977\,
            I => \N__46969\
        );

    \I__10880\ : InMux
    port map (
            O => \N__46976\,
            I => \N__46963\
        );

    \I__10879\ : InMux
    port map (
            O => \N__46975\,
            I => \N__46963\
        );

    \I__10878\ : Span4Mux_v
    port map (
            O => \N__46972\,
            I => \N__46960\
        );

    \I__10877\ : Span4Mux_h
    port map (
            O => \N__46969\,
            I => \N__46957\
        );

    \I__10876\ : InMux
    port map (
            O => \N__46968\,
            I => \N__46953\
        );

    \I__10875\ : LocalMux
    port map (
            O => \N__46963\,
            I => \N__46946\
        );

    \I__10874\ : Span4Mux_h
    port map (
            O => \N__46960\,
            I => \N__46946\
        );

    \I__10873\ : Span4Mux_h
    port map (
            O => \N__46957\,
            I => \N__46946\
        );

    \I__10872\ : InMux
    port map (
            O => \N__46956\,
            I => \N__46943\
        );

    \I__10871\ : LocalMux
    port map (
            O => \N__46953\,
            I => \iac_raw_buf_N_728\
        );

    \I__10870\ : Odrv4
    port map (
            O => \N__46946\,
            I => \iac_raw_buf_N_728\
        );

    \I__10869\ : LocalMux
    port map (
            O => \N__46943\,
            I => \iac_raw_buf_N_728\
        );

    \I__10868\ : InMux
    port map (
            O => \N__46936\,
            I => \N__46932\
        );

    \I__10867\ : InMux
    port map (
            O => \N__46935\,
            I => \N__46929\
        );

    \I__10866\ : LocalMux
    port map (
            O => \N__46932\,
            I => \N__46923\
        );

    \I__10865\ : LocalMux
    port map (
            O => \N__46929\,
            I => \N__46923\
        );

    \I__10864\ : InMux
    port map (
            O => \N__46928\,
            I => \N__46920\
        );

    \I__10863\ : Span4Mux_h
    port map (
            O => \N__46923\,
            I => \N__46917\
        );

    \I__10862\ : LocalMux
    port map (
            O => \N__46920\,
            I => data_cntvec_0
        );

    \I__10861\ : Odrv4
    port map (
            O => \N__46917\,
            I => data_cntvec_0
        );

    \I__10860\ : InMux
    port map (
            O => \N__46912\,
            I => \N__46909\
        );

    \I__10859\ : LocalMux
    port map (
            O => \N__46909\,
            I => \N__46904\
        );

    \I__10858\ : InMux
    port map (
            O => \N__46908\,
            I => \N__46901\
        );

    \I__10857\ : InMux
    port map (
            O => \N__46907\,
            I => \N__46898\
        );

    \I__10856\ : Span4Mux_h
    port map (
            O => \N__46904\,
            I => \N__46895\
        );

    \I__10855\ : LocalMux
    port map (
            O => \N__46901\,
            I => \N__46892\
        );

    \I__10854\ : LocalMux
    port map (
            O => \N__46898\,
            I => data_cntvec_1
        );

    \I__10853\ : Odrv4
    port map (
            O => \N__46895\,
            I => data_cntvec_1
        );

    \I__10852\ : Odrv12
    port map (
            O => \N__46892\,
            I => data_cntvec_1
        );

    \I__10851\ : InMux
    port map (
            O => \N__46885\,
            I => n19296
        );

    \I__10850\ : InMux
    port map (
            O => \N__46882\,
            I => \N__46878\
        );

    \I__10849\ : InMux
    port map (
            O => \N__46881\,
            I => \N__46875\
        );

    \I__10848\ : LocalMux
    port map (
            O => \N__46878\,
            I => \N__46872\
        );

    \I__10847\ : LocalMux
    port map (
            O => \N__46875\,
            I => \N__46866\
        );

    \I__10846\ : Span4Mux_h
    port map (
            O => \N__46872\,
            I => \N__46866\
        );

    \I__10845\ : InMux
    port map (
            O => \N__46871\,
            I => \N__46863\
        );

    \I__10844\ : Span4Mux_h
    port map (
            O => \N__46866\,
            I => \N__46860\
        );

    \I__10843\ : LocalMux
    port map (
            O => \N__46863\,
            I => data_cntvec_2
        );

    \I__10842\ : Odrv4
    port map (
            O => \N__46860\,
            I => data_cntvec_2
        );

    \I__10841\ : InMux
    port map (
            O => \N__46855\,
            I => n19297
        );

    \I__10840\ : InMux
    port map (
            O => \N__46852\,
            I => \N__46848\
        );

    \I__10839\ : InMux
    port map (
            O => \N__46851\,
            I => \N__46845\
        );

    \I__10838\ : LocalMux
    port map (
            O => \N__46848\,
            I => \N__46842\
        );

    \I__10837\ : LocalMux
    port map (
            O => \N__46845\,
            I => \N__46839\
        );

    \I__10836\ : Span4Mux_v
    port map (
            O => \N__46842\,
            I => \N__46835\
        );

    \I__10835\ : Span4Mux_h
    port map (
            O => \N__46839\,
            I => \N__46832\
        );

    \I__10834\ : InMux
    port map (
            O => \N__46838\,
            I => \N__46829\
        );

    \I__10833\ : Span4Mux_h
    port map (
            O => \N__46835\,
            I => \N__46826\
        );

    \I__10832\ : Span4Mux_h
    port map (
            O => \N__46832\,
            I => \N__46823\
        );

    \I__10831\ : LocalMux
    port map (
            O => \N__46829\,
            I => data_cntvec_3
        );

    \I__10830\ : Odrv4
    port map (
            O => \N__46826\,
            I => data_cntvec_3
        );

    \I__10829\ : Odrv4
    port map (
            O => \N__46823\,
            I => data_cntvec_3
        );

    \I__10828\ : InMux
    port map (
            O => \N__46816\,
            I => n19298
        );

    \I__10827\ : InMux
    port map (
            O => \N__46813\,
            I => \N__46809\
        );

    \I__10826\ : InMux
    port map (
            O => \N__46812\,
            I => \N__46806\
        );

    \I__10825\ : LocalMux
    port map (
            O => \N__46809\,
            I => \N__46803\
        );

    \I__10824\ : LocalMux
    port map (
            O => \N__46806\,
            I => \N__46797\
        );

    \I__10823\ : Span4Mux_h
    port map (
            O => \N__46803\,
            I => \N__46797\
        );

    \I__10822\ : InMux
    port map (
            O => \N__46802\,
            I => \N__46794\
        );

    \I__10821\ : Span4Mux_h
    port map (
            O => \N__46797\,
            I => \N__46791\
        );

    \I__10820\ : LocalMux
    port map (
            O => \N__46794\,
            I => data_cntvec_4
        );

    \I__10819\ : Odrv4
    port map (
            O => \N__46791\,
            I => data_cntvec_4
        );

    \I__10818\ : InMux
    port map (
            O => \N__46786\,
            I => n19299
        );

    \I__10817\ : InMux
    port map (
            O => \N__46783\,
            I => \N__46779\
        );

    \I__10816\ : InMux
    port map (
            O => \N__46782\,
            I => \N__46776\
        );

    \I__10815\ : LocalMux
    port map (
            O => \N__46779\,
            I => \N__46773\
        );

    \I__10814\ : LocalMux
    port map (
            O => \N__46776\,
            I => \N__46767\
        );

    \I__10813\ : Span4Mux_h
    port map (
            O => \N__46773\,
            I => \N__46767\
        );

    \I__10812\ : InMux
    port map (
            O => \N__46772\,
            I => \N__46764\
        );

    \I__10811\ : Span4Mux_h
    port map (
            O => \N__46767\,
            I => \N__46761\
        );

    \I__10810\ : LocalMux
    port map (
            O => \N__46764\,
            I => data_cntvec_5
        );

    \I__10809\ : Odrv4
    port map (
            O => \N__46761\,
            I => data_cntvec_5
        );

    \I__10808\ : InMux
    port map (
            O => \N__46756\,
            I => n19300
        );

    \I__10807\ : InMux
    port map (
            O => \N__46753\,
            I => \N__46750\
        );

    \I__10806\ : LocalMux
    port map (
            O => \N__46750\,
            I => \N__46747\
        );

    \I__10805\ : Span4Mux_h
    port map (
            O => \N__46747\,
            I => \N__46744\
        );

    \I__10804\ : Odrv4
    port map (
            O => \N__46744\,
            I => n4_adj_1566
        );

    \I__10803\ : CascadeMux
    port map (
            O => \N__46741\,
            I => \n22063_cascade_\
        );

    \I__10802\ : InMux
    port map (
            O => \N__46738\,
            I => \N__46735\
        );

    \I__10801\ : LocalMux
    port map (
            O => \N__46735\,
            I => \N__46731\
        );

    \I__10800\ : InMux
    port map (
            O => \N__46734\,
            I => \N__46728\
        );

    \I__10799\ : Span4Mux_h
    port map (
            O => \N__46731\,
            I => \N__46725\
        );

    \I__10798\ : LocalMux
    port map (
            O => \N__46728\,
            I => \N__46720\
        );

    \I__10797\ : Span4Mux_h
    port map (
            O => \N__46725\,
            I => \N__46720\
        );

    \I__10796\ : Odrv4
    port map (
            O => \N__46720\,
            I => comm_buf_6_4
        );

    \I__10795\ : CascadeMux
    port map (
            O => \N__46717\,
            I => \N__46714\
        );

    \I__10794\ : InMux
    port map (
            O => \N__46714\,
            I => \N__46711\
        );

    \I__10793\ : LocalMux
    port map (
            O => \N__46711\,
            I => n21081
        );

    \I__10792\ : CascadeMux
    port map (
            O => \N__46708\,
            I => \N__46704\
        );

    \I__10791\ : InMux
    port map (
            O => \N__46707\,
            I => \N__46701\
        );

    \I__10790\ : InMux
    port map (
            O => \N__46704\,
            I => \N__46697\
        );

    \I__10789\ : LocalMux
    port map (
            O => \N__46701\,
            I => \N__46694\
        );

    \I__10788\ : InMux
    port map (
            O => \N__46700\,
            I => \N__46691\
        );

    \I__10787\ : LocalMux
    port map (
            O => \N__46697\,
            I => \N__46688\
        );

    \I__10786\ : Span4Mux_v
    port map (
            O => \N__46694\,
            I => \N__46683\
        );

    \I__10785\ : LocalMux
    port map (
            O => \N__46691\,
            I => \N__46683\
        );

    \I__10784\ : Span4Mux_v
    port map (
            O => \N__46688\,
            I => \N__46680\
        );

    \I__10783\ : Sp12to4
    port map (
            O => \N__46683\,
            I => \N__46677\
        );

    \I__10782\ : Span4Mux_h
    port map (
            O => \N__46680\,
            I => \N__46674\
        );

    \I__10781\ : Span12Mux_h
    port map (
            O => \N__46677\,
            I => \N__46671\
        );

    \I__10780\ : Odrv4
    port map (
            O => \N__46674\,
            I => comm_buf_0_4
        );

    \I__10779\ : Odrv12
    port map (
            O => \N__46671\,
            I => comm_buf_0_4
        );

    \I__10778\ : InMux
    port map (
            O => \N__46666\,
            I => \N__46661\
        );

    \I__10777\ : CascadeMux
    port map (
            O => \N__46665\,
            I => \N__46658\
        );

    \I__10776\ : InMux
    port map (
            O => \N__46664\,
            I => \N__46655\
        );

    \I__10775\ : LocalMux
    port map (
            O => \N__46661\,
            I => \N__46651\
        );

    \I__10774\ : InMux
    port map (
            O => \N__46658\,
            I => \N__46648\
        );

    \I__10773\ : LocalMux
    port map (
            O => \N__46655\,
            I => \N__46643\
        );

    \I__10772\ : InMux
    port map (
            O => \N__46654\,
            I => \N__46640\
        );

    \I__10771\ : Span4Mux_v
    port map (
            O => \N__46651\,
            I => \N__46637\
        );

    \I__10770\ : LocalMux
    port map (
            O => \N__46648\,
            I => \N__46634\
        );

    \I__10769\ : InMux
    port map (
            O => \N__46647\,
            I => \N__46631\
        );

    \I__10768\ : InMux
    port map (
            O => \N__46646\,
            I => \N__46628\
        );

    \I__10767\ : Span4Mux_v
    port map (
            O => \N__46643\,
            I => \N__46625\
        );

    \I__10766\ : LocalMux
    port map (
            O => \N__46640\,
            I => \N__46622\
        );

    \I__10765\ : Span4Mux_h
    port map (
            O => \N__46637\,
            I => \N__46619\
        );

    \I__10764\ : Span4Mux_h
    port map (
            O => \N__46634\,
            I => \N__46614\
        );

    \I__10763\ : LocalMux
    port map (
            O => \N__46631\,
            I => \N__46614\
        );

    \I__10762\ : LocalMux
    port map (
            O => \N__46628\,
            I => \N__46611\
        );

    \I__10761\ : Span4Mux_h
    port map (
            O => \N__46625\,
            I => \N__46606\
        );

    \I__10760\ : Span4Mux_h
    port map (
            O => \N__46622\,
            I => \N__46606\
        );

    \I__10759\ : Odrv4
    port map (
            O => \N__46619\,
            I => comm_buf_1_4
        );

    \I__10758\ : Odrv4
    port map (
            O => \N__46614\,
            I => comm_buf_1_4
        );

    \I__10757\ : Odrv12
    port map (
            O => \N__46611\,
            I => comm_buf_1_4
        );

    \I__10756\ : Odrv4
    port map (
            O => \N__46606\,
            I => comm_buf_1_4
        );

    \I__10755\ : InMux
    port map (
            O => \N__46597\,
            I => \N__46594\
        );

    \I__10754\ : LocalMux
    port map (
            O => \N__46594\,
            I => n1_adj_1564
        );

    \I__10753\ : CascadeMux
    port map (
            O => \N__46591\,
            I => \n18824_cascade_\
        );

    \I__10752\ : InMux
    port map (
            O => \N__46588\,
            I => \N__46585\
        );

    \I__10751\ : LocalMux
    port map (
            O => \N__46585\,
            I => \N__46582\
        );

    \I__10750\ : Span4Mux_v
    port map (
            O => \N__46582\,
            I => \N__46578\
        );

    \I__10749\ : InMux
    port map (
            O => \N__46581\,
            I => \N__46575\
        );

    \I__10748\ : Span4Mux_h
    port map (
            O => \N__46578\,
            I => \N__46570\
        );

    \I__10747\ : LocalMux
    port map (
            O => \N__46575\,
            I => \N__46570\
        );

    \I__10746\ : Odrv4
    port map (
            O => \N__46570\,
            I => n20507
        );

    \I__10745\ : CascadeMux
    port map (
            O => \N__46567\,
            I => \N__46564\
        );

    \I__10744\ : InMux
    port map (
            O => \N__46564\,
            I => \N__46561\
        );

    \I__10743\ : LocalMux
    port map (
            O => \N__46561\,
            I => \N__46558\
        );

    \I__10742\ : Span4Mux_h
    port map (
            O => \N__46558\,
            I => \N__46555\
        );

    \I__10741\ : Odrv4
    port map (
            O => \N__46555\,
            I => comm_buf_2_4
        );

    \I__10740\ : InMux
    port map (
            O => \N__46552\,
            I => \N__46549\
        );

    \I__10739\ : LocalMux
    port map (
            O => \N__46549\,
            I => \N__46546\
        );

    \I__10738\ : Span4Mux_v
    port map (
            O => \N__46546\,
            I => \N__46543\
        );

    \I__10737\ : Span4Mux_h
    port map (
            O => \N__46543\,
            I => \N__46540\
        );

    \I__10736\ : Odrv4
    port map (
            O => \N__46540\,
            I => comm_buf_3_4
        );

    \I__10735\ : InMux
    port map (
            O => \N__46537\,
            I => \N__46534\
        );

    \I__10734\ : LocalMux
    port map (
            O => \N__46534\,
            I => n2_adj_1565
        );

    \I__10733\ : InMux
    port map (
            O => \N__46531\,
            I => \N__46528\
        );

    \I__10732\ : LocalMux
    port map (
            O => \N__46528\,
            I => \N__46525\
        );

    \I__10731\ : Odrv12
    port map (
            O => \N__46525\,
            I => comm_buf_5_1
        );

    \I__10730\ : InMux
    port map (
            O => \N__46522\,
            I => \N__46519\
        );

    \I__10729\ : LocalMux
    port map (
            O => \N__46519\,
            I => \N__46516\
        );

    \I__10728\ : Span4Mux_h
    port map (
            O => \N__46516\,
            I => \N__46513\
        );

    \I__10727\ : Odrv4
    port map (
            O => \N__46513\,
            I => comm_buf_4_1
        );

    \I__10726\ : CascadeMux
    port map (
            O => \N__46510\,
            I => \n4_adj_1483_cascade_\
        );

    \I__10725\ : InMux
    port map (
            O => \N__46507\,
            I => \N__46504\
        );

    \I__10724\ : LocalMux
    port map (
            O => \N__46504\,
            I => \N__46501\
        );

    \I__10723\ : Span4Mux_h
    port map (
            O => \N__46501\,
            I => \N__46497\
        );

    \I__10722\ : InMux
    port map (
            O => \N__46500\,
            I => \N__46494\
        );

    \I__10721\ : Span4Mux_h
    port map (
            O => \N__46497\,
            I => \N__46491\
        );

    \I__10720\ : LocalMux
    port map (
            O => \N__46494\,
            I => \N__46488\
        );

    \I__10719\ : Odrv4
    port map (
            O => \N__46491\,
            I => n12205
        );

    \I__10718\ : Odrv4
    port map (
            O => \N__46488\,
            I => n12205
        );

    \I__10717\ : InMux
    port map (
            O => \N__46483\,
            I => \N__46480\
        );

    \I__10716\ : LocalMux
    port map (
            O => \N__46480\,
            I => \N__46477\
        );

    \I__10715\ : Span12Mux_v
    port map (
            O => \N__46477\,
            I => \N__46474\
        );

    \I__10714\ : Odrv12
    port map (
            O => \N__46474\,
            I => n4
        );

    \I__10713\ : CascadeMux
    port map (
            O => \N__46471\,
            I => \n20510_cascade_\
        );

    \I__10712\ : InMux
    port map (
            O => \N__46468\,
            I => \N__46462\
        );

    \I__10711\ : InMux
    port map (
            O => \N__46467\,
            I => \N__46462\
        );

    \I__10710\ : LocalMux
    port map (
            O => \N__46462\,
            I => \N__46459\
        );

    \I__10709\ : Span4Mux_v
    port map (
            O => \N__46459\,
            I => \N__46456\
        );

    \I__10708\ : Odrv4
    port map (
            O => \N__46456\,
            I => n3
        );

    \I__10707\ : CEMux
    port map (
            O => \N__46453\,
            I => \N__46450\
        );

    \I__10706\ : LocalMux
    port map (
            O => \N__46450\,
            I => \N__46447\
        );

    \I__10705\ : Span4Mux_h
    port map (
            O => \N__46447\,
            I => \N__46444\
        );

    \I__10704\ : Span4Mux_h
    port map (
            O => \N__46444\,
            I => \N__46441\
        );

    \I__10703\ : Odrv4
    port map (
            O => \N__46441\,
            I => n20534
        );

    \I__10702\ : InMux
    port map (
            O => \N__46438\,
            I => \N__46435\
        );

    \I__10701\ : LocalMux
    port map (
            O => \N__46435\,
            I => n11810
        );

    \I__10700\ : CascadeMux
    port map (
            O => \N__46432\,
            I => \n11810_cascade_\
        );

    \I__10699\ : InMux
    port map (
            O => \N__46429\,
            I => \N__46426\
        );

    \I__10698\ : LocalMux
    port map (
            O => \N__46426\,
            I => \N__46423\
        );

    \I__10697\ : Span4Mux_v
    port map (
            O => \N__46423\,
            I => \N__46419\
        );

    \I__10696\ : InMux
    port map (
            O => \N__46422\,
            I => \N__46416\
        );

    \I__10695\ : Span4Mux_h
    port map (
            O => \N__46419\,
            I => \N__46413\
        );

    \I__10694\ : LocalMux
    port map (
            O => \N__46416\,
            I => n20650
        );

    \I__10693\ : Odrv4
    port map (
            O => \N__46413\,
            I => n20650
        );

    \I__10692\ : CascadeMux
    port map (
            O => \N__46408\,
            I => \n20672_cascade_\
        );

    \I__10691\ : InMux
    port map (
            O => \N__46405\,
            I => \N__46402\
        );

    \I__10690\ : LocalMux
    port map (
            O => \N__46402\,
            I => n20510
        );

    \I__10689\ : InMux
    port map (
            O => \N__46399\,
            I => \N__46395\
        );

    \I__10688\ : InMux
    port map (
            O => \N__46398\,
            I => \N__46392\
        );

    \I__10687\ : LocalMux
    port map (
            O => \N__46395\,
            I => n20585
        );

    \I__10686\ : LocalMux
    port map (
            O => \N__46392\,
            I => n20585
        );

    \I__10685\ : InMux
    port map (
            O => \N__46387\,
            I => \N__46384\
        );

    \I__10684\ : LocalMux
    port map (
            O => \N__46384\,
            I => n11824
        );

    \I__10683\ : InMux
    port map (
            O => \N__46381\,
            I => \N__46378\
        );

    \I__10682\ : LocalMux
    port map (
            O => \N__46378\,
            I => \N__46367\
        );

    \I__10681\ : InMux
    port map (
            O => \N__46377\,
            I => \N__46364\
        );

    \I__10680\ : InMux
    port map (
            O => \N__46376\,
            I => \N__46349\
        );

    \I__10679\ : InMux
    port map (
            O => \N__46375\,
            I => \N__46349\
        );

    \I__10678\ : InMux
    port map (
            O => \N__46374\,
            I => \N__46349\
        );

    \I__10677\ : InMux
    port map (
            O => \N__46373\,
            I => \N__46349\
        );

    \I__10676\ : InMux
    port map (
            O => \N__46372\,
            I => \N__46349\
        );

    \I__10675\ : InMux
    port map (
            O => \N__46371\,
            I => \N__46349\
        );

    \I__10674\ : InMux
    port map (
            O => \N__46370\,
            I => \N__46349\
        );

    \I__10673\ : Odrv12
    port map (
            O => \N__46367\,
            I => \comm_spi.bit_cnt_3\
        );

    \I__10672\ : LocalMux
    port map (
            O => \N__46364\,
            I => \comm_spi.bit_cnt_3\
        );

    \I__10671\ : LocalMux
    port map (
            O => \N__46349\,
            I => \comm_spi.bit_cnt_3\
        );

    \I__10670\ : InMux
    port map (
            O => \N__46342\,
            I => \N__46339\
        );

    \I__10669\ : LocalMux
    port map (
            O => \N__46339\,
            I => \N__46336\
        );

    \I__10668\ : Span4Mux_h
    port map (
            O => \N__46336\,
            I => \N__46333\
        );

    \I__10667\ : Span4Mux_h
    port map (
            O => \N__46333\,
            I => \N__46323\
        );

    \I__10666\ : InMux
    port map (
            O => \N__46332\,
            I => \N__46308\
        );

    \I__10665\ : InMux
    port map (
            O => \N__46331\,
            I => \N__46308\
        );

    \I__10664\ : InMux
    port map (
            O => \N__46330\,
            I => \N__46308\
        );

    \I__10663\ : InMux
    port map (
            O => \N__46329\,
            I => \N__46308\
        );

    \I__10662\ : InMux
    port map (
            O => \N__46328\,
            I => \N__46308\
        );

    \I__10661\ : InMux
    port map (
            O => \N__46327\,
            I => \N__46308\
        );

    \I__10660\ : InMux
    port map (
            O => \N__46326\,
            I => \N__46308\
        );

    \I__10659\ : Odrv4
    port map (
            O => \N__46323\,
            I => \comm_spi.n16858\
        );

    \I__10658\ : LocalMux
    port map (
            O => \N__46308\,
            I => \comm_spi.n16858\
        );

    \I__10657\ : InMux
    port map (
            O => \N__46303\,
            I => \N__46300\
        );

    \I__10656\ : LocalMux
    port map (
            O => \N__46300\,
            I => \N__46297\
        );

    \I__10655\ : Odrv4
    port map (
            O => \N__46297\,
            I => n21087
        );

    \I__10654\ : InMux
    port map (
            O => \N__46294\,
            I => \N__46290\
        );

    \I__10653\ : InMux
    port map (
            O => \N__46293\,
            I => \N__46287\
        );

    \I__10652\ : LocalMux
    port map (
            O => \N__46290\,
            I => \comm_spi.n14620\
        );

    \I__10651\ : LocalMux
    port map (
            O => \N__46287\,
            I => \comm_spi.n14620\
        );

    \I__10650\ : SRMux
    port map (
            O => \N__46282\,
            I => \N__46279\
        );

    \I__10649\ : LocalMux
    port map (
            O => \N__46279\,
            I => \N__46276\
        );

    \I__10648\ : Odrv12
    port map (
            O => \N__46276\,
            I => \comm_spi.data_tx_7__N_772\
        );

    \I__10647\ : InMux
    port map (
            O => \N__46273\,
            I => \N__46270\
        );

    \I__10646\ : LocalMux
    port map (
            O => \N__46270\,
            I => \N__46266\
        );

    \I__10645\ : InMux
    port map (
            O => \N__46269\,
            I => \N__46263\
        );

    \I__10644\ : Span4Mux_v
    port map (
            O => \N__46266\,
            I => \N__46258\
        );

    \I__10643\ : LocalMux
    port map (
            O => \N__46263\,
            I => \N__46258\
        );

    \I__10642\ : Span4Mux_h
    port map (
            O => \N__46258\,
            I => \N__46254\
        );

    \I__10641\ : InMux
    port map (
            O => \N__46257\,
            I => \N__46251\
        );

    \I__10640\ : Odrv4
    port map (
            O => \N__46254\,
            I => \comm_spi.n22638\
        );

    \I__10639\ : LocalMux
    port map (
            O => \N__46251\,
            I => \comm_spi.n22638\
        );

    \I__10638\ : InMux
    port map (
            O => \N__46246\,
            I => \N__46243\
        );

    \I__10637\ : LocalMux
    port map (
            O => \N__46243\,
            I => \N__46239\
        );

    \I__10636\ : InMux
    port map (
            O => \N__46242\,
            I => \N__46236\
        );

    \I__10635\ : Odrv4
    port map (
            O => \N__46239\,
            I => \comm_spi.n14619\
        );

    \I__10634\ : LocalMux
    port map (
            O => \N__46236\,
            I => \comm_spi.n14619\
        );

    \I__10633\ : InMux
    port map (
            O => \N__46231\,
            I => \N__46228\
        );

    \I__10632\ : LocalMux
    port map (
            O => \N__46228\,
            I => \N__46224\
        );

    \I__10631\ : InMux
    port map (
            O => \N__46227\,
            I => \N__46221\
        );

    \I__10630\ : Odrv4
    port map (
            O => \N__46224\,
            I => \comm_spi.n14615\
        );

    \I__10629\ : LocalMux
    port map (
            O => \N__46221\,
            I => \comm_spi.n14615\
        );

    \I__10628\ : SRMux
    port map (
            O => \N__46216\,
            I => \N__46213\
        );

    \I__10627\ : LocalMux
    port map (
            O => \N__46213\,
            I => \N__46210\
        );

    \I__10626\ : Odrv12
    port map (
            O => \N__46210\,
            I => \comm_spi.data_tx_7__N_761\
        );

    \I__10625\ : InMux
    port map (
            O => \N__46207\,
            I => \N__46203\
        );

    \I__10624\ : InMux
    port map (
            O => \N__46206\,
            I => \N__46200\
        );

    \I__10623\ : LocalMux
    port map (
            O => \N__46203\,
            I => \N__46195\
        );

    \I__10622\ : LocalMux
    port map (
            O => \N__46200\,
            I => \N__46195\
        );

    \I__10621\ : Span4Mux_v
    port map (
            O => \N__46195\,
            I => \N__46192\
        );

    \I__10620\ : Sp12to4
    port map (
            O => \N__46192\,
            I => \N__46188\
        );

    \I__10619\ : InMux
    port map (
            O => \N__46191\,
            I => \N__46185\
        );

    \I__10618\ : Odrv12
    port map (
            O => \N__46188\,
            I => \comm_spi.n22641\
        );

    \I__10617\ : LocalMux
    port map (
            O => \N__46185\,
            I => \comm_spi.n22641\
        );

    \I__10616\ : InMux
    port map (
            O => \N__46180\,
            I => \N__46176\
        );

    \I__10615\ : InMux
    port map (
            O => \N__46179\,
            I => \N__46173\
        );

    \I__10614\ : LocalMux
    port map (
            O => \N__46176\,
            I => \N__46168\
        );

    \I__10613\ : LocalMux
    port map (
            O => \N__46173\,
            I => \N__46168\
        );

    \I__10612\ : Span4Mux_v
    port map (
            O => \N__46168\,
            I => \N__46165\
        );

    \I__10611\ : Sp12to4
    port map (
            O => \N__46165\,
            I => \N__46162\
        );

    \I__10610\ : Odrv12
    port map (
            O => \N__46162\,
            I => \comm_spi.n14611\
        );

    \I__10609\ : InMux
    port map (
            O => \N__46159\,
            I => \N__46156\
        );

    \I__10608\ : LocalMux
    port map (
            O => \N__46156\,
            I => \N__46152\
        );

    \I__10607\ : InMux
    port map (
            O => \N__46155\,
            I => \N__46149\
        );

    \I__10606\ : Span4Mux_v
    port map (
            O => \N__46152\,
            I => \N__46146\
        );

    \I__10605\ : LocalMux
    port map (
            O => \N__46149\,
            I => \N__46143\
        );

    \I__10604\ : Odrv4
    port map (
            O => \N__46146\,
            I => \comm_spi.n14612\
        );

    \I__10603\ : Odrv12
    port map (
            O => \N__46143\,
            I => \comm_spi.n14612\
        );

    \I__10602\ : InMux
    port map (
            O => \N__46138\,
            I => \N__46134\
        );

    \I__10601\ : InMux
    port map (
            O => \N__46137\,
            I => \N__46131\
        );

    \I__10600\ : LocalMux
    port map (
            O => \N__46134\,
            I => \N__46128\
        );

    \I__10599\ : LocalMux
    port map (
            O => \N__46131\,
            I => \N__46125\
        );

    \I__10598\ : Odrv4
    port map (
            O => \N__46128\,
            I => \comm_spi.n14616\
        );

    \I__10597\ : Odrv4
    port map (
            O => \N__46125\,
            I => \comm_spi.n14616\
        );

    \I__10596\ : InMux
    port map (
            O => \N__46120\,
            I => \N__46117\
        );

    \I__10595\ : LocalMux
    port map (
            O => \N__46117\,
            I => \N__46114\
        );

    \I__10594\ : Odrv4
    port map (
            O => \N__46114\,
            I => n20641
        );

    \I__10593\ : CascadeMux
    port map (
            O => \N__46111\,
            I => \N__46108\
        );

    \I__10592\ : InMux
    port map (
            O => \N__46108\,
            I => \N__46105\
        );

    \I__10591\ : LocalMux
    port map (
            O => \N__46105\,
            I => \N__46102\
        );

    \I__10590\ : Span4Mux_h
    port map (
            O => \N__46102\,
            I => \N__46099\
        );

    \I__10589\ : Odrv4
    port map (
            O => \N__46099\,
            I => n17656
        );

    \I__10588\ : InMux
    port map (
            O => \N__46096\,
            I => \N__46093\
        );

    \I__10587\ : LocalMux
    port map (
            O => \N__46093\,
            I => \N__46090\
        );

    \I__10586\ : Odrv4
    port map (
            O => \N__46090\,
            I => n21162
        );

    \I__10585\ : CascadeMux
    port map (
            O => \N__46087\,
            I => \n17658_cascade_\
        );

    \I__10584\ : InMux
    port map (
            O => \N__46084\,
            I => \N__46081\
        );

    \I__10583\ : LocalMux
    port map (
            O => \N__46081\,
            I => \N__46078\
        );

    \I__10582\ : Span4Mux_v
    port map (
            O => \N__46078\,
            I => \N__46074\
        );

    \I__10581\ : InMux
    port map (
            O => \N__46077\,
            I => \N__46071\
        );

    \I__10580\ : Sp12to4
    port map (
            O => \N__46074\,
            I => \N__46066\
        );

    \I__10579\ : LocalMux
    port map (
            O => \N__46071\,
            I => \N__46066\
        );

    \I__10578\ : Odrv12
    port map (
            O => \N__46066\,
            I => n20653
        );

    \I__10577\ : CascadeMux
    port map (
            O => \N__46063\,
            I => \n12220_cascade_\
        );

    \I__10576\ : InMux
    port map (
            O => \N__46060\,
            I => \N__46057\
        );

    \I__10575\ : LocalMux
    port map (
            O => \N__46057\,
            I => n17338
        );

    \I__10574\ : InMux
    port map (
            O => \N__46054\,
            I => \N__46050\
        );

    \I__10573\ : InMux
    port map (
            O => \N__46053\,
            I => \N__46047\
        );

    \I__10572\ : LocalMux
    port map (
            O => \N__46050\,
            I => n17336
        );

    \I__10571\ : LocalMux
    port map (
            O => \N__46047\,
            I => n17336
        );

    \I__10570\ : InMux
    port map (
            O => \N__46042\,
            I => \N__46039\
        );

    \I__10569\ : LocalMux
    port map (
            O => \N__46039\,
            I => \N__46034\
        );

    \I__10568\ : InMux
    port map (
            O => \N__46038\,
            I => \N__46031\
        );

    \I__10567\ : InMux
    port map (
            O => \N__46037\,
            I => \N__46028\
        );

    \I__10566\ : Odrv4
    port map (
            O => \N__46034\,
            I => data_index_5
        );

    \I__10565\ : LocalMux
    port map (
            O => \N__46031\,
            I => data_index_5
        );

    \I__10564\ : LocalMux
    port map (
            O => \N__46028\,
            I => data_index_5
        );

    \I__10563\ : InMux
    port map (
            O => \N__46021\,
            I => \N__46010\
        );

    \I__10562\ : InMux
    port map (
            O => \N__46020\,
            I => \N__46007\
        );

    \I__10561\ : InMux
    port map (
            O => \N__46019\,
            I => \N__45994\
        );

    \I__10560\ : InMux
    port map (
            O => \N__46018\,
            I => \N__45994\
        );

    \I__10559\ : InMux
    port map (
            O => \N__46017\,
            I => \N__45994\
        );

    \I__10558\ : InMux
    port map (
            O => \N__46016\,
            I => \N__45994\
        );

    \I__10557\ : InMux
    port map (
            O => \N__46015\,
            I => \N__45994\
        );

    \I__10556\ : InMux
    port map (
            O => \N__46014\,
            I => \N__45991\
        );

    \I__10555\ : InMux
    port map (
            O => \N__46013\,
            I => \N__45988\
        );

    \I__10554\ : LocalMux
    port map (
            O => \N__46010\,
            I => \N__45982\
        );

    \I__10553\ : LocalMux
    port map (
            O => \N__46007\,
            I => \N__45982\
        );

    \I__10552\ : InMux
    port map (
            O => \N__46006\,
            I => \N__45977\
        );

    \I__10551\ : InMux
    port map (
            O => \N__46005\,
            I => \N__45977\
        );

    \I__10550\ : LocalMux
    port map (
            O => \N__45994\,
            I => \N__45974\
        );

    \I__10549\ : LocalMux
    port map (
            O => \N__45991\,
            I => \N__45969\
        );

    \I__10548\ : LocalMux
    port map (
            O => \N__45988\,
            I => \N__45969\
        );

    \I__10547\ : InMux
    port map (
            O => \N__45987\,
            I => \N__45966\
        );

    \I__10546\ : Span4Mux_v
    port map (
            O => \N__45982\,
            I => \N__45960\
        );

    \I__10545\ : LocalMux
    port map (
            O => \N__45977\,
            I => \N__45960\
        );

    \I__10544\ : Span4Mux_h
    port map (
            O => \N__45974\,
            I => \N__45953\
        );

    \I__10543\ : Span4Mux_v
    port map (
            O => \N__45969\,
            I => \N__45953\
        );

    \I__10542\ : LocalMux
    port map (
            O => \N__45966\,
            I => \N__45953\
        );

    \I__10541\ : InMux
    port map (
            O => \N__45965\,
            I => \N__45950\
        );

    \I__10540\ : Sp12to4
    port map (
            O => \N__45960\,
            I => \N__45947\
        );

    \I__10539\ : Span4Mux_h
    port map (
            O => \N__45953\,
            I => \N__45942\
        );

    \I__10538\ : LocalMux
    port map (
            O => \N__45950\,
            I => \N__45942\
        );

    \I__10537\ : Odrv12
    port map (
            O => \N__45947\,
            I => n16708
        );

    \I__10536\ : Odrv4
    port map (
            O => \N__45942\,
            I => n16708
        );

    \I__10535\ : InMux
    port map (
            O => \N__45937\,
            I => \N__45934\
        );

    \I__10534\ : LocalMux
    port map (
            O => \N__45934\,
            I => \N__45930\
        );

    \I__10533\ : InMux
    port map (
            O => \N__45933\,
            I => \N__45927\
        );

    \I__10532\ : Span4Mux_h
    port map (
            O => \N__45930\,
            I => \N__45924\
        );

    \I__10531\ : LocalMux
    port map (
            O => \N__45927\,
            I => \N__45921\
        );

    \I__10530\ : Odrv4
    port map (
            O => \N__45924\,
            I => n20626
        );

    \I__10529\ : Odrv12
    port map (
            O => \N__45921\,
            I => n20626
        );

    \I__10528\ : CascadeMux
    port map (
            O => \N__45916\,
            I => \N__45908\
        );

    \I__10527\ : CascadeMux
    port map (
            O => \N__45915\,
            I => \N__45905\
        );

    \I__10526\ : CascadeMux
    port map (
            O => \N__45914\,
            I => \N__45902\
        );

    \I__10525\ : CascadeMux
    port map (
            O => \N__45913\,
            I => \N__45897\
        );

    \I__10524\ : InMux
    port map (
            O => \N__45912\,
            I => \N__45892\
        );

    \I__10523\ : InMux
    port map (
            O => \N__45911\,
            I => \N__45888\
        );

    \I__10522\ : InMux
    port map (
            O => \N__45908\,
            I => \N__45877\
        );

    \I__10521\ : InMux
    port map (
            O => \N__45905\,
            I => \N__45877\
        );

    \I__10520\ : InMux
    port map (
            O => \N__45902\,
            I => \N__45877\
        );

    \I__10519\ : InMux
    port map (
            O => \N__45901\,
            I => \N__45877\
        );

    \I__10518\ : InMux
    port map (
            O => \N__45900\,
            I => \N__45877\
        );

    \I__10517\ : InMux
    port map (
            O => \N__45897\,
            I => \N__45871\
        );

    \I__10516\ : InMux
    port map (
            O => \N__45896\,
            I => \N__45871\
        );

    \I__10515\ : InMux
    port map (
            O => \N__45895\,
            I => \N__45868\
        );

    \I__10514\ : LocalMux
    port map (
            O => \N__45892\,
            I => \N__45865\
        );

    \I__10513\ : InMux
    port map (
            O => \N__45891\,
            I => \N__45862\
        );

    \I__10512\ : LocalMux
    port map (
            O => \N__45888\,
            I => \N__45859\
        );

    \I__10511\ : LocalMux
    port map (
            O => \N__45877\,
            I => \N__45856\
        );

    \I__10510\ : InMux
    port map (
            O => \N__45876\,
            I => \N__45853\
        );

    \I__10509\ : LocalMux
    port map (
            O => \N__45871\,
            I => \N__45850\
        );

    \I__10508\ : LocalMux
    port map (
            O => \N__45868\,
            I => \N__45847\
        );

    \I__10507\ : Span4Mux_h
    port map (
            O => \N__45865\,
            I => \N__45844\
        );

    \I__10506\ : LocalMux
    port map (
            O => \N__45862\,
            I => \N__45841\
        );

    \I__10505\ : Span4Mux_v
    port map (
            O => \N__45859\,
            I => \N__45835\
        );

    \I__10504\ : Span4Mux_h
    port map (
            O => \N__45856\,
            I => \N__45830\
        );

    \I__10503\ : LocalMux
    port map (
            O => \N__45853\,
            I => \N__45830\
        );

    \I__10502\ : Span4Mux_h
    port map (
            O => \N__45850\,
            I => \N__45822\
        );

    \I__10501\ : Span4Mux_v
    port map (
            O => \N__45847\,
            I => \N__45822\
        );

    \I__10500\ : Span4Mux_v
    port map (
            O => \N__45844\,
            I => \N__45822\
        );

    \I__10499\ : Span4Mux_h
    port map (
            O => \N__45841\,
            I => \N__45819\
        );

    \I__10498\ : InMux
    port map (
            O => \N__45840\,
            I => \N__45816\
        );

    \I__10497\ : InMux
    port map (
            O => \N__45839\,
            I => \N__45811\
        );

    \I__10496\ : InMux
    port map (
            O => \N__45838\,
            I => \N__45811\
        );

    \I__10495\ : Span4Mux_h
    port map (
            O => \N__45835\,
            I => \N__45807\
        );

    \I__10494\ : Span4Mux_h
    port map (
            O => \N__45830\,
            I => \N__45804\
        );

    \I__10493\ : InMux
    port map (
            O => \N__45829\,
            I => \N__45801\
        );

    \I__10492\ : Span4Mux_h
    port map (
            O => \N__45822\,
            I => \N__45798\
        );

    \I__10491\ : Span4Mux_h
    port map (
            O => \N__45819\,
            I => \N__45795\
        );

    \I__10490\ : LocalMux
    port map (
            O => \N__45816\,
            I => \N__45790\
        );

    \I__10489\ : LocalMux
    port map (
            O => \N__45811\,
            I => \N__45790\
        );

    \I__10488\ : InMux
    port map (
            O => \N__45810\,
            I => \N__45787\
        );

    \I__10487\ : Odrv4
    port map (
            O => \N__45807\,
            I => n11805
        );

    \I__10486\ : Odrv4
    port map (
            O => \N__45804\,
            I => n11805
        );

    \I__10485\ : LocalMux
    port map (
            O => \N__45801\,
            I => n11805
        );

    \I__10484\ : Odrv4
    port map (
            O => \N__45798\,
            I => n11805
        );

    \I__10483\ : Odrv4
    port map (
            O => \N__45795\,
            I => n11805
        );

    \I__10482\ : Odrv12
    port map (
            O => \N__45790\,
            I => n11805
        );

    \I__10481\ : LocalMux
    port map (
            O => \N__45787\,
            I => n11805
        );

    \I__10480\ : CascadeMux
    port map (
            O => \N__45772\,
            I => \N__45769\
        );

    \I__10479\ : InMux
    port map (
            O => \N__45769\,
            I => \N__45762\
        );

    \I__10478\ : CascadeMux
    port map (
            O => \N__45768\,
            I => \N__45759\
        );

    \I__10477\ : InMux
    port map (
            O => \N__45767\,
            I => \N__45756\
        );

    \I__10476\ : InMux
    port map (
            O => \N__45766\,
            I => \N__45753\
        );

    \I__10475\ : InMux
    port map (
            O => \N__45765\,
            I => \N__45750\
        );

    \I__10474\ : LocalMux
    port map (
            O => \N__45762\,
            I => \N__45747\
        );

    \I__10473\ : InMux
    port map (
            O => \N__45759\,
            I => \N__45744\
        );

    \I__10472\ : LocalMux
    port map (
            O => \N__45756\,
            I => \N__45741\
        );

    \I__10471\ : LocalMux
    port map (
            O => \N__45753\,
            I => \N__45738\
        );

    \I__10470\ : LocalMux
    port map (
            O => \N__45750\,
            I => \N__45735\
        );

    \I__10469\ : Span4Mux_h
    port map (
            O => \N__45747\,
            I => \N__45728\
        );

    \I__10468\ : LocalMux
    port map (
            O => \N__45744\,
            I => \N__45728\
        );

    \I__10467\ : Span4Mux_v
    port map (
            O => \N__45741\,
            I => \N__45728\
        );

    \I__10466\ : Span4Mux_h
    port map (
            O => \N__45738\,
            I => \N__45724\
        );

    \I__10465\ : Span4Mux_v
    port map (
            O => \N__45735\,
            I => \N__45721\
        );

    \I__10464\ : Span4Mux_h
    port map (
            O => \N__45728\,
            I => \N__45718\
        );

    \I__10463\ : InMux
    port map (
            O => \N__45727\,
            I => \N__45715\
        );

    \I__10462\ : Span4Mux_v
    port map (
            O => \N__45724\,
            I => \N__45712\
        );

    \I__10461\ : Span4Mux_v
    port map (
            O => \N__45721\,
            I => \N__45709\
        );

    \I__10460\ : Span4Mux_h
    port map (
            O => \N__45718\,
            I => \N__45706\
        );

    \I__10459\ : LocalMux
    port map (
            O => \N__45715\,
            I => n14_adj_1523
        );

    \I__10458\ : Odrv4
    port map (
            O => \N__45712\,
            I => n14_adj_1523
        );

    \I__10457\ : Odrv4
    port map (
            O => \N__45709\,
            I => n14_adj_1523
        );

    \I__10456\ : Odrv4
    port map (
            O => \N__45706\,
            I => n14_adj_1523
        );

    \I__10455\ : InMux
    port map (
            O => \N__45697\,
            I => \N__45688\
        );

    \I__10454\ : InMux
    port map (
            O => \N__45696\,
            I => \N__45681\
        );

    \I__10453\ : InMux
    port map (
            O => \N__45695\,
            I => \N__45681\
        );

    \I__10452\ : InMux
    port map (
            O => \N__45694\,
            I => \N__45681\
        );

    \I__10451\ : InMux
    port map (
            O => \N__45693\,
            I => \N__45678\
        );

    \I__10450\ : InMux
    port map (
            O => \N__45692\,
            I => \N__45668\
        );

    \I__10449\ : InMux
    port map (
            O => \N__45691\,
            I => \N__45668\
        );

    \I__10448\ : LocalMux
    port map (
            O => \N__45688\,
            I => \N__45661\
        );

    \I__10447\ : LocalMux
    port map (
            O => \N__45681\,
            I => \N__45661\
        );

    \I__10446\ : LocalMux
    port map (
            O => \N__45678\,
            I => \N__45661\
        );

    \I__10445\ : InMux
    port map (
            O => \N__45677\,
            I => \N__45658\
        );

    \I__10444\ : InMux
    port map (
            O => \N__45676\,
            I => \N__45650\
        );

    \I__10443\ : InMux
    port map (
            O => \N__45675\,
            I => \N__45650\
        );

    \I__10442\ : InMux
    port map (
            O => \N__45674\,
            I => \N__45647\
        );

    \I__10441\ : InMux
    port map (
            O => \N__45673\,
            I => \N__45644\
        );

    \I__10440\ : LocalMux
    port map (
            O => \N__45668\,
            I => \N__45641\
        );

    \I__10439\ : Span4Mux_v
    port map (
            O => \N__45661\,
            I => \N__45638\
        );

    \I__10438\ : LocalMux
    port map (
            O => \N__45658\,
            I => \N__45635\
        );

    \I__10437\ : InMux
    port map (
            O => \N__45657\,
            I => \N__45632\
        );

    \I__10436\ : InMux
    port map (
            O => \N__45656\,
            I => \N__45629\
        );

    \I__10435\ : InMux
    port map (
            O => \N__45655\,
            I => \N__45626\
        );

    \I__10434\ : LocalMux
    port map (
            O => \N__45650\,
            I => \N__45621\
        );

    \I__10433\ : LocalMux
    port map (
            O => \N__45647\,
            I => \N__45621\
        );

    \I__10432\ : LocalMux
    port map (
            O => \N__45644\,
            I => \N__45616\
        );

    \I__10431\ : Span4Mux_v
    port map (
            O => \N__45641\,
            I => \N__45616\
        );

    \I__10430\ : Span4Mux_h
    port map (
            O => \N__45638\,
            I => \N__45611\
        );

    \I__10429\ : Span4Mux_h
    port map (
            O => \N__45635\,
            I => \N__45611\
        );

    \I__10428\ : LocalMux
    port map (
            O => \N__45632\,
            I => \N__45608\
        );

    \I__10427\ : LocalMux
    port map (
            O => \N__45629\,
            I => n12353
        );

    \I__10426\ : LocalMux
    port map (
            O => \N__45626\,
            I => n12353
        );

    \I__10425\ : Odrv12
    port map (
            O => \N__45621\,
            I => n12353
        );

    \I__10424\ : Odrv4
    port map (
            O => \N__45616\,
            I => n12353
        );

    \I__10423\ : Odrv4
    port map (
            O => \N__45611\,
            I => n12353
        );

    \I__10422\ : Odrv4
    port map (
            O => \N__45608\,
            I => n12353
        );

    \I__10421\ : CascadeMux
    port map (
            O => \N__45595\,
            I => \N__45592\
        );

    \I__10420\ : InMux
    port map (
            O => \N__45592\,
            I => \N__45588\
        );

    \I__10419\ : InMux
    port map (
            O => \N__45591\,
            I => \N__45585\
        );

    \I__10418\ : LocalMux
    port map (
            O => \N__45588\,
            I => \N__45582\
        );

    \I__10417\ : LocalMux
    port map (
            O => \N__45585\,
            I => \N__45578\
        );

    \I__10416\ : Span4Mux_v
    port map (
            O => \N__45582\,
            I => \N__45575\
        );

    \I__10415\ : InMux
    port map (
            O => \N__45581\,
            I => \N__45572\
        );

    \I__10414\ : Span4Mux_v
    port map (
            O => \N__45578\,
            I => \N__45567\
        );

    \I__10413\ : Span4Mux_h
    port map (
            O => \N__45575\,
            I => \N__45567\
        );

    \I__10412\ : LocalMux
    port map (
            O => \N__45572\,
            I => buf_dds0_15
        );

    \I__10411\ : Odrv4
    port map (
            O => \N__45567\,
            I => buf_dds0_15
        );

    \I__10410\ : InMux
    port map (
            O => \N__45562\,
            I => \N__45558\
        );

    \I__10409\ : InMux
    port map (
            O => \N__45561\,
            I => \N__45555\
        );

    \I__10408\ : LocalMux
    port map (
            O => \N__45558\,
            I => \N__45552\
        );

    \I__10407\ : LocalMux
    port map (
            O => \N__45555\,
            I => \N__45549\
        );

    \I__10406\ : Span4Mux_v
    port map (
            O => \N__45552\,
            I => \N__45546\
        );

    \I__10405\ : Span4Mux_h
    port map (
            O => \N__45549\,
            I => \N__45543\
        );

    \I__10404\ : Odrv4
    port map (
            O => \N__45546\,
            I => n9
        );

    \I__10403\ : Odrv4
    port map (
            O => \N__45543\,
            I => n9
        );

    \I__10402\ : CEMux
    port map (
            O => \N__45538\,
            I => \N__45535\
        );

    \I__10401\ : LocalMux
    port map (
            O => \N__45535\,
            I => \N__45531\
        );

    \I__10400\ : CEMux
    port map (
            O => \N__45534\,
            I => \N__45528\
        );

    \I__10399\ : Span4Mux_v
    port map (
            O => \N__45531\,
            I => \N__45525\
        );

    \I__10398\ : LocalMux
    port map (
            O => \N__45528\,
            I => \N__45522\
        );

    \I__10397\ : Span4Mux_h
    port map (
            O => \N__45525\,
            I => \N__45519\
        );

    \I__10396\ : Span4Mux_h
    port map (
            O => \N__45522\,
            I => \N__45516\
        );

    \I__10395\ : Odrv4
    port map (
            O => \N__45519\,
            I => \SIG_DDS.n9\
        );

    \I__10394\ : Odrv4
    port map (
            O => \N__45516\,
            I => \SIG_DDS.n9\
        );

    \I__10393\ : IoInMux
    port map (
            O => \N__45511\,
            I => \N__45507\
        );

    \I__10392\ : InMux
    port map (
            O => \N__45510\,
            I => \N__45504\
        );

    \I__10391\ : LocalMux
    port map (
            O => \N__45507\,
            I => \N__45501\
        );

    \I__10390\ : LocalMux
    port map (
            O => \N__45504\,
            I => \N__45498\
        );

    \I__10389\ : Span4Mux_s1_v
    port map (
            O => \N__45501\,
            I => \N__45494\
        );

    \I__10388\ : Span4Mux_h
    port map (
            O => \N__45498\,
            I => \N__45491\
        );

    \I__10387\ : InMux
    port map (
            O => \N__45497\,
            I => \N__45488\
        );

    \I__10386\ : Span4Mux_v
    port map (
            O => \N__45494\,
            I => \N__45483\
        );

    \I__10385\ : Span4Mux_v
    port map (
            O => \N__45491\,
            I => \N__45483\
        );

    \I__10384\ : LocalMux
    port map (
            O => \N__45488\,
            I => \SELIRNG1\
        );

    \I__10383\ : Odrv4
    port map (
            O => \N__45483\,
            I => \SELIRNG1\
        );

    \I__10382\ : InMux
    port map (
            O => \N__45478\,
            I => \N__45474\
        );

    \I__10381\ : CascadeMux
    port map (
            O => \N__45477\,
            I => \N__45471\
        );

    \I__10380\ : LocalMux
    port map (
            O => \N__45474\,
            I => \N__45467\
        );

    \I__10379\ : InMux
    port map (
            O => \N__45471\,
            I => \N__45464\
        );

    \I__10378\ : InMux
    port map (
            O => \N__45470\,
            I => \N__45461\
        );

    \I__10377\ : Span4Mux_h
    port map (
            O => \N__45467\,
            I => \N__45456\
        );

    \I__10376\ : LocalMux
    port map (
            O => \N__45464\,
            I => \N__45456\
        );

    \I__10375\ : LocalMux
    port map (
            O => \N__45461\,
            I => \acadc_skipCount_11\
        );

    \I__10374\ : Odrv4
    port map (
            O => \N__45456\,
            I => \acadc_skipCount_11\
        );

    \I__10373\ : InMux
    port map (
            O => \N__45451\,
            I => \N__45448\
        );

    \I__10372\ : LocalMux
    port map (
            O => \N__45448\,
            I => n23_adj_1518
        );

    \I__10371\ : InMux
    port map (
            O => \N__45445\,
            I => \N__45442\
        );

    \I__10370\ : LocalMux
    port map (
            O => \N__45442\,
            I => comm_length_0
        );

    \I__10369\ : CEMux
    port map (
            O => \N__45439\,
            I => \N__45436\
        );

    \I__10368\ : LocalMux
    port map (
            O => \N__45436\,
            I => \N__45433\
        );

    \I__10367\ : Span4Mux_v
    port map (
            O => \N__45433\,
            I => \N__45428\
        );

    \I__10366\ : InMux
    port map (
            O => \N__45432\,
            I => \N__45425\
        );

    \I__10365\ : InMux
    port map (
            O => \N__45431\,
            I => \N__45422\
        );

    \I__10364\ : Span4Mux_h
    port map (
            O => \N__45428\,
            I => \N__45419\
        );

    \I__10363\ : LocalMux
    port map (
            O => \N__45425\,
            I => \N__45414\
        );

    \I__10362\ : LocalMux
    port map (
            O => \N__45422\,
            I => \N__45414\
        );

    \I__10361\ : Span4Mux_h
    port map (
            O => \N__45419\,
            I => \N__45411\
        );

    \I__10360\ : Span4Mux_h
    port map (
            O => \N__45414\,
            I => \N__45408\
        );

    \I__10359\ : Odrv4
    port map (
            O => \N__45411\,
            I => n11846
        );

    \I__10358\ : Odrv4
    port map (
            O => \N__45408\,
            I => n11846
        );

    \I__10357\ : SRMux
    port map (
            O => \N__45403\,
            I => \N__45400\
        );

    \I__10356\ : LocalMux
    port map (
            O => \N__45400\,
            I => \N__45397\
        );

    \I__10355\ : Odrv12
    port map (
            O => \N__45397\,
            I => n14652
        );

    \I__10354\ : CascadeMux
    port map (
            O => \N__45394\,
            I => \N__45391\
        );

    \I__10353\ : InMux
    port map (
            O => \N__45391\,
            I => \N__45388\
        );

    \I__10352\ : LocalMux
    port map (
            O => \N__45388\,
            I => \N__45385\
        );

    \I__10351\ : Odrv4
    port map (
            O => \N__45385\,
            I => n10553
        );

    \I__10350\ : CascadeMux
    port map (
            O => \N__45382\,
            I => \N__45377\
        );

    \I__10349\ : CascadeMux
    port map (
            O => \N__45381\,
            I => \N__45373\
        );

    \I__10348\ : InMux
    port map (
            O => \N__45380\,
            I => \N__45370\
        );

    \I__10347\ : InMux
    port map (
            O => \N__45377\,
            I => \N__45367\
        );

    \I__10346\ : InMux
    port map (
            O => \N__45376\,
            I => \N__45364\
        );

    \I__10345\ : InMux
    port map (
            O => \N__45373\,
            I => \N__45361\
        );

    \I__10344\ : LocalMux
    port map (
            O => \N__45370\,
            I => \N__45356\
        );

    \I__10343\ : LocalMux
    port map (
            O => \N__45367\,
            I => \N__45356\
        );

    \I__10342\ : LocalMux
    port map (
            O => \N__45364\,
            I => \N__45353\
        );

    \I__10341\ : LocalMux
    port map (
            O => \N__45361\,
            I => \N__45350\
        );

    \I__10340\ : Span4Mux_h
    port map (
            O => \N__45356\,
            I => \N__45347\
        );

    \I__10339\ : Span12Mux_h
    port map (
            O => \N__45353\,
            I => \N__45344\
        );

    \I__10338\ : Span4Mux_h
    port map (
            O => \N__45350\,
            I => \N__45341\
        );

    \I__10337\ : Span4Mux_v
    port map (
            O => \N__45347\,
            I => \N__45338\
        );

    \I__10336\ : Odrv12
    port map (
            O => \N__45344\,
            I => n20622
        );

    \I__10335\ : Odrv4
    port map (
            O => \N__45341\,
            I => n20622
        );

    \I__10334\ : Odrv4
    port map (
            O => \N__45338\,
            I => n20622
        );

    \I__10333\ : InMux
    port map (
            O => \N__45331\,
            I => \N__45324\
        );

    \I__10332\ : InMux
    port map (
            O => \N__45330\,
            I => \N__45317\
        );

    \I__10331\ : InMux
    port map (
            O => \N__45329\,
            I => \N__45317\
        );

    \I__10330\ : InMux
    port map (
            O => \N__45328\,
            I => \N__45317\
        );

    \I__10329\ : InMux
    port map (
            O => \N__45327\,
            I => \N__45314\
        );

    \I__10328\ : LocalMux
    port map (
            O => \N__45324\,
            I => \N__45311\
        );

    \I__10327\ : LocalMux
    port map (
            O => \N__45317\,
            I => \N__45307\
        );

    \I__10326\ : LocalMux
    port map (
            O => \N__45314\,
            I => \N__45304\
        );

    \I__10325\ : Span4Mux_v
    port map (
            O => \N__45311\,
            I => \N__45301\
        );

    \I__10324\ : InMux
    port map (
            O => \N__45310\,
            I => \N__45298\
        );

    \I__10323\ : Span4Mux_h
    port map (
            O => \N__45307\,
            I => \N__45293\
        );

    \I__10322\ : Span4Mux_v
    port map (
            O => \N__45304\,
            I => \N__45293\
        );

    \I__10321\ : Sp12to4
    port map (
            O => \N__45301\,
            I => \N__45289\
        );

    \I__10320\ : LocalMux
    port map (
            O => \N__45298\,
            I => \N__45286\
        );

    \I__10319\ : Span4Mux_h
    port map (
            O => \N__45293\,
            I => \N__45283\
        );

    \I__10318\ : InMux
    port map (
            O => \N__45292\,
            I => \N__45280\
        );

    \I__10317\ : Span12Mux_h
    port map (
            O => \N__45289\,
            I => \N__45276\
        );

    \I__10316\ : Span12Mux_v
    port map (
            O => \N__45286\,
            I => \N__45273\
        );

    \I__10315\ : Span4Mux_h
    port map (
            O => \N__45283\,
            I => \N__45268\
        );

    \I__10314\ : LocalMux
    port map (
            O => \N__45280\,
            I => \N__45268\
        );

    \I__10313\ : InMux
    port map (
            O => \N__45279\,
            I => \N__45265\
        );

    \I__10312\ : Odrv12
    port map (
            O => \N__45276\,
            I => n12381
        );

    \I__10311\ : Odrv12
    port map (
            O => \N__45273\,
            I => n12381
        );

    \I__10310\ : Odrv4
    port map (
            O => \N__45268\,
            I => n12381
        );

    \I__10309\ : LocalMux
    port map (
            O => \N__45265\,
            I => n12381
        );

    \I__10308\ : CascadeMux
    port map (
            O => \N__45256\,
            I => \N__45251\
        );

    \I__10307\ : InMux
    port map (
            O => \N__45255\,
            I => \N__45248\
        );

    \I__10306\ : InMux
    port map (
            O => \N__45254\,
            I => \N__45245\
        );

    \I__10305\ : InMux
    port map (
            O => \N__45251\,
            I => \N__45242\
        );

    \I__10304\ : LocalMux
    port map (
            O => \N__45248\,
            I => req_data_cnt_11
        );

    \I__10303\ : LocalMux
    port map (
            O => \N__45245\,
            I => req_data_cnt_11
        );

    \I__10302\ : LocalMux
    port map (
            O => \N__45242\,
            I => req_data_cnt_11
        );

    \I__10301\ : InMux
    port map (
            O => \N__45235\,
            I => \N__45232\
        );

    \I__10300\ : LocalMux
    port map (
            O => \N__45232\,
            I => \N__45228\
        );

    \I__10299\ : InMux
    port map (
            O => \N__45231\,
            I => \N__45224\
        );

    \I__10298\ : Span12Mux_h
    port map (
            O => \N__45228\,
            I => \N__45221\
        );

    \I__10297\ : InMux
    port map (
            O => \N__45227\,
            I => \N__45218\
        );

    \I__10296\ : LocalMux
    port map (
            O => \N__45224\,
            I => req_data_cnt_14
        );

    \I__10295\ : Odrv12
    port map (
            O => \N__45221\,
            I => req_data_cnt_14
        );

    \I__10294\ : LocalMux
    port map (
            O => \N__45218\,
            I => req_data_cnt_14
        );

    \I__10293\ : InMux
    port map (
            O => \N__45211\,
            I => \N__45208\
        );

    \I__10292\ : LocalMux
    port map (
            O => \N__45208\,
            I => n23_adj_1491
        );

    \I__10291\ : CascadeMux
    port map (
            O => \N__45205\,
            I => \N__45202\
        );

    \I__10290\ : InMux
    port map (
            O => \N__45202\,
            I => \N__45198\
        );

    \I__10289\ : CascadeMux
    port map (
            O => \N__45201\,
            I => \N__45195\
        );

    \I__10288\ : LocalMux
    port map (
            O => \N__45198\,
            I => \N__45192\
        );

    \I__10287\ : InMux
    port map (
            O => \N__45195\,
            I => \N__45189\
        );

    \I__10286\ : Span4Mux_v
    port map (
            O => \N__45192\,
            I => \N__45186\
        );

    \I__10285\ : LocalMux
    port map (
            O => \N__45189\,
            I => \N__45183\
        );

    \I__10284\ : Span4Mux_h
    port map (
            O => \N__45186\,
            I => \N__45180\
        );

    \I__10283\ : Span4Mux_v
    port map (
            O => \N__45183\,
            I => \N__45176\
        );

    \I__10282\ : Span4Mux_h
    port map (
            O => \N__45180\,
            I => \N__45173\
        );

    \I__10281\ : InMux
    port map (
            O => \N__45179\,
            I => \N__45170\
        );

    \I__10280\ : Odrv4
    port map (
            O => \N__45176\,
            I => cmd_rdadctmp_15_adj_1428
        );

    \I__10279\ : Odrv4
    port map (
            O => \N__45173\,
            I => cmd_rdadctmp_15_adj_1428
        );

    \I__10278\ : LocalMux
    port map (
            O => \N__45170\,
            I => cmd_rdadctmp_15_adj_1428
        );

    \I__10277\ : CascadeMux
    port map (
            O => \N__45163\,
            I => \N__45160\
        );

    \I__10276\ : InMux
    port map (
            O => \N__45160\,
            I => \N__45156\
        );

    \I__10275\ : CascadeMux
    port map (
            O => \N__45159\,
            I => \N__45152\
        );

    \I__10274\ : LocalMux
    port map (
            O => \N__45156\,
            I => \N__45149\
        );

    \I__10273\ : InMux
    port map (
            O => \N__45155\,
            I => \N__45144\
        );

    \I__10272\ : InMux
    port map (
            O => \N__45152\,
            I => \N__45144\
        );

    \I__10271\ : Odrv4
    port map (
            O => \N__45149\,
            I => cmd_rdadctmp_15
        );

    \I__10270\ : LocalMux
    port map (
            O => \N__45144\,
            I => cmd_rdadctmp_15
        );

    \I__10269\ : CascadeMux
    port map (
            O => \N__45139\,
            I => \N__45135\
        );

    \I__10268\ : CascadeMux
    port map (
            O => \N__45138\,
            I => \N__45132\
        );

    \I__10267\ : InMux
    port map (
            O => \N__45135\,
            I => \N__45129\
        );

    \I__10266\ : InMux
    port map (
            O => \N__45132\,
            I => \N__45126\
        );

    \I__10265\ : LocalMux
    port map (
            O => \N__45129\,
            I => \N__45123\
        );

    \I__10264\ : LocalMux
    port map (
            O => \N__45126\,
            I => \N__45120\
        );

    \I__10263\ : Span4Mux_h
    port map (
            O => \N__45123\,
            I => \N__45117\
        );

    \I__10262\ : Span4Mux_v
    port map (
            O => \N__45120\,
            I => \N__45114\
        );

    \I__10261\ : Span4Mux_h
    port map (
            O => \N__45117\,
            I => \N__45110\
        );

    \I__10260\ : Sp12to4
    port map (
            O => \N__45114\,
            I => \N__45107\
        );

    \I__10259\ : InMux
    port map (
            O => \N__45113\,
            I => \N__45104\
        );

    \I__10258\ : Span4Mux_h
    port map (
            O => \N__45110\,
            I => \N__45101\
        );

    \I__10257\ : Span12Mux_h
    port map (
            O => \N__45107\,
            I => \N__45098\
        );

    \I__10256\ : LocalMux
    port map (
            O => \N__45104\,
            I => cmd_rdadctmp_16
        );

    \I__10255\ : Odrv4
    port map (
            O => \N__45101\,
            I => cmd_rdadctmp_16
        );

    \I__10254\ : Odrv12
    port map (
            O => \N__45098\,
            I => cmd_rdadctmp_16
        );

    \I__10253\ : CascadeMux
    port map (
            O => \N__45091\,
            I => \N__45088\
        );

    \I__10252\ : InMux
    port map (
            O => \N__45088\,
            I => \N__45083\
        );

    \I__10251\ : InMux
    port map (
            O => \N__45087\,
            I => \N__45080\
        );

    \I__10250\ : InMux
    port map (
            O => \N__45086\,
            I => \N__45077\
        );

    \I__10249\ : LocalMux
    port map (
            O => \N__45083\,
            I => \N__45074\
        );

    \I__10248\ : LocalMux
    port map (
            O => \N__45080\,
            I => req_data_cnt_13
        );

    \I__10247\ : LocalMux
    port map (
            O => \N__45077\,
            I => req_data_cnt_13
        );

    \I__10246\ : Odrv4
    port map (
            O => \N__45074\,
            I => req_data_cnt_13
        );

    \I__10245\ : InMux
    port map (
            O => \N__45067\,
            I => \N__45064\
        );

    \I__10244\ : LocalMux
    port map (
            O => \N__45064\,
            I => \N__45061\
        );

    \I__10243\ : Odrv12
    port map (
            O => \N__45061\,
            I => n21022
        );

    \I__10242\ : CascadeMux
    port map (
            O => \N__45058\,
            I => \N__45055\
        );

    \I__10241\ : InMux
    port map (
            O => \N__45055\,
            I => \N__45052\
        );

    \I__10240\ : LocalMux
    port map (
            O => \N__45052\,
            I => \N__45049\
        );

    \I__10239\ : Span4Mux_v
    port map (
            O => \N__45049\,
            I => \N__45046\
        );

    \I__10238\ : Span4Mux_h
    port map (
            O => \N__45046\,
            I => \N__45043\
        );

    \I__10237\ : Odrv4
    port map (
            O => \N__45043\,
            I => n21049
        );

    \I__10236\ : InMux
    port map (
            O => \N__45040\,
            I => \N__45034\
        );

    \I__10235\ : InMux
    port map (
            O => \N__45039\,
            I => \N__45034\
        );

    \I__10234\ : LocalMux
    port map (
            O => \N__45034\,
            I => comm_length_2
        );

    \I__10233\ : CascadeMux
    port map (
            O => \N__45031\,
            I => \n21955_cascade_\
        );

    \I__10232\ : InMux
    port map (
            O => \N__45028\,
            I => \N__45025\
        );

    \I__10231\ : LocalMux
    port map (
            O => \N__45025\,
            I => n21958
        );

    \I__10230\ : InMux
    port map (
            O => \N__45022\,
            I => \N__45019\
        );

    \I__10229\ : LocalMux
    port map (
            O => \N__45019\,
            I => n21024
        );

    \I__10228\ : InMux
    port map (
            O => \N__45016\,
            I => \N__45013\
        );

    \I__10227\ : LocalMux
    port map (
            O => \N__45013\,
            I => \N__45010\
        );

    \I__10226\ : Span4Mux_v
    port map (
            O => \N__45010\,
            I => \N__45007\
        );

    \I__10225\ : Sp12to4
    port map (
            O => \N__45007\,
            I => \N__45004\
        );

    \I__10224\ : Span12Mux_h
    port map (
            O => \N__45004\,
            I => \N__45001\
        );

    \I__10223\ : Odrv12
    port map (
            O => \N__45001\,
            I => buf_data_iac_19
        );

    \I__10222\ : InMux
    port map (
            O => \N__44998\,
            I => \N__44995\
        );

    \I__10221\ : LocalMux
    port map (
            O => \N__44995\,
            I => n20950
        );

    \I__10220\ : InMux
    port map (
            O => \N__44992\,
            I => \N__44989\
        );

    \I__10219\ : LocalMux
    port map (
            O => \N__44989\,
            I => \N__44985\
        );

    \I__10218\ : InMux
    port map (
            O => \N__44988\,
            I => \N__44982\
        );

    \I__10217\ : Span4Mux_h
    port map (
            O => \N__44985\,
            I => \N__44979\
        );

    \I__10216\ : LocalMux
    port map (
            O => \N__44982\,
            I => data_idxvec_11
        );

    \I__10215\ : Odrv4
    port map (
            O => \N__44979\,
            I => data_idxvec_11
        );

    \I__10214\ : InMux
    port map (
            O => \N__44974\,
            I => \N__44971\
        );

    \I__10213\ : LocalMux
    port map (
            O => \N__44971\,
            I => n26_adj_1519
        );

    \I__10212\ : InMux
    port map (
            O => \N__44968\,
            I => \N__44964\
        );

    \I__10211\ : InMux
    port map (
            O => \N__44967\,
            I => \N__44961\
        );

    \I__10210\ : LocalMux
    port map (
            O => \N__44964\,
            I => secclk_cnt_17
        );

    \I__10209\ : LocalMux
    port map (
            O => \N__44961\,
            I => secclk_cnt_17
        );

    \I__10208\ : InMux
    port map (
            O => \N__44956\,
            I => n19463
        );

    \I__10207\ : InMux
    port map (
            O => \N__44953\,
            I => \N__44949\
        );

    \I__10206\ : InMux
    port map (
            O => \N__44952\,
            I => \N__44946\
        );

    \I__10205\ : LocalMux
    port map (
            O => \N__44949\,
            I => \N__44943\
        );

    \I__10204\ : LocalMux
    port map (
            O => \N__44946\,
            I => secclk_cnt_18
        );

    \I__10203\ : Odrv4
    port map (
            O => \N__44943\,
            I => secclk_cnt_18
        );

    \I__10202\ : InMux
    port map (
            O => \N__44938\,
            I => n19464
        );

    \I__10201\ : InMux
    port map (
            O => \N__44935\,
            I => n19465
        );

    \I__10200\ : InMux
    port map (
            O => \N__44932\,
            I => \N__44928\
        );

    \I__10199\ : InMux
    port map (
            O => \N__44931\,
            I => \N__44925\
        );

    \I__10198\ : LocalMux
    port map (
            O => \N__44928\,
            I => secclk_cnt_20
        );

    \I__10197\ : LocalMux
    port map (
            O => \N__44925\,
            I => secclk_cnt_20
        );

    \I__10196\ : InMux
    port map (
            O => \N__44920\,
            I => n19466
        );

    \I__10195\ : InMux
    port map (
            O => \N__44917\,
            I => n19467
        );

    \I__10194\ : InMux
    port map (
            O => \N__44914\,
            I => n19468
        );

    \I__10193\ : SRMux
    port map (
            O => \N__44911\,
            I => \N__44907\
        );

    \I__10192\ : SRMux
    port map (
            O => \N__44910\,
            I => \N__44903\
        );

    \I__10191\ : LocalMux
    port map (
            O => \N__44907\,
            I => \N__44899\
        );

    \I__10190\ : SRMux
    port map (
            O => \N__44906\,
            I => \N__44896\
        );

    \I__10189\ : LocalMux
    port map (
            O => \N__44903\,
            I => \N__44893\
        );

    \I__10188\ : InMux
    port map (
            O => \N__44902\,
            I => \N__44890\
        );

    \I__10187\ : Span4Mux_v
    port map (
            O => \N__44899\,
            I => \N__44887\
        );

    \I__10186\ : LocalMux
    port map (
            O => \N__44896\,
            I => \N__44884\
        );

    \I__10185\ : Span4Mux_h
    port map (
            O => \N__44893\,
            I => \N__44879\
        );

    \I__10184\ : LocalMux
    port map (
            O => \N__44890\,
            I => \N__44879\
        );

    \I__10183\ : Odrv4
    port map (
            O => \N__44887\,
            I => n14700
        );

    \I__10182\ : Odrv4
    port map (
            O => \N__44884\,
            I => n14700
        );

    \I__10181\ : Odrv4
    port map (
            O => \N__44879\,
            I => n14700
        );

    \I__10180\ : InMux
    port map (
            O => \N__44872\,
            I => \N__44868\
        );

    \I__10179\ : InMux
    port map (
            O => \N__44871\,
            I => \N__44865\
        );

    \I__10178\ : LocalMux
    port map (
            O => \N__44868\,
            I => \N__44862\
        );

    \I__10177\ : LocalMux
    port map (
            O => \N__44865\,
            I => \N__44857\
        );

    \I__10176\ : Span4Mux_h
    port map (
            O => \N__44862\,
            I => \N__44857\
        );

    \I__10175\ : Span4Mux_h
    port map (
            O => \N__44857\,
            I => \N__44854\
        );

    \I__10174\ : Odrv4
    port map (
            O => \N__44854\,
            I => comm_buf_0_5
        );

    \I__10173\ : CascadeMux
    port map (
            O => \N__44851\,
            I => \N__44843\
        );

    \I__10172\ : InMux
    port map (
            O => \N__44850\,
            I => \N__44840\
        );

    \I__10171\ : InMux
    port map (
            O => \N__44849\,
            I => \N__44837\
        );

    \I__10170\ : InMux
    port map (
            O => \N__44848\,
            I => \N__44834\
        );

    \I__10169\ : InMux
    port map (
            O => \N__44847\,
            I => \N__44831\
        );

    \I__10168\ : InMux
    port map (
            O => \N__44846\,
            I => \N__44828\
        );

    \I__10167\ : InMux
    port map (
            O => \N__44843\,
            I => \N__44825\
        );

    \I__10166\ : LocalMux
    port map (
            O => \N__44840\,
            I => \N__44822\
        );

    \I__10165\ : LocalMux
    port map (
            O => \N__44837\,
            I => \N__44819\
        );

    \I__10164\ : LocalMux
    port map (
            O => \N__44834\,
            I => \N__44812\
        );

    \I__10163\ : LocalMux
    port map (
            O => \N__44831\,
            I => \N__44812\
        );

    \I__10162\ : LocalMux
    port map (
            O => \N__44828\,
            I => \N__44812\
        );

    \I__10161\ : LocalMux
    port map (
            O => \N__44825\,
            I => \N__44809\
        );

    \I__10160\ : Span4Mux_h
    port map (
            O => \N__44822\,
            I => \N__44806\
        );

    \I__10159\ : Span4Mux_v
    port map (
            O => \N__44819\,
            I => \N__44801\
        );

    \I__10158\ : Span4Mux_h
    port map (
            O => \N__44812\,
            I => \N__44801\
        );

    \I__10157\ : Span4Mux_v
    port map (
            O => \N__44809\,
            I => \N__44796\
        );

    \I__10156\ : Sp12to4
    port map (
            O => \N__44806\,
            I => \N__44793\
        );

    \I__10155\ : Span4Mux_h
    port map (
            O => \N__44801\,
            I => \N__44790\
        );

    \I__10154\ : InMux
    port map (
            O => \N__44800\,
            I => \N__44785\
        );

    \I__10153\ : InMux
    port map (
            O => \N__44799\,
            I => \N__44785\
        );

    \I__10152\ : Span4Mux_h
    port map (
            O => \N__44796\,
            I => \N__44782\
        );

    \I__10151\ : Span12Mux_v
    port map (
            O => \N__44793\,
            I => \N__44779\
        );

    \I__10150\ : Span4Mux_v
    port map (
            O => \N__44790\,
            I => \N__44776\
        );

    \I__10149\ : LocalMux
    port map (
            O => \N__44785\,
            I => n14_adj_1556
        );

    \I__10148\ : Odrv4
    port map (
            O => \N__44782\,
            I => n14_adj_1556
        );

    \I__10147\ : Odrv12
    port map (
            O => \N__44779\,
            I => n14_adj_1556
        );

    \I__10146\ : Odrv4
    port map (
            O => \N__44776\,
            I => n14_adj_1556
        );

    \I__10145\ : IoInMux
    port map (
            O => \N__44767\,
            I => \N__44764\
        );

    \I__10144\ : LocalMux
    port map (
            O => \N__44764\,
            I => \N__44761\
        );

    \I__10143\ : IoSpan4Mux
    port map (
            O => \N__44761\,
            I => \N__44758\
        );

    \I__10142\ : Span4Mux_s1_h
    port map (
            O => \N__44758\,
            I => \N__44755\
        );

    \I__10141\ : Sp12to4
    port map (
            O => \N__44755\,
            I => \N__44751\
        );

    \I__10140\ : InMux
    port map (
            O => \N__44754\,
            I => \N__44748\
        );

    \I__10139\ : Span12Mux_v
    port map (
            O => \N__44751\,
            I => \N__44745\
        );

    \I__10138\ : LocalMux
    port map (
            O => \N__44748\,
            I => \N__44741\
        );

    \I__10137\ : Span12Mux_h
    port map (
            O => \N__44745\,
            I => \N__44738\
        );

    \I__10136\ : InMux
    port map (
            O => \N__44744\,
            I => \N__44735\
        );

    \I__10135\ : Span4Mux_h
    port map (
            O => \N__44741\,
            I => \N__44732\
        );

    \I__10134\ : Odrv12
    port map (
            O => \N__44738\,
            I => \VDC_RNG0\
        );

    \I__10133\ : LocalMux
    port map (
            O => \N__44735\,
            I => \VDC_RNG0\
        );

    \I__10132\ : Odrv4
    port map (
            O => \N__44732\,
            I => \VDC_RNG0\
        );

    \I__10131\ : InMux
    port map (
            O => \N__44725\,
            I => \N__44722\
        );

    \I__10130\ : LocalMux
    port map (
            O => \N__44722\,
            I => \N__44719\
        );

    \I__10129\ : Span4Mux_h
    port map (
            O => \N__44719\,
            I => \N__44714\
        );

    \I__10128\ : InMux
    port map (
            O => \N__44718\,
            I => \N__44709\
        );

    \I__10127\ : InMux
    port map (
            O => \N__44717\,
            I => \N__44709\
        );

    \I__10126\ : Odrv4
    port map (
            O => \N__44714\,
            I => \acadc_skipCount_12\
        );

    \I__10125\ : LocalMux
    port map (
            O => \N__44709\,
            I => \acadc_skipCount_12\
        );

    \I__10124\ : InMux
    port map (
            O => \N__44704\,
            I => \N__44700\
        );

    \I__10123\ : InMux
    port map (
            O => \N__44703\,
            I => \N__44697\
        );

    \I__10122\ : LocalMux
    port map (
            O => \N__44700\,
            I => secclk_cnt_9
        );

    \I__10121\ : LocalMux
    port map (
            O => \N__44697\,
            I => secclk_cnt_9
        );

    \I__10120\ : InMux
    port map (
            O => \N__44692\,
            I => n19455
        );

    \I__10119\ : CascadeMux
    port map (
            O => \N__44689\,
            I => \N__44685\
        );

    \I__10118\ : InMux
    port map (
            O => \N__44688\,
            I => \N__44682\
        );

    \I__10117\ : InMux
    port map (
            O => \N__44685\,
            I => \N__44679\
        );

    \I__10116\ : LocalMux
    port map (
            O => \N__44682\,
            I => secclk_cnt_10
        );

    \I__10115\ : LocalMux
    port map (
            O => \N__44679\,
            I => secclk_cnt_10
        );

    \I__10114\ : InMux
    port map (
            O => \N__44674\,
            I => n19456
        );

    \I__10113\ : CascadeMux
    port map (
            O => \N__44671\,
            I => \N__44667\
        );

    \I__10112\ : InMux
    port map (
            O => \N__44670\,
            I => \N__44664\
        );

    \I__10111\ : InMux
    port map (
            O => \N__44667\,
            I => \N__44661\
        );

    \I__10110\ : LocalMux
    port map (
            O => \N__44664\,
            I => secclk_cnt_11
        );

    \I__10109\ : LocalMux
    port map (
            O => \N__44661\,
            I => secclk_cnt_11
        );

    \I__10108\ : InMux
    port map (
            O => \N__44656\,
            I => n19457
        );

    \I__10107\ : InMux
    port map (
            O => \N__44653\,
            I => n19458
        );

    \I__10106\ : CascadeMux
    port map (
            O => \N__44650\,
            I => \N__44646\
        );

    \I__10105\ : InMux
    port map (
            O => \N__44649\,
            I => \N__44643\
        );

    \I__10104\ : InMux
    port map (
            O => \N__44646\,
            I => \N__44640\
        );

    \I__10103\ : LocalMux
    port map (
            O => \N__44643\,
            I => secclk_cnt_13
        );

    \I__10102\ : LocalMux
    port map (
            O => \N__44640\,
            I => secclk_cnt_13
        );

    \I__10101\ : InMux
    port map (
            O => \N__44635\,
            I => n19459
        );

    \I__10100\ : InMux
    port map (
            O => \N__44632\,
            I => \N__44628\
        );

    \I__10099\ : InMux
    port map (
            O => \N__44631\,
            I => \N__44625\
        );

    \I__10098\ : LocalMux
    port map (
            O => \N__44628\,
            I => secclk_cnt_14
        );

    \I__10097\ : LocalMux
    port map (
            O => \N__44625\,
            I => secclk_cnt_14
        );

    \I__10096\ : InMux
    port map (
            O => \N__44620\,
            I => n19460
        );

    \I__10095\ : InMux
    port map (
            O => \N__44617\,
            I => \N__44613\
        );

    \I__10094\ : InMux
    port map (
            O => \N__44616\,
            I => \N__44610\
        );

    \I__10093\ : LocalMux
    port map (
            O => \N__44613\,
            I => secclk_cnt_15
        );

    \I__10092\ : LocalMux
    port map (
            O => \N__44610\,
            I => secclk_cnt_15
        );

    \I__10091\ : InMux
    port map (
            O => \N__44605\,
            I => n19461
        );

    \I__10090\ : InMux
    port map (
            O => \N__44602\,
            I => \N__44598\
        );

    \I__10089\ : InMux
    port map (
            O => \N__44601\,
            I => \N__44595\
        );

    \I__10088\ : LocalMux
    port map (
            O => \N__44598\,
            I => secclk_cnt_16
        );

    \I__10087\ : LocalMux
    port map (
            O => \N__44595\,
            I => secclk_cnt_16
        );

    \I__10086\ : InMux
    port map (
            O => \N__44590\,
            I => \bfn_17_11_0_\
        );

    \I__10085\ : InMux
    port map (
            O => \N__44587\,
            I => \N__44583\
        );

    \I__10084\ : InMux
    port map (
            O => \N__44586\,
            I => \N__44580\
        );

    \I__10083\ : LocalMux
    port map (
            O => \N__44583\,
            I => secclk_cnt_0
        );

    \I__10082\ : LocalMux
    port map (
            O => \N__44580\,
            I => secclk_cnt_0
        );

    \I__10081\ : InMux
    port map (
            O => \N__44575\,
            I => \bfn_17_9_0_\
        );

    \I__10080\ : CascadeMux
    port map (
            O => \N__44572\,
            I => \N__44568\
        );

    \I__10079\ : InMux
    port map (
            O => \N__44571\,
            I => \N__44565\
        );

    \I__10078\ : InMux
    port map (
            O => \N__44568\,
            I => \N__44562\
        );

    \I__10077\ : LocalMux
    port map (
            O => \N__44565\,
            I => secclk_cnt_1
        );

    \I__10076\ : LocalMux
    port map (
            O => \N__44562\,
            I => secclk_cnt_1
        );

    \I__10075\ : InMux
    port map (
            O => \N__44557\,
            I => n19447
        );

    \I__10074\ : InMux
    port map (
            O => \N__44554\,
            I => \N__44550\
        );

    \I__10073\ : InMux
    port map (
            O => \N__44553\,
            I => \N__44547\
        );

    \I__10072\ : LocalMux
    port map (
            O => \N__44550\,
            I => secclk_cnt_2
        );

    \I__10071\ : LocalMux
    port map (
            O => \N__44547\,
            I => secclk_cnt_2
        );

    \I__10070\ : InMux
    port map (
            O => \N__44542\,
            I => n19448
        );

    \I__10069\ : InMux
    port map (
            O => \N__44539\,
            I => \N__44536\
        );

    \I__10068\ : LocalMux
    port map (
            O => \N__44536\,
            I => \N__44532\
        );

    \I__10067\ : InMux
    port map (
            O => \N__44535\,
            I => \N__44529\
        );

    \I__10066\ : Odrv4
    port map (
            O => \N__44532\,
            I => secclk_cnt_3
        );

    \I__10065\ : LocalMux
    port map (
            O => \N__44529\,
            I => secclk_cnt_3
        );

    \I__10064\ : InMux
    port map (
            O => \N__44524\,
            I => n19449
        );

    \I__10063\ : InMux
    port map (
            O => \N__44521\,
            I => \N__44517\
        );

    \I__10062\ : InMux
    port map (
            O => \N__44520\,
            I => \N__44514\
        );

    \I__10061\ : LocalMux
    port map (
            O => \N__44517\,
            I => secclk_cnt_4
        );

    \I__10060\ : LocalMux
    port map (
            O => \N__44514\,
            I => secclk_cnt_4
        );

    \I__10059\ : InMux
    port map (
            O => \N__44509\,
            I => n19450
        );

    \I__10058\ : InMux
    port map (
            O => \N__44506\,
            I => \N__44502\
        );

    \I__10057\ : InMux
    port map (
            O => \N__44505\,
            I => \N__44499\
        );

    \I__10056\ : LocalMux
    port map (
            O => \N__44502\,
            I => \N__44496\
        );

    \I__10055\ : LocalMux
    port map (
            O => \N__44499\,
            I => secclk_cnt_5
        );

    \I__10054\ : Odrv4
    port map (
            O => \N__44496\,
            I => secclk_cnt_5
        );

    \I__10053\ : InMux
    port map (
            O => \N__44491\,
            I => n19451
        );

    \I__10052\ : InMux
    port map (
            O => \N__44488\,
            I => \N__44484\
        );

    \I__10051\ : InMux
    port map (
            O => \N__44487\,
            I => \N__44481\
        );

    \I__10050\ : LocalMux
    port map (
            O => \N__44484\,
            I => secclk_cnt_6
        );

    \I__10049\ : LocalMux
    port map (
            O => \N__44481\,
            I => secclk_cnt_6
        );

    \I__10048\ : InMux
    port map (
            O => \N__44476\,
            I => n19452
        );

    \I__10047\ : InMux
    port map (
            O => \N__44473\,
            I => \N__44469\
        );

    \I__10046\ : InMux
    port map (
            O => \N__44472\,
            I => \N__44466\
        );

    \I__10045\ : LocalMux
    port map (
            O => \N__44469\,
            I => \N__44463\
        );

    \I__10044\ : LocalMux
    port map (
            O => \N__44466\,
            I => secclk_cnt_7
        );

    \I__10043\ : Odrv4
    port map (
            O => \N__44463\,
            I => secclk_cnt_7
        );

    \I__10042\ : InMux
    port map (
            O => \N__44458\,
            I => n19453
        );

    \I__10041\ : InMux
    port map (
            O => \N__44455\,
            I => \N__44451\
        );

    \I__10040\ : InMux
    port map (
            O => \N__44454\,
            I => \N__44448\
        );

    \I__10039\ : LocalMux
    port map (
            O => \N__44451\,
            I => secclk_cnt_8
        );

    \I__10038\ : LocalMux
    port map (
            O => \N__44448\,
            I => secclk_cnt_8
        );

    \I__10037\ : InMux
    port map (
            O => \N__44443\,
            I => \bfn_17_10_0_\
        );

    \I__10036\ : InMux
    port map (
            O => \N__44440\,
            I => \N__44437\
        );

    \I__10035\ : LocalMux
    port map (
            O => \N__44437\,
            I => \comm_state_3_N_412_3\
        );

    \I__10034\ : InMux
    port map (
            O => \N__44434\,
            I => \N__44431\
        );

    \I__10033\ : LocalMux
    port map (
            O => \N__44431\,
            I => n1252
        );

    \I__10032\ : InMux
    port map (
            O => \N__44428\,
            I => \N__44425\
        );

    \I__10031\ : LocalMux
    port map (
            O => \N__44425\,
            I => n8_adj_1555
        );

    \I__10030\ : CascadeMux
    port map (
            O => \N__44422\,
            I => \n2342_cascade_\
        );

    \I__10029\ : InMux
    port map (
            O => \N__44419\,
            I => \N__44415\
        );

    \I__10028\ : InMux
    port map (
            O => \N__44418\,
            I => \N__44412\
        );

    \I__10027\ : LocalMux
    port map (
            O => \N__44415\,
            I => \N__44408\
        );

    \I__10026\ : LocalMux
    port map (
            O => \N__44412\,
            I => \N__44405\
        );

    \I__10025\ : InMux
    port map (
            O => \N__44411\,
            I => \N__44402\
        );

    \I__10024\ : Span4Mux_v
    port map (
            O => \N__44408\,
            I => \N__44397\
        );

    \I__10023\ : Span12Mux_v
    port map (
            O => \N__44405\,
            I => \N__44392\
        );

    \I__10022\ : LocalMux
    port map (
            O => \N__44402\,
            I => \N__44392\
        );

    \I__10021\ : InMux
    port map (
            O => \N__44401\,
            I => \N__44389\
        );

    \I__10020\ : InMux
    port map (
            O => \N__44400\,
            I => \N__44386\
        );

    \I__10019\ : Sp12to4
    port map (
            O => \N__44397\,
            I => \N__44379\
        );

    \I__10018\ : Span12Mux_v
    port map (
            O => \N__44392\,
            I => \N__44379\
        );

    \I__10017\ : LocalMux
    port map (
            O => \N__44389\,
            I => \N__44379\
        );

    \I__10016\ : LocalMux
    port map (
            O => \N__44386\,
            I => \comm_state_3_N_428_2\
        );

    \I__10015\ : Odrv12
    port map (
            O => \N__44379\,
            I => \comm_state_3_N_428_2\
        );

    \I__10014\ : CascadeMux
    port map (
            O => \N__44374\,
            I => \n15_adj_1602_cascade_\
        );

    \I__10013\ : InMux
    port map (
            O => \N__44371\,
            I => \N__44368\
        );

    \I__10012\ : LocalMux
    port map (
            O => \N__44368\,
            I => n20571
        );

    \I__10011\ : CascadeMux
    port map (
            O => \N__44365\,
            I => \n20641_cascade_\
        );

    \I__10010\ : InMux
    port map (
            O => \N__44362\,
            I => \N__44359\
        );

    \I__10009\ : LocalMux
    port map (
            O => \N__44359\,
            I => n12_adj_1603
        );

    \I__10008\ : InMux
    port map (
            O => \N__44356\,
            I => \N__44353\
        );

    \I__10007\ : LocalMux
    port map (
            O => \N__44353\,
            I => \N__44350\
        );

    \I__10006\ : Span4Mux_h
    port map (
            O => \N__44350\,
            I => \N__44347\
        );

    \I__10005\ : Span4Mux_h
    port map (
            O => \N__44347\,
            I => \N__44344\
        );

    \I__10004\ : Odrv4
    port map (
            O => \N__44344\,
            I => n7_adj_1588
        );

    \I__10003\ : SRMux
    port map (
            O => \N__44341\,
            I => \N__44338\
        );

    \I__10002\ : LocalMux
    port map (
            O => \N__44338\,
            I => \N__44335\
        );

    \I__10001\ : Span4Mux_v
    port map (
            O => \N__44335\,
            I => \N__44332\
        );

    \I__10000\ : Span4Mux_h
    port map (
            O => \N__44332\,
            I => \N__44329\
        );

    \I__9999\ : Span4Mux_v
    port map (
            O => \N__44329\,
            I => \N__44326\
        );

    \I__9998\ : Odrv4
    port map (
            O => \N__44326\,
            I => \comm_spi.data_tx_7__N_759\
        );

    \I__9997\ : InMux
    port map (
            O => \N__44323\,
            I => \N__44319\
        );

    \I__9996\ : InMux
    port map (
            O => \N__44322\,
            I => \N__44316\
        );

    \I__9995\ : LocalMux
    port map (
            O => \N__44319\,
            I => \comm_spi.n14596\
        );

    \I__9994\ : LocalMux
    port map (
            O => \N__44316\,
            I => \comm_spi.n14596\
        );

    \I__9993\ : InMux
    port map (
            O => \N__44311\,
            I => \N__44307\
        );

    \I__9992\ : InMux
    port map (
            O => \N__44310\,
            I => \N__44304\
        );

    \I__9991\ : LocalMux
    port map (
            O => \N__44307\,
            I => \N__44301\
        );

    \I__9990\ : LocalMux
    port map (
            O => \N__44304\,
            I => \N__44298\
        );

    \I__9989\ : Span4Mux_v
    port map (
            O => \N__44301\,
            I => \N__44295\
        );

    \I__9988\ : Span4Mux_v
    port map (
            O => \N__44298\,
            I => \N__44292\
        );

    \I__9987\ : Odrv4
    port map (
            O => \N__44295\,
            I => \comm_spi.n14595\
        );

    \I__9986\ : Odrv4
    port map (
            O => \N__44292\,
            I => \comm_spi.n14595\
        );

    \I__9985\ : InMux
    port map (
            O => \N__44287\,
            I => \N__44284\
        );

    \I__9984\ : LocalMux
    port map (
            O => \N__44284\,
            I => \N__44279\
        );

    \I__9983\ : InMux
    port map (
            O => \N__44283\,
            I => \N__44276\
        );

    \I__9982\ : InMux
    port map (
            O => \N__44282\,
            I => \N__44273\
        );

    \I__9981\ : Span4Mux_v
    port map (
            O => \N__44279\,
            I => \N__44263\
        );

    \I__9980\ : LocalMux
    port map (
            O => \N__44276\,
            I => \N__44263\
        );

    \I__9979\ : LocalMux
    port map (
            O => \N__44273\,
            I => \N__44263\
        );

    \I__9978\ : InMux
    port map (
            O => \N__44272\,
            I => \N__44260\
        );

    \I__9977\ : InMux
    port map (
            O => \N__44271\,
            I => \N__44257\
        );

    \I__9976\ : InMux
    port map (
            O => \N__44270\,
            I => \N__44254\
        );

    \I__9975\ : Span4Mux_h
    port map (
            O => \N__44263\,
            I => \N__44251\
        );

    \I__9974\ : LocalMux
    port map (
            O => \N__44260\,
            I => \comm_spi.n14588\
        );

    \I__9973\ : LocalMux
    port map (
            O => \N__44257\,
            I => \comm_spi.n14588\
        );

    \I__9972\ : LocalMux
    port map (
            O => \N__44254\,
            I => \comm_spi.n14588\
        );

    \I__9971\ : Odrv4
    port map (
            O => \N__44251\,
            I => \comm_spi.n14588\
        );

    \I__9970\ : InMux
    port map (
            O => \N__44242\,
            I => \N__44239\
        );

    \I__9969\ : LocalMux
    port map (
            O => \N__44239\,
            I => \N__44236\
        );

    \I__9968\ : Odrv4
    port map (
            O => \N__44236\,
            I => \comm_spi.n14590\
        );

    \I__9967\ : SRMux
    port map (
            O => \N__44233\,
            I => \N__44228\
        );

    \I__9966\ : SRMux
    port map (
            O => \N__44232\,
            I => \N__44225\
        );

    \I__9965\ : SRMux
    port map (
            O => \N__44231\,
            I => \N__44222\
        );

    \I__9964\ : LocalMux
    port map (
            O => \N__44228\,
            I => \N__44219\
        );

    \I__9963\ : LocalMux
    port map (
            O => \N__44225\,
            I => \N__44216\
        );

    \I__9962\ : LocalMux
    port map (
            O => \N__44222\,
            I => \N__44213\
        );

    \I__9961\ : Span4Mux_h
    port map (
            O => \N__44219\,
            I => \N__44210\
        );

    \I__9960\ : Span4Mux_v
    port map (
            O => \N__44216\,
            I => \N__44207\
        );

    \I__9959\ : Span4Mux_v
    port map (
            O => \N__44213\,
            I => \N__44204\
        );

    \I__9958\ : Odrv4
    port map (
            O => \N__44210\,
            I => \comm_spi.data_tx_7__N_766\
        );

    \I__9957\ : Odrv4
    port map (
            O => \N__44207\,
            I => \comm_spi.data_tx_7__N_766\
        );

    \I__9956\ : Odrv4
    port map (
            O => \N__44204\,
            I => \comm_spi.data_tx_7__N_766\
        );

    \I__9955\ : InMux
    port map (
            O => \N__44197\,
            I => \N__44194\
        );

    \I__9954\ : LocalMux
    port map (
            O => \N__44194\,
            I => \N__44191\
        );

    \I__9953\ : Span4Mux_h
    port map (
            O => \N__44191\,
            I => \N__44188\
        );

    \I__9952\ : Span4Mux_h
    port map (
            O => \N__44188\,
            I => \N__44185\
        );

    \I__9951\ : Odrv4
    port map (
            O => \N__44185\,
            I => n20931
        );

    \I__9950\ : CascadeMux
    port map (
            O => \N__44182\,
            I => \n21913_cascade_\
        );

    \I__9949\ : InMux
    port map (
            O => \N__44179\,
            I => \N__44176\
        );

    \I__9948\ : LocalMux
    port map (
            O => \N__44176\,
            I => n21916
        );

    \I__9947\ : CascadeMux
    port map (
            O => \N__44173\,
            I => \n1252_cascade_\
        );

    \I__9946\ : InMux
    port map (
            O => \N__44170\,
            I => \N__44167\
        );

    \I__9945\ : LocalMux
    port map (
            O => \N__44167\,
            I => n2
        );

    \I__9944\ : CascadeMux
    port map (
            O => \N__44164\,
            I => \n21088_cascade_\
        );

    \I__9943\ : CEMux
    port map (
            O => \N__44161\,
            I => \N__44158\
        );

    \I__9942\ : LocalMux
    port map (
            O => \N__44158\,
            I => \N__44155\
        );

    \I__9941\ : Span4Mux_v
    port map (
            O => \N__44155\,
            I => \N__44152\
        );

    \I__9940\ : Odrv4
    port map (
            O => \N__44152\,
            I => n14_adj_1497
        );

    \I__9939\ : CascadeMux
    port map (
            O => \N__44149\,
            I => \N__44143\
        );

    \I__9938\ : CascadeMux
    port map (
            O => \N__44148\,
            I => \N__44140\
        );

    \I__9937\ : CascadeMux
    port map (
            O => \N__44147\,
            I => \N__44137\
        );

    \I__9936\ : CascadeMux
    port map (
            O => \N__44146\,
            I => \N__44134\
        );

    \I__9935\ : InMux
    port map (
            O => \N__44143\,
            I => \N__44131\
        );

    \I__9934\ : InMux
    port map (
            O => \N__44140\,
            I => \N__44128\
        );

    \I__9933\ : InMux
    port map (
            O => \N__44137\,
            I => \N__44124\
        );

    \I__9932\ : InMux
    port map (
            O => \N__44134\,
            I => \N__44121\
        );

    \I__9931\ : LocalMux
    port map (
            O => \N__44131\,
            I => \N__44116\
        );

    \I__9930\ : LocalMux
    port map (
            O => \N__44128\,
            I => \N__44116\
        );

    \I__9929\ : InMux
    port map (
            O => \N__44127\,
            I => \N__44113\
        );

    \I__9928\ : LocalMux
    port map (
            O => \N__44124\,
            I => \N__44109\
        );

    \I__9927\ : LocalMux
    port map (
            O => \N__44121\,
            I => \N__44104\
        );

    \I__9926\ : Span4Mux_v
    port map (
            O => \N__44116\,
            I => \N__44101\
        );

    \I__9925\ : LocalMux
    port map (
            O => \N__44113\,
            I => \N__44098\
        );

    \I__9924\ : InMux
    port map (
            O => \N__44112\,
            I => \N__44095\
        );

    \I__9923\ : Span4Mux_v
    port map (
            O => \N__44109\,
            I => \N__44092\
        );

    \I__9922\ : InMux
    port map (
            O => \N__44108\,
            I => \N__44089\
        );

    \I__9921\ : InMux
    port map (
            O => \N__44107\,
            I => \N__44086\
        );

    \I__9920\ : Span4Mux_v
    port map (
            O => \N__44104\,
            I => \N__44081\
        );

    \I__9919\ : Span4Mux_h
    port map (
            O => \N__44101\,
            I => \N__44076\
        );

    \I__9918\ : Span4Mux_v
    port map (
            O => \N__44098\,
            I => \N__44076\
        );

    \I__9917\ : LocalMux
    port map (
            O => \N__44095\,
            I => \N__44073\
        );

    \I__9916\ : Span4Mux_h
    port map (
            O => \N__44092\,
            I => \N__44066\
        );

    \I__9915\ : LocalMux
    port map (
            O => \N__44089\,
            I => \N__44066\
        );

    \I__9914\ : LocalMux
    port map (
            O => \N__44086\,
            I => \N__44066\
        );

    \I__9913\ : InMux
    port map (
            O => \N__44085\,
            I => \N__44061\
        );

    \I__9912\ : InMux
    port map (
            O => \N__44084\,
            I => \N__44061\
        );

    \I__9911\ : Sp12to4
    port map (
            O => \N__44081\,
            I => \N__44058\
        );

    \I__9910\ : Span4Mux_v
    port map (
            O => \N__44076\,
            I => \N__44053\
        );

    \I__9909\ : Span4Mux_v
    port map (
            O => \N__44073\,
            I => \N__44053\
        );

    \I__9908\ : Span4Mux_v
    port map (
            O => \N__44066\,
            I => \N__44050\
        );

    \I__9907\ : LocalMux
    port map (
            O => \N__44061\,
            I => \N__44047\
        );

    \I__9906\ : Span12Mux_v
    port map (
            O => \N__44058\,
            I => \N__44040\
        );

    \I__9905\ : Sp12to4
    port map (
            O => \N__44053\,
            I => \N__44040\
        );

    \I__9904\ : Sp12to4
    port map (
            O => \N__44050\,
            I => \N__44040\
        );

    \I__9903\ : Odrv4
    port map (
            O => \N__44047\,
            I => comm_buf_0_1
        );

    \I__9902\ : Odrv12
    port map (
            O => \N__44040\,
            I => comm_buf_0_1
        );

    \I__9901\ : IoInMux
    port map (
            O => \N__44035\,
            I => \N__44032\
        );

    \I__9900\ : LocalMux
    port map (
            O => \N__44032\,
            I => \N__44028\
        );

    \I__9899\ : InMux
    port map (
            O => \N__44031\,
            I => \N__44025\
        );

    \I__9898\ : IoSpan4Mux
    port map (
            O => \N__44028\,
            I => \N__44022\
        );

    \I__9897\ : LocalMux
    port map (
            O => \N__44025\,
            I => \N__44019\
        );

    \I__9896\ : IoSpan4Mux
    port map (
            O => \N__44022\,
            I => \N__44016\
        );

    \I__9895\ : Span4Mux_h
    port map (
            O => \N__44019\,
            I => \N__44013\
        );

    \I__9894\ : Span4Mux_s3_v
    port map (
            O => \N__44016\,
            I => \N__44010\
        );

    \I__9893\ : Span4Mux_v
    port map (
            O => \N__44013\,
            I => \N__44006\
        );

    \I__9892\ : Span4Mux_v
    port map (
            O => \N__44010\,
            I => \N__44003\
        );

    \I__9891\ : InMux
    port map (
            O => \N__44009\,
            I => \N__44000\
        );

    \I__9890\ : Span4Mux_h
    port map (
            O => \N__44006\,
            I => \N__43997\
        );

    \I__9889\ : Odrv4
    port map (
            O => \N__44003\,
            I => \DDS_RNG_0\
        );

    \I__9888\ : LocalMux
    port map (
            O => \N__44000\,
            I => \DDS_RNG_0\
        );

    \I__9887\ : Odrv4
    port map (
            O => \N__43997\,
            I => \DDS_RNG_0\
        );

    \I__9886\ : InMux
    port map (
            O => \N__43990\,
            I => \N__43987\
        );

    \I__9885\ : LocalMux
    port map (
            O => \N__43987\,
            I => \N__43984\
        );

    \I__9884\ : Odrv4
    port map (
            O => \N__43984\,
            I => n8_adj_1538
        );

    \I__9883\ : InMux
    port map (
            O => \N__43981\,
            I => \N__43977\
        );

    \I__9882\ : InMux
    port map (
            O => \N__43980\,
            I => \N__43974\
        );

    \I__9881\ : LocalMux
    port map (
            O => \N__43977\,
            I => \N__43969\
        );

    \I__9880\ : LocalMux
    port map (
            O => \N__43974\,
            I => \N__43969\
        );

    \I__9879\ : Odrv12
    port map (
            O => \N__43969\,
            I => n7_adj_1537
        );

    \I__9878\ : CascadeMux
    port map (
            O => \N__43966\,
            I => \N__43963\
        );

    \I__9877\ : CascadeBuf
    port map (
            O => \N__43963\,
            I => \N__43960\
        );

    \I__9876\ : CascadeMux
    port map (
            O => \N__43960\,
            I => \N__43957\
        );

    \I__9875\ : CascadeBuf
    port map (
            O => \N__43957\,
            I => \N__43954\
        );

    \I__9874\ : CascadeMux
    port map (
            O => \N__43954\,
            I => \N__43951\
        );

    \I__9873\ : CascadeBuf
    port map (
            O => \N__43951\,
            I => \N__43948\
        );

    \I__9872\ : CascadeMux
    port map (
            O => \N__43948\,
            I => \N__43945\
        );

    \I__9871\ : CascadeBuf
    port map (
            O => \N__43945\,
            I => \N__43942\
        );

    \I__9870\ : CascadeMux
    port map (
            O => \N__43942\,
            I => \N__43939\
        );

    \I__9869\ : CascadeBuf
    port map (
            O => \N__43939\,
            I => \N__43936\
        );

    \I__9868\ : CascadeMux
    port map (
            O => \N__43936\,
            I => \N__43933\
        );

    \I__9867\ : CascadeBuf
    port map (
            O => \N__43933\,
            I => \N__43930\
        );

    \I__9866\ : CascadeMux
    port map (
            O => \N__43930\,
            I => \N__43927\
        );

    \I__9865\ : CascadeBuf
    port map (
            O => \N__43927\,
            I => \N__43924\
        );

    \I__9864\ : CascadeMux
    port map (
            O => \N__43924\,
            I => \N__43920\
        );

    \I__9863\ : CascadeMux
    port map (
            O => \N__43923\,
            I => \N__43917\
        );

    \I__9862\ : CascadeBuf
    port map (
            O => \N__43920\,
            I => \N__43914\
        );

    \I__9861\ : CascadeBuf
    port map (
            O => \N__43917\,
            I => \N__43911\
        );

    \I__9860\ : CascadeMux
    port map (
            O => \N__43914\,
            I => \N__43908\
        );

    \I__9859\ : CascadeMux
    port map (
            O => \N__43911\,
            I => \N__43905\
        );

    \I__9858\ : CascadeBuf
    port map (
            O => \N__43908\,
            I => \N__43902\
        );

    \I__9857\ : InMux
    port map (
            O => \N__43905\,
            I => \N__43899\
        );

    \I__9856\ : CascadeMux
    port map (
            O => \N__43902\,
            I => \N__43896\
        );

    \I__9855\ : LocalMux
    port map (
            O => \N__43899\,
            I => \N__43893\
        );

    \I__9854\ : InMux
    port map (
            O => \N__43896\,
            I => \N__43890\
        );

    \I__9853\ : Span4Mux_v
    port map (
            O => \N__43893\,
            I => \N__43887\
        );

    \I__9852\ : LocalMux
    port map (
            O => \N__43890\,
            I => \N__43884\
        );

    \I__9851\ : Span4Mux_h
    port map (
            O => \N__43887\,
            I => \N__43881\
        );

    \I__9850\ : Span12Mux_h
    port map (
            O => \N__43884\,
            I => \N__43878\
        );

    \I__9849\ : Odrv4
    port map (
            O => \N__43881\,
            I => \data_index_9_N_212_6\
        );

    \I__9848\ : Odrv12
    port map (
            O => \N__43878\,
            I => \data_index_9_N_212_6\
        );

    \I__9847\ : InMux
    port map (
            O => \N__43873\,
            I => \N__43866\
        );

    \I__9846\ : InMux
    port map (
            O => \N__43872\,
            I => \N__43866\
        );

    \I__9845\ : InMux
    port map (
            O => \N__43871\,
            I => \N__43861\
        );

    \I__9844\ : LocalMux
    port map (
            O => \N__43866\,
            I => \N__43858\
        );

    \I__9843\ : InMux
    port map (
            O => \N__43865\,
            I => \N__43855\
        );

    \I__9842\ : InMux
    port map (
            O => \N__43864\,
            I => \N__43852\
        );

    \I__9841\ : LocalMux
    port map (
            O => \N__43861\,
            I => \N__43849\
        );

    \I__9840\ : Span4Mux_v
    port map (
            O => \N__43858\,
            I => \N__43842\
        );

    \I__9839\ : LocalMux
    port map (
            O => \N__43855\,
            I => \N__43842\
        );

    \I__9838\ : LocalMux
    port map (
            O => \N__43852\,
            I => \N__43837\
        );

    \I__9837\ : Span4Mux_h
    port map (
            O => \N__43849\,
            I => \N__43837\
        );

    \I__9836\ : InMux
    port map (
            O => \N__43848\,
            I => \N__43834\
        );

    \I__9835\ : InMux
    port map (
            O => \N__43847\,
            I => \N__43831\
        );

    \I__9834\ : Odrv4
    port map (
            O => \N__43842\,
            I => n11901
        );

    \I__9833\ : Odrv4
    port map (
            O => \N__43837\,
            I => n11901
        );

    \I__9832\ : LocalMux
    port map (
            O => \N__43834\,
            I => n11901
        );

    \I__9831\ : LocalMux
    port map (
            O => \N__43831\,
            I => n11901
        );

    \I__9830\ : CascadeMux
    port map (
            O => \N__43822\,
            I => \N__43818\
        );

    \I__9829\ : InMux
    port map (
            O => \N__43821\,
            I => \N__43813\
        );

    \I__9828\ : InMux
    port map (
            O => \N__43818\,
            I => \N__43810\
        );

    \I__9827\ : InMux
    port map (
            O => \N__43817\,
            I => \N__43807\
        );

    \I__9826\ : CascadeMux
    port map (
            O => \N__43816\,
            I => \N__43803\
        );

    \I__9825\ : LocalMux
    port map (
            O => \N__43813\,
            I => \N__43797\
        );

    \I__9824\ : LocalMux
    port map (
            O => \N__43810\,
            I => \N__43797\
        );

    \I__9823\ : LocalMux
    port map (
            O => \N__43807\,
            I => \N__43793\
        );

    \I__9822\ : CascadeMux
    port map (
            O => \N__43806\,
            I => \N__43790\
        );

    \I__9821\ : InMux
    port map (
            O => \N__43803\,
            I => \N__43787\
        );

    \I__9820\ : InMux
    port map (
            O => \N__43802\,
            I => \N__43784\
        );

    \I__9819\ : Span4Mux_v
    port map (
            O => \N__43797\,
            I => \N__43781\
        );

    \I__9818\ : InMux
    port map (
            O => \N__43796\,
            I => \N__43778\
        );

    \I__9817\ : Span4Mux_h
    port map (
            O => \N__43793\,
            I => \N__43775\
        );

    \I__9816\ : InMux
    port map (
            O => \N__43790\,
            I => \N__43772\
        );

    \I__9815\ : LocalMux
    port map (
            O => \N__43787\,
            I => \N__43769\
        );

    \I__9814\ : LocalMux
    port map (
            O => \N__43784\,
            I => \N__43761\
        );

    \I__9813\ : Span4Mux_v
    port map (
            O => \N__43781\,
            I => \N__43761\
        );

    \I__9812\ : LocalMux
    port map (
            O => \N__43778\,
            I => \N__43761\
        );

    \I__9811\ : Span4Mux_v
    port map (
            O => \N__43775\,
            I => \N__43755\
        );

    \I__9810\ : LocalMux
    port map (
            O => \N__43772\,
            I => \N__43755\
        );

    \I__9809\ : Span4Mux_h
    port map (
            O => \N__43769\,
            I => \N__43752\
        );

    \I__9808\ : InMux
    port map (
            O => \N__43768\,
            I => \N__43749\
        );

    \I__9807\ : Span4Mux_h
    port map (
            O => \N__43761\,
            I => \N__43746\
        );

    \I__9806\ : CascadeMux
    port map (
            O => \N__43760\,
            I => \N__43743\
        );

    \I__9805\ : Span4Mux_h
    port map (
            O => \N__43755\,
            I => \N__43740\
        );

    \I__9804\ : Span4Mux_v
    port map (
            O => \N__43752\,
            I => \N__43735\
        );

    \I__9803\ : LocalMux
    port map (
            O => \N__43749\,
            I => \N__43735\
        );

    \I__9802\ : Span4Mux_h
    port map (
            O => \N__43746\,
            I => \N__43732\
        );

    \I__9801\ : InMux
    port map (
            O => \N__43743\,
            I => \N__43729\
        );

    \I__9800\ : Span4Mux_h
    port map (
            O => \N__43740\,
            I => \N__43726\
        );

    \I__9799\ : Span4Mux_h
    port map (
            O => \N__43735\,
            I => \N__43723\
        );

    \I__9798\ : Sp12to4
    port map (
            O => \N__43732\,
            I => \N__43720\
        );

    \I__9797\ : LocalMux
    port map (
            O => \N__43729\,
            I => comm_buf_0_3
        );

    \I__9796\ : Odrv4
    port map (
            O => \N__43726\,
            I => comm_buf_0_3
        );

    \I__9795\ : Odrv4
    port map (
            O => \N__43723\,
            I => comm_buf_0_3
        );

    \I__9794\ : Odrv12
    port map (
            O => \N__43720\,
            I => comm_buf_0_3
        );

    \I__9793\ : SRMux
    port map (
            O => \N__43711\,
            I => \N__43707\
        );

    \I__9792\ : InMux
    port map (
            O => \N__43710\,
            I => \N__43704\
        );

    \I__9791\ : LocalMux
    port map (
            O => \N__43707\,
            I => \N__43701\
        );

    \I__9790\ : LocalMux
    port map (
            O => \N__43704\,
            I => \N__43698\
        );

    \I__9789\ : Span4Mux_h
    port map (
            O => \N__43701\,
            I => \N__43695\
        );

    \I__9788\ : Span4Mux_v
    port map (
            O => \N__43698\,
            I => \N__43692\
        );

    \I__9787\ : Odrv4
    port map (
            O => \N__43695\,
            I => n14869
        );

    \I__9786\ : Odrv4
    port map (
            O => \N__43692\,
            I => n14869
        );

    \I__9785\ : InMux
    port map (
            O => \N__43687\,
            I => \N__43678\
        );

    \I__9784\ : InMux
    port map (
            O => \N__43686\,
            I => \N__43678\
        );

    \I__9783\ : InMux
    port map (
            O => \N__43685\,
            I => \N__43678\
        );

    \I__9782\ : LocalMux
    port map (
            O => \N__43678\,
            I => \N__43674\
        );

    \I__9781\ : InMux
    port map (
            O => \N__43677\,
            I => \N__43670\
        );

    \I__9780\ : Span4Mux_h
    port map (
            O => \N__43674\,
            I => \N__43667\
        );

    \I__9779\ : CascadeMux
    port map (
            O => \N__43673\,
            I => \N__43664\
        );

    \I__9778\ : LocalMux
    port map (
            O => \N__43670\,
            I => \N__43661\
        );

    \I__9777\ : Span4Mux_v
    port map (
            O => \N__43667\,
            I => \N__43658\
        );

    \I__9776\ : InMux
    port map (
            O => \N__43664\,
            I => \N__43655\
        );

    \I__9775\ : Span12Mux_h
    port map (
            O => \N__43661\,
            I => \N__43652\
        );

    \I__9774\ : Odrv4
    port map (
            O => \N__43658\,
            I => bit_cnt_0
        );

    \I__9773\ : LocalMux
    port map (
            O => \N__43655\,
            I => bit_cnt_0
        );

    \I__9772\ : Odrv12
    port map (
            O => \N__43652\,
            I => bit_cnt_0
        );

    \I__9771\ : InMux
    port map (
            O => \N__43645\,
            I => \N__43642\
        );

    \I__9770\ : LocalMux
    port map (
            O => \N__43642\,
            I => \N__43638\
        );

    \I__9769\ : InMux
    port map (
            O => \N__43641\,
            I => \N__43635\
        );

    \I__9768\ : Odrv4
    port map (
            O => \N__43638\,
            I => \comm_spi.n14624\
        );

    \I__9767\ : LocalMux
    port map (
            O => \N__43635\,
            I => \comm_spi.n14624\
        );

    \I__9766\ : SRMux
    port map (
            O => \N__43630\,
            I => \N__43627\
        );

    \I__9765\ : LocalMux
    port map (
            O => \N__43627\,
            I => \N__43624\
        );

    \I__9764\ : Span4Mux_v
    port map (
            O => \N__43624\,
            I => \N__43621\
        );

    \I__9763\ : Span4Mux_h
    port map (
            O => \N__43621\,
            I => \N__43618\
        );

    \I__9762\ : Span4Mux_v
    port map (
            O => \N__43618\,
            I => \N__43615\
        );

    \I__9761\ : Odrv4
    port map (
            O => \N__43615\,
            I => \comm_spi.data_tx_7__N_769\
        );

    \I__9760\ : InMux
    port map (
            O => \N__43612\,
            I => \N__43609\
        );

    \I__9759\ : LocalMux
    port map (
            O => \N__43609\,
            I => \comm_spi.n22626\
        );

    \I__9758\ : CascadeMux
    port map (
            O => \N__43606\,
            I => \comm_spi.n22626_cascade_\
        );

    \I__9757\ : InMux
    port map (
            O => \N__43603\,
            I => \N__43600\
        );

    \I__9756\ : LocalMux
    port map (
            O => \N__43600\,
            I => \N__43597\
        );

    \I__9755\ : Span4Mux_v
    port map (
            O => \N__43597\,
            I => \N__43594\
        );

    \I__9754\ : Odrv4
    port map (
            O => \N__43594\,
            I => \comm_spi.n14589\
        );

    \I__9753\ : IoInMux
    port map (
            O => \N__43591\,
            I => \N__43588\
        );

    \I__9752\ : LocalMux
    port map (
            O => \N__43588\,
            I => \N__43585\
        );

    \I__9751\ : Span4Mux_s1_h
    port map (
            O => \N__43585\,
            I => \N__43582\
        );

    \I__9750\ : Sp12to4
    port map (
            O => \N__43582\,
            I => \N__43579\
        );

    \I__9749\ : Span12Mux_s9_v
    port map (
            O => \N__43579\,
            I => \N__43576\
        );

    \I__9748\ : Odrv12
    port map (
            O => \N__43576\,
            I => \ICE_SPI_MISO\
        );

    \I__9747\ : InMux
    port map (
            O => \N__43573\,
            I => \N__43570\
        );

    \I__9746\ : LocalMux
    port map (
            O => \N__43570\,
            I => \N__43566\
        );

    \I__9745\ : InMux
    port map (
            O => \N__43569\,
            I => \N__43563\
        );

    \I__9744\ : Span4Mux_v
    port map (
            O => \N__43566\,
            I => \N__43559\
        );

    \I__9743\ : LocalMux
    port map (
            O => \N__43563\,
            I => \N__43556\
        );

    \I__9742\ : InMux
    port map (
            O => \N__43562\,
            I => \N__43553\
        );

    \I__9741\ : Odrv4
    port map (
            O => \N__43559\,
            I => \comm_spi.n22635\
        );

    \I__9740\ : Odrv12
    port map (
            O => \N__43556\,
            I => \comm_spi.n22635\
        );

    \I__9739\ : LocalMux
    port map (
            O => \N__43553\,
            I => \comm_spi.n22635\
        );

    \I__9738\ : InMux
    port map (
            O => \N__43546\,
            I => \N__43542\
        );

    \I__9737\ : InMux
    port map (
            O => \N__43545\,
            I => \N__43539\
        );

    \I__9736\ : LocalMux
    port map (
            O => \N__43542\,
            I => \comm_spi.n14623\
        );

    \I__9735\ : LocalMux
    port map (
            O => \N__43539\,
            I => \comm_spi.n14623\
        );

    \I__9734\ : CascadeMux
    port map (
            O => \N__43534\,
            I => \N__43529\
        );

    \I__9733\ : CascadeMux
    port map (
            O => \N__43533\,
            I => \N__43526\
        );

    \I__9732\ : CascadeMux
    port map (
            O => \N__43532\,
            I => \N__43521\
        );

    \I__9731\ : InMux
    port map (
            O => \N__43529\,
            I => \N__43517\
        );

    \I__9730\ : InMux
    port map (
            O => \N__43526\,
            I => \N__43514\
        );

    \I__9729\ : CascadeMux
    port map (
            O => \N__43525\,
            I => \N__43511\
        );

    \I__9728\ : InMux
    port map (
            O => \N__43524\,
            I => \N__43508\
        );

    \I__9727\ : InMux
    port map (
            O => \N__43521\,
            I => \N__43505\
        );

    \I__9726\ : InMux
    port map (
            O => \N__43520\,
            I => \N__43501\
        );

    \I__9725\ : LocalMux
    port map (
            O => \N__43517\,
            I => \N__43496\
        );

    \I__9724\ : LocalMux
    port map (
            O => \N__43514\,
            I => \N__43496\
        );

    \I__9723\ : InMux
    port map (
            O => \N__43511\,
            I => \N__43493\
        );

    \I__9722\ : LocalMux
    port map (
            O => \N__43508\,
            I => \N__43488\
        );

    \I__9721\ : LocalMux
    port map (
            O => \N__43505\,
            I => \N__43488\
        );

    \I__9720\ : CascadeMux
    port map (
            O => \N__43504\,
            I => \N__43484\
        );

    \I__9719\ : LocalMux
    port map (
            O => \N__43501\,
            I => \N__43481\
        );

    \I__9718\ : Span4Mux_v
    port map (
            O => \N__43496\,
            I => \N__43478\
        );

    \I__9717\ : LocalMux
    port map (
            O => \N__43493\,
            I => \N__43475\
        );

    \I__9716\ : Span4Mux_v
    port map (
            O => \N__43488\,
            I => \N__43471\
        );

    \I__9715\ : InMux
    port map (
            O => \N__43487\,
            I => \N__43468\
        );

    \I__9714\ : InMux
    port map (
            O => \N__43484\,
            I => \N__43465\
        );

    \I__9713\ : Span4Mux_h
    port map (
            O => \N__43481\,
            I => \N__43462\
        );

    \I__9712\ : Span4Mux_v
    port map (
            O => \N__43478\,
            I => \N__43456\
        );

    \I__9711\ : Span4Mux_h
    port map (
            O => \N__43475\,
            I => \N__43456\
        );

    \I__9710\ : InMux
    port map (
            O => \N__43474\,
            I => \N__43453\
        );

    \I__9709\ : Sp12to4
    port map (
            O => \N__43471\,
            I => \N__43450\
        );

    \I__9708\ : LocalMux
    port map (
            O => \N__43468\,
            I => \N__43447\
        );

    \I__9707\ : LocalMux
    port map (
            O => \N__43465\,
            I => \N__43444\
        );

    \I__9706\ : Span4Mux_v
    port map (
            O => \N__43462\,
            I => \N__43441\
        );

    \I__9705\ : InMux
    port map (
            O => \N__43461\,
            I => \N__43438\
        );

    \I__9704\ : Span4Mux_h
    port map (
            O => \N__43456\,
            I => \N__43435\
        );

    \I__9703\ : LocalMux
    port map (
            O => \N__43453\,
            I => \N__43428\
        );

    \I__9702\ : Span12Mux_h
    port map (
            O => \N__43450\,
            I => \N__43428\
        );

    \I__9701\ : Sp12to4
    port map (
            O => \N__43447\,
            I => \N__43428\
        );

    \I__9700\ : Odrv4
    port map (
            O => \N__43444\,
            I => comm_buf_0_0
        );

    \I__9699\ : Odrv4
    port map (
            O => \N__43441\,
            I => comm_buf_0_0
        );

    \I__9698\ : LocalMux
    port map (
            O => \N__43438\,
            I => comm_buf_0_0
        );

    \I__9697\ : Odrv4
    port map (
            O => \N__43435\,
            I => comm_buf_0_0
        );

    \I__9696\ : Odrv12
    port map (
            O => \N__43428\,
            I => comm_buf_0_0
        );

    \I__9695\ : InMux
    port map (
            O => \N__43417\,
            I => \N__43414\
        );

    \I__9694\ : LocalMux
    port map (
            O => \N__43414\,
            I => \N__43410\
        );

    \I__9693\ : InMux
    port map (
            O => \N__43413\,
            I => \N__43406\
        );

    \I__9692\ : Span4Mux_v
    port map (
            O => \N__43410\,
            I => \N__43403\
        );

    \I__9691\ : InMux
    port map (
            O => \N__43409\,
            I => \N__43400\
        );

    \I__9690\ : LocalMux
    port map (
            O => \N__43406\,
            I => \N__43397\
        );

    \I__9689\ : Odrv4
    port map (
            O => \N__43403\,
            I => buf_dds0_8
        );

    \I__9688\ : LocalMux
    port map (
            O => \N__43400\,
            I => buf_dds0_8
        );

    \I__9687\ : Odrv12
    port map (
            O => \N__43397\,
            I => buf_dds0_8
        );

    \I__9686\ : InMux
    port map (
            O => \N__43390\,
            I => \N__43387\
        );

    \I__9685\ : LocalMux
    port map (
            O => \N__43387\,
            I => \N__43384\
        );

    \I__9684\ : Span4Mux_v
    port map (
            O => \N__43384\,
            I => \N__43379\
        );

    \I__9683\ : InMux
    port map (
            O => \N__43383\,
            I => \N__43376\
        );

    \I__9682\ : InMux
    port map (
            O => \N__43382\,
            I => \N__43371\
        );

    \I__9681\ : Span4Mux_v
    port map (
            O => \N__43379\,
            I => \N__43366\
        );

    \I__9680\ : LocalMux
    port map (
            O => \N__43376\,
            I => \N__43366\
        );

    \I__9679\ : InMux
    port map (
            O => \N__43375\,
            I => \N__43363\
        );

    \I__9678\ : InMux
    port map (
            O => \N__43374\,
            I => \N__43360\
        );

    \I__9677\ : LocalMux
    port map (
            O => \N__43371\,
            I => \N__43357\
        );

    \I__9676\ : Span4Mux_v
    port map (
            O => \N__43366\,
            I => \N__43354\
        );

    \I__9675\ : LocalMux
    port map (
            O => \N__43363\,
            I => \N__43351\
        );

    \I__9674\ : LocalMux
    port map (
            O => \N__43360\,
            I => \N__43348\
        );

    \I__9673\ : Span4Mux_h
    port map (
            O => \N__43357\,
            I => \N__43344\
        );

    \I__9672\ : Span4Mux_h
    port map (
            O => \N__43354\,
            I => \N__43339\
        );

    \I__9671\ : Span4Mux_v
    port map (
            O => \N__43351\,
            I => \N__43339\
        );

    \I__9670\ : Span4Mux_v
    port map (
            O => \N__43348\,
            I => \N__43336\
        );

    \I__9669\ : InMux
    port map (
            O => \N__43347\,
            I => \N__43333\
        );

    \I__9668\ : Span4Mux_v
    port map (
            O => \N__43344\,
            I => \N__43328\
        );

    \I__9667\ : Span4Mux_v
    port map (
            O => \N__43339\,
            I => \N__43328\
        );

    \I__9666\ : Odrv4
    port map (
            O => \N__43336\,
            I => comm_buf_1_1
        );

    \I__9665\ : LocalMux
    port map (
            O => \N__43333\,
            I => comm_buf_1_1
        );

    \I__9664\ : Odrv4
    port map (
            O => \N__43328\,
            I => comm_buf_1_1
        );

    \I__9663\ : InMux
    port map (
            O => \N__43321\,
            I => \N__43316\
        );

    \I__9662\ : InMux
    port map (
            O => \N__43320\,
            I => \N__43313\
        );

    \I__9661\ : InMux
    port map (
            O => \N__43319\,
            I => \N__43310\
        );

    \I__9660\ : LocalMux
    port map (
            O => \N__43316\,
            I => \N__43305\
        );

    \I__9659\ : LocalMux
    port map (
            O => \N__43313\,
            I => \N__43305\
        );

    \I__9658\ : LocalMux
    port map (
            O => \N__43310\,
            I => data_index_1
        );

    \I__9657\ : Odrv4
    port map (
            O => \N__43305\,
            I => data_index_1
        );

    \I__9656\ : InMux
    port map (
            O => \N__43300\,
            I => \N__43296\
        );

    \I__9655\ : InMux
    port map (
            O => \N__43299\,
            I => \N__43292\
        );

    \I__9654\ : LocalMux
    port map (
            O => \N__43296\,
            I => \N__43288\
        );

    \I__9653\ : InMux
    port map (
            O => \N__43295\,
            I => \N__43285\
        );

    \I__9652\ : LocalMux
    port map (
            O => \N__43292\,
            I => \N__43281\
        );

    \I__9651\ : InMux
    port map (
            O => \N__43291\,
            I => \N__43278\
        );

    \I__9650\ : Span4Mux_h
    port map (
            O => \N__43288\,
            I => \N__43268\
        );

    \I__9649\ : LocalMux
    port map (
            O => \N__43285\,
            I => \N__43268\
        );

    \I__9648\ : InMux
    port map (
            O => \N__43284\,
            I => \N__43265\
        );

    \I__9647\ : Span4Mux_v
    port map (
            O => \N__43281\,
            I => \N__43260\
        );

    \I__9646\ : LocalMux
    port map (
            O => \N__43278\,
            I => \N__43260\
        );

    \I__9645\ : InMux
    port map (
            O => \N__43277\,
            I => \N__43257\
        );

    \I__9644\ : InMux
    port map (
            O => \N__43276\,
            I => \N__43254\
        );

    \I__9643\ : InMux
    port map (
            O => \N__43275\,
            I => \N__43249\
        );

    \I__9642\ : InMux
    port map (
            O => \N__43274\,
            I => \N__43249\
        );

    \I__9641\ : InMux
    port map (
            O => \N__43273\,
            I => \N__43246\
        );

    \I__9640\ : Span4Mux_h
    port map (
            O => \N__43268\,
            I => \N__43243\
        );

    \I__9639\ : LocalMux
    port map (
            O => \N__43265\,
            I => n8780
        );

    \I__9638\ : Odrv4
    port map (
            O => \N__43260\,
            I => n8780
        );

    \I__9637\ : LocalMux
    port map (
            O => \N__43257\,
            I => n8780
        );

    \I__9636\ : LocalMux
    port map (
            O => \N__43254\,
            I => n8780
        );

    \I__9635\ : LocalMux
    port map (
            O => \N__43249\,
            I => n8780
        );

    \I__9634\ : LocalMux
    port map (
            O => \N__43246\,
            I => n8780
        );

    \I__9633\ : Odrv4
    port map (
            O => \N__43243\,
            I => n8780
        );

    \I__9632\ : InMux
    port map (
            O => \N__43228\,
            I => \N__43225\
        );

    \I__9631\ : LocalMux
    port map (
            O => \N__43225\,
            I => n8_adj_1547
        );

    \I__9630\ : CascadeMux
    port map (
            O => \N__43222\,
            I => \n8_adj_1547_cascade_\
        );

    \I__9629\ : InMux
    port map (
            O => \N__43219\,
            I => \N__43213\
        );

    \I__9628\ : InMux
    port map (
            O => \N__43218\,
            I => \N__43213\
        );

    \I__9627\ : LocalMux
    port map (
            O => \N__43213\,
            I => \N__43210\
        );

    \I__9626\ : Odrv12
    port map (
            O => \N__43210\,
            I => n7_adj_1546
        );

    \I__9625\ : CascadeMux
    port map (
            O => \N__43207\,
            I => \N__43204\
        );

    \I__9624\ : CascadeBuf
    port map (
            O => \N__43204\,
            I => \N__43201\
        );

    \I__9623\ : CascadeMux
    port map (
            O => \N__43201\,
            I => \N__43198\
        );

    \I__9622\ : CascadeBuf
    port map (
            O => \N__43198\,
            I => \N__43195\
        );

    \I__9621\ : CascadeMux
    port map (
            O => \N__43195\,
            I => \N__43192\
        );

    \I__9620\ : CascadeBuf
    port map (
            O => \N__43192\,
            I => \N__43189\
        );

    \I__9619\ : CascadeMux
    port map (
            O => \N__43189\,
            I => \N__43186\
        );

    \I__9618\ : CascadeBuf
    port map (
            O => \N__43186\,
            I => \N__43183\
        );

    \I__9617\ : CascadeMux
    port map (
            O => \N__43183\,
            I => \N__43180\
        );

    \I__9616\ : CascadeBuf
    port map (
            O => \N__43180\,
            I => \N__43177\
        );

    \I__9615\ : CascadeMux
    port map (
            O => \N__43177\,
            I => \N__43174\
        );

    \I__9614\ : CascadeBuf
    port map (
            O => \N__43174\,
            I => \N__43171\
        );

    \I__9613\ : CascadeMux
    port map (
            O => \N__43171\,
            I => \N__43168\
        );

    \I__9612\ : CascadeBuf
    port map (
            O => \N__43168\,
            I => \N__43165\
        );

    \I__9611\ : CascadeMux
    port map (
            O => \N__43165\,
            I => \N__43162\
        );

    \I__9610\ : CascadeBuf
    port map (
            O => \N__43162\,
            I => \N__43159\
        );

    \I__9609\ : CascadeMux
    port map (
            O => \N__43159\,
            I => \N__43155\
        );

    \I__9608\ : CascadeMux
    port map (
            O => \N__43158\,
            I => \N__43152\
        );

    \I__9607\ : CascadeBuf
    port map (
            O => \N__43155\,
            I => \N__43149\
        );

    \I__9606\ : CascadeBuf
    port map (
            O => \N__43152\,
            I => \N__43146\
        );

    \I__9605\ : CascadeMux
    port map (
            O => \N__43149\,
            I => \N__43143\
        );

    \I__9604\ : CascadeMux
    port map (
            O => \N__43146\,
            I => \N__43140\
        );

    \I__9603\ : InMux
    port map (
            O => \N__43143\,
            I => \N__43137\
        );

    \I__9602\ : InMux
    port map (
            O => \N__43140\,
            I => \N__43134\
        );

    \I__9601\ : LocalMux
    port map (
            O => \N__43137\,
            I => \N__43131\
        );

    \I__9600\ : LocalMux
    port map (
            O => \N__43134\,
            I => \N__43128\
        );

    \I__9599\ : Span4Mux_v
    port map (
            O => \N__43131\,
            I => \N__43125\
        );

    \I__9598\ : Span4Mux_v
    port map (
            O => \N__43128\,
            I => \N__43122\
        );

    \I__9597\ : Span4Mux_h
    port map (
            O => \N__43125\,
            I => \N__43119\
        );

    \I__9596\ : Span4Mux_h
    port map (
            O => \N__43122\,
            I => \N__43116\
        );

    \I__9595\ : Span4Mux_h
    port map (
            O => \N__43119\,
            I => \N__43113\
        );

    \I__9594\ : Odrv4
    port map (
            O => \N__43116\,
            I => \data_index_9_N_212_1\
        );

    \I__9593\ : Odrv4
    port map (
            O => \N__43113\,
            I => \data_index_9_N_212_1\
        );

    \I__9592\ : CascadeMux
    port map (
            O => \N__43108\,
            I => \N__43105\
        );

    \I__9591\ : InMux
    port map (
            O => \N__43105\,
            I => \N__43101\
        );

    \I__9590\ : CascadeMux
    port map (
            O => \N__43104\,
            I => \N__43098\
        );

    \I__9589\ : LocalMux
    port map (
            O => \N__43101\,
            I => \N__43094\
        );

    \I__9588\ : InMux
    port map (
            O => \N__43098\,
            I => \N__43091\
        );

    \I__9587\ : CascadeMux
    port map (
            O => \N__43097\,
            I => \N__43088\
        );

    \I__9586\ : Span4Mux_v
    port map (
            O => \N__43094\,
            I => \N__43085\
        );

    \I__9585\ : LocalMux
    port map (
            O => \N__43091\,
            I => \N__43082\
        );

    \I__9584\ : InMux
    port map (
            O => \N__43088\,
            I => \N__43079\
        );

    \I__9583\ : Span4Mux_h
    port map (
            O => \N__43085\,
            I => \N__43076\
        );

    \I__9582\ : Span12Mux_h
    port map (
            O => \N__43082\,
            I => \N__43073\
        );

    \I__9581\ : LocalMux
    port map (
            O => \N__43079\,
            I => buf_dds0_11
        );

    \I__9580\ : Odrv4
    port map (
            O => \N__43076\,
            I => buf_dds0_11
        );

    \I__9579\ : Odrv12
    port map (
            O => \N__43073\,
            I => buf_dds0_11
        );

    \I__9578\ : InMux
    port map (
            O => \N__43066\,
            I => \N__43062\
        );

    \I__9577\ : InMux
    port map (
            O => \N__43065\,
            I => \N__43059\
        );

    \I__9576\ : LocalMux
    port map (
            O => \N__43062\,
            I => \N__43056\
        );

    \I__9575\ : LocalMux
    port map (
            O => \N__43059\,
            I => \N__43050\
        );

    \I__9574\ : Span4Mux_h
    port map (
            O => \N__43056\,
            I => \N__43050\
        );

    \I__9573\ : InMux
    port map (
            O => \N__43055\,
            I => \N__43047\
        );

    \I__9572\ : Span4Mux_h
    port map (
            O => \N__43050\,
            I => \N__43044\
        );

    \I__9571\ : LocalMux
    port map (
            O => \N__43047\,
            I => buf_dds0_5
        );

    \I__9570\ : Odrv4
    port map (
            O => \N__43044\,
            I => buf_dds0_5
        );

    \I__9569\ : InMux
    port map (
            O => \N__43039\,
            I => \N__43035\
        );

    \I__9568\ : InMux
    port map (
            O => \N__43038\,
            I => \N__43032\
        );

    \I__9567\ : LocalMux
    port map (
            O => \N__43035\,
            I => \N__43029\
        );

    \I__9566\ : LocalMux
    port map (
            O => \N__43032\,
            I => n8_adj_1532
        );

    \I__9565\ : Odrv4
    port map (
            O => \N__43029\,
            I => n8_adj_1532
        );

    \I__9564\ : InMux
    port map (
            O => \N__43024\,
            I => \N__43020\
        );

    \I__9563\ : InMux
    port map (
            O => \N__43023\,
            I => \N__43017\
        );

    \I__9562\ : LocalMux
    port map (
            O => \N__43020\,
            I => \N__43014\
        );

    \I__9561\ : LocalMux
    port map (
            O => \N__43017\,
            I => n7_adj_1531
        );

    \I__9560\ : Odrv12
    port map (
            O => \N__43014\,
            I => n7_adj_1531
        );

    \I__9559\ : CascadeMux
    port map (
            O => \N__43009\,
            I => \N__43006\
        );

    \I__9558\ : CascadeBuf
    port map (
            O => \N__43006\,
            I => \N__43003\
        );

    \I__9557\ : CascadeMux
    port map (
            O => \N__43003\,
            I => \N__43000\
        );

    \I__9556\ : CascadeBuf
    port map (
            O => \N__43000\,
            I => \N__42997\
        );

    \I__9555\ : CascadeMux
    port map (
            O => \N__42997\,
            I => \N__42994\
        );

    \I__9554\ : CascadeBuf
    port map (
            O => \N__42994\,
            I => \N__42991\
        );

    \I__9553\ : CascadeMux
    port map (
            O => \N__42991\,
            I => \N__42988\
        );

    \I__9552\ : CascadeBuf
    port map (
            O => \N__42988\,
            I => \N__42985\
        );

    \I__9551\ : CascadeMux
    port map (
            O => \N__42985\,
            I => \N__42982\
        );

    \I__9550\ : CascadeBuf
    port map (
            O => \N__42982\,
            I => \N__42979\
        );

    \I__9549\ : CascadeMux
    port map (
            O => \N__42979\,
            I => \N__42976\
        );

    \I__9548\ : CascadeBuf
    port map (
            O => \N__42976\,
            I => \N__42973\
        );

    \I__9547\ : CascadeMux
    port map (
            O => \N__42973\,
            I => \N__42970\
        );

    \I__9546\ : CascadeBuf
    port map (
            O => \N__42970\,
            I => \N__42967\
        );

    \I__9545\ : CascadeMux
    port map (
            O => \N__42967\,
            I => \N__42963\
        );

    \I__9544\ : CascadeMux
    port map (
            O => \N__42966\,
            I => \N__42960\
        );

    \I__9543\ : CascadeBuf
    port map (
            O => \N__42963\,
            I => \N__42957\
        );

    \I__9542\ : CascadeBuf
    port map (
            O => \N__42960\,
            I => \N__42954\
        );

    \I__9541\ : CascadeMux
    port map (
            O => \N__42957\,
            I => \N__42951\
        );

    \I__9540\ : CascadeMux
    port map (
            O => \N__42954\,
            I => \N__42948\
        );

    \I__9539\ : CascadeBuf
    port map (
            O => \N__42951\,
            I => \N__42945\
        );

    \I__9538\ : InMux
    port map (
            O => \N__42948\,
            I => \N__42942\
        );

    \I__9537\ : CascadeMux
    port map (
            O => \N__42945\,
            I => \N__42939\
        );

    \I__9536\ : LocalMux
    port map (
            O => \N__42942\,
            I => \N__42936\
        );

    \I__9535\ : InMux
    port map (
            O => \N__42939\,
            I => \N__42933\
        );

    \I__9534\ : Span4Mux_v
    port map (
            O => \N__42936\,
            I => \N__42930\
        );

    \I__9533\ : LocalMux
    port map (
            O => \N__42933\,
            I => \N__42927\
        );

    \I__9532\ : Span4Mux_h
    port map (
            O => \N__42930\,
            I => \N__42924\
        );

    \I__9531\ : Span12Mux_h
    port map (
            O => \N__42927\,
            I => \N__42921\
        );

    \I__9530\ : Odrv4
    port map (
            O => \N__42924\,
            I => \data_index_9_N_212_9\
        );

    \I__9529\ : Odrv12
    port map (
            O => \N__42921\,
            I => \data_index_9_N_212_9\
        );

    \I__9528\ : CascadeMux
    port map (
            O => \N__42916\,
            I => \N__42912\
        );

    \I__9527\ : InMux
    port map (
            O => \N__42915\,
            I => \N__42909\
        );

    \I__9526\ : InMux
    port map (
            O => \N__42912\,
            I => \N__42906\
        );

    \I__9525\ : LocalMux
    port map (
            O => \N__42909\,
            I => tmp_buf_15
        );

    \I__9524\ : LocalMux
    port map (
            O => \N__42906\,
            I => tmp_buf_15
        );

    \I__9523\ : IoInMux
    port map (
            O => \N__42901\,
            I => \N__42898\
        );

    \I__9522\ : LocalMux
    port map (
            O => \N__42898\,
            I => \N__42895\
        );

    \I__9521\ : IoSpan4Mux
    port map (
            O => \N__42895\,
            I => \N__42892\
        );

    \I__9520\ : Span4Mux_s3_v
    port map (
            O => \N__42892\,
            I => \N__42889\
        );

    \I__9519\ : Span4Mux_h
    port map (
            O => \N__42889\,
            I => \N__42886\
        );

    \I__9518\ : Span4Mux_v
    port map (
            O => \N__42886\,
            I => \N__42882\
        );

    \I__9517\ : InMux
    port map (
            O => \N__42885\,
            I => \N__42879\
        );

    \I__9516\ : Odrv4
    port map (
            O => \N__42882\,
            I => \DDS_MOSI\
        );

    \I__9515\ : LocalMux
    port map (
            O => \N__42879\,
            I => \DDS_MOSI\
        );

    \I__9514\ : InMux
    port map (
            O => \N__42874\,
            I => \N__42870\
        );

    \I__9513\ : InMux
    port map (
            O => \N__42873\,
            I => \N__42867\
        );

    \I__9512\ : LocalMux
    port map (
            O => \N__42870\,
            I => \N__42864\
        );

    \I__9511\ : LocalMux
    port map (
            O => \N__42867\,
            I => n7_adj_1515
        );

    \I__9510\ : Odrv12
    port map (
            O => \N__42864\,
            I => n7_adj_1515
        );

    \I__9509\ : InMux
    port map (
            O => \N__42859\,
            I => \N__42856\
        );

    \I__9508\ : LocalMux
    port map (
            O => \N__42856\,
            I => \N__42852\
        );

    \I__9507\ : InMux
    port map (
            O => \N__42855\,
            I => \N__42849\
        );

    \I__9506\ : Span4Mux_h
    port map (
            O => \N__42852\,
            I => \N__42846\
        );

    \I__9505\ : LocalMux
    port map (
            O => \N__42849\,
            I => n17314
        );

    \I__9504\ : Odrv4
    port map (
            O => \N__42846\,
            I => n17314
        );

    \I__9503\ : InMux
    port map (
            O => \N__42841\,
            I => \N__42836\
        );

    \I__9502\ : InMux
    port map (
            O => \N__42840\,
            I => \N__42833\
        );

    \I__9501\ : InMux
    port map (
            O => \N__42839\,
            I => \N__42830\
        );

    \I__9500\ : LocalMux
    port map (
            O => \N__42836\,
            I => data_index_0
        );

    \I__9499\ : LocalMux
    port map (
            O => \N__42833\,
            I => data_index_0
        );

    \I__9498\ : LocalMux
    port map (
            O => \N__42830\,
            I => data_index_0
        );

    \I__9497\ : CascadeMux
    port map (
            O => \N__42823\,
            I => \N__42819\
        );

    \I__9496\ : CascadeMux
    port map (
            O => \N__42822\,
            I => \N__42816\
        );

    \I__9495\ : InMux
    port map (
            O => \N__42819\,
            I => \N__42812\
        );

    \I__9494\ : InMux
    port map (
            O => \N__42816\,
            I => \N__42809\
        );

    \I__9493\ : InMux
    port map (
            O => \N__42815\,
            I => \N__42805\
        );

    \I__9492\ : LocalMux
    port map (
            O => \N__42812\,
            I => \N__42801\
        );

    \I__9491\ : LocalMux
    port map (
            O => \N__42809\,
            I => \N__42798\
        );

    \I__9490\ : CascadeMux
    port map (
            O => \N__42808\,
            I => \N__42795\
        );

    \I__9489\ : LocalMux
    port map (
            O => \N__42805\,
            I => \N__42792\
        );

    \I__9488\ : InMux
    port map (
            O => \N__42804\,
            I => \N__42789\
        );

    \I__9487\ : Span4Mux_v
    port map (
            O => \N__42801\,
            I => \N__42785\
        );

    \I__9486\ : Span4Mux_h
    port map (
            O => \N__42798\,
            I => \N__42782\
        );

    \I__9485\ : InMux
    port map (
            O => \N__42795\,
            I => \N__42779\
        );

    \I__9484\ : Span4Mux_h
    port map (
            O => \N__42792\,
            I => \N__42774\
        );

    \I__9483\ : LocalMux
    port map (
            O => \N__42789\,
            I => \N__42774\
        );

    \I__9482\ : InMux
    port map (
            O => \N__42788\,
            I => \N__42771\
        );

    \I__9481\ : Sp12to4
    port map (
            O => \N__42785\,
            I => \N__42768\
        );

    \I__9480\ : Span4Mux_v
    port map (
            O => \N__42782\,
            I => \N__42759\
        );

    \I__9479\ : LocalMux
    port map (
            O => \N__42779\,
            I => \N__42759\
        );

    \I__9478\ : Span4Mux_v
    port map (
            O => \N__42774\,
            I => \N__42759\
        );

    \I__9477\ : LocalMux
    port map (
            O => \N__42771\,
            I => \N__42759\
        );

    \I__9476\ : Odrv12
    port map (
            O => \N__42768\,
            I => comm_buf_1_2
        );

    \I__9475\ : Odrv4
    port map (
            O => \N__42759\,
            I => comm_buf_1_2
        );

    \I__9474\ : InMux
    port map (
            O => \N__42754\,
            I => \N__42750\
        );

    \I__9473\ : InMux
    port map (
            O => \N__42753\,
            I => \N__42747\
        );

    \I__9472\ : LocalMux
    port map (
            O => \N__42750\,
            I => \N__42743\
        );

    \I__9471\ : LocalMux
    port map (
            O => \N__42747\,
            I => \N__42740\
        );

    \I__9470\ : InMux
    port map (
            O => \N__42746\,
            I => \N__42737\
        );

    \I__9469\ : Span4Mux_v
    port map (
            O => \N__42743\,
            I => \N__42732\
        );

    \I__9468\ : Span4Mux_h
    port map (
            O => \N__42740\,
            I => \N__42732\
        );

    \I__9467\ : LocalMux
    port map (
            O => \N__42737\,
            I => buf_dds0_2
        );

    \I__9466\ : Odrv4
    port map (
            O => \N__42732\,
            I => buf_dds0_2
        );

    \I__9465\ : InMux
    port map (
            O => \N__42727\,
            I => \N__42720\
        );

    \I__9464\ : InMux
    port map (
            O => \N__42726\,
            I => \N__42720\
        );

    \I__9463\ : InMux
    port map (
            O => \N__42725\,
            I => \N__42717\
        );

    \I__9462\ : LocalMux
    port map (
            O => \N__42720\,
            I => data_index_9
        );

    \I__9461\ : LocalMux
    port map (
            O => \N__42717\,
            I => data_index_9
        );

    \I__9460\ : InMux
    port map (
            O => \N__42712\,
            I => \N__42708\
        );

    \I__9459\ : InMux
    port map (
            O => \N__42711\,
            I => \N__42705\
        );

    \I__9458\ : LocalMux
    port map (
            O => \N__42708\,
            I => \N__42702\
        );

    \I__9457\ : LocalMux
    port map (
            O => \N__42705\,
            I => \N__42698\
        );

    \I__9456\ : Span4Mux_h
    port map (
            O => \N__42702\,
            I => \N__42695\
        );

    \I__9455\ : InMux
    port map (
            O => \N__42701\,
            I => \N__42692\
        );

    \I__9454\ : Span4Mux_h
    port map (
            O => \N__42698\,
            I => \N__42689\
        );

    \I__9453\ : Odrv4
    port map (
            O => \N__42695\,
            I => buf_dds0_4
        );

    \I__9452\ : LocalMux
    port map (
            O => \N__42692\,
            I => buf_dds0_4
        );

    \I__9451\ : Odrv4
    port map (
            O => \N__42689\,
            I => buf_dds0_4
        );

    \I__9450\ : CascadeMux
    port map (
            O => \N__42682\,
            I => \n8_adj_1538_cascade_\
        );

    \I__9449\ : InMux
    port map (
            O => \N__42679\,
            I => \N__42674\
        );

    \I__9448\ : InMux
    port map (
            O => \N__42678\,
            I => \N__42671\
        );

    \I__9447\ : InMux
    port map (
            O => \N__42677\,
            I => \N__42668\
        );

    \I__9446\ : LocalMux
    port map (
            O => \N__42674\,
            I => \N__42663\
        );

    \I__9445\ : LocalMux
    port map (
            O => \N__42671\,
            I => \N__42663\
        );

    \I__9444\ : LocalMux
    port map (
            O => \N__42668\,
            I => data_index_6
        );

    \I__9443\ : Odrv4
    port map (
            O => \N__42663\,
            I => data_index_6
        );

    \I__9442\ : InMux
    port map (
            O => \N__42658\,
            I => \N__42655\
        );

    \I__9441\ : LocalMux
    port map (
            O => \N__42655\,
            I => \N__42651\
        );

    \I__9440\ : InMux
    port map (
            O => \N__42654\,
            I => \N__42648\
        );

    \I__9439\ : Span4Mux_h
    port map (
            O => \N__42651\,
            I => \N__42645\
        );

    \I__9438\ : LocalMux
    port map (
            O => \N__42648\,
            I => \N__42641\
        );

    \I__9437\ : Sp12to4
    port map (
            O => \N__42645\,
            I => \N__42638\
        );

    \I__9436\ : InMux
    port map (
            O => \N__42644\,
            I => \N__42635\
        );

    \I__9435\ : Span4Mux_h
    port map (
            O => \N__42641\,
            I => \N__42632\
        );

    \I__9434\ : Odrv12
    port map (
            O => \N__42638\,
            I => buf_dds0_6
        );

    \I__9433\ : LocalMux
    port map (
            O => \N__42635\,
            I => buf_dds0_6
        );

    \I__9432\ : Odrv4
    port map (
            O => \N__42632\,
            I => buf_dds0_6
        );

    \I__9431\ : CascadeMux
    port map (
            O => \N__42625\,
            I => \N__42620\
        );

    \I__9430\ : InMux
    port map (
            O => \N__42624\,
            I => \N__42616\
        );

    \I__9429\ : InMux
    port map (
            O => \N__42623\,
            I => \N__42612\
        );

    \I__9428\ : InMux
    port map (
            O => \N__42620\,
            I => \N__42609\
        );

    \I__9427\ : CascadeMux
    port map (
            O => \N__42619\,
            I => \N__42606\
        );

    \I__9426\ : LocalMux
    port map (
            O => \N__42616\,
            I => \N__42603\
        );

    \I__9425\ : CascadeMux
    port map (
            O => \N__42615\,
            I => \N__42600\
        );

    \I__9424\ : LocalMux
    port map (
            O => \N__42612\,
            I => \N__42597\
        );

    \I__9423\ : LocalMux
    port map (
            O => \N__42609\,
            I => \N__42593\
        );

    \I__9422\ : InMux
    port map (
            O => \N__42606\,
            I => \N__42590\
        );

    \I__9421\ : Span4Mux_h
    port map (
            O => \N__42603\,
            I => \N__42587\
        );

    \I__9420\ : InMux
    port map (
            O => \N__42600\,
            I => \N__42584\
        );

    \I__9419\ : Span4Mux_v
    port map (
            O => \N__42597\,
            I => \N__42581\
        );

    \I__9418\ : InMux
    port map (
            O => \N__42596\,
            I => \N__42578\
        );

    \I__9417\ : Span4Mux_v
    port map (
            O => \N__42593\,
            I => \N__42575\
        );

    \I__9416\ : LocalMux
    port map (
            O => \N__42590\,
            I => \N__42570\
        );

    \I__9415\ : Span4Mux_v
    port map (
            O => \N__42587\,
            I => \N__42570\
        );

    \I__9414\ : LocalMux
    port map (
            O => \N__42584\,
            I => \N__42567\
        );

    \I__9413\ : Span4Mux_v
    port map (
            O => \N__42581\,
            I => \N__42562\
        );

    \I__9412\ : LocalMux
    port map (
            O => \N__42578\,
            I => \N__42562\
        );

    \I__9411\ : Span4Mux_h
    port map (
            O => \N__42575\,
            I => \N__42559\
        );

    \I__9410\ : Span4Mux_v
    port map (
            O => \N__42570\,
            I => \N__42556\
        );

    \I__9409\ : Span4Mux_h
    port map (
            O => \N__42567\,
            I => \N__42551\
        );

    \I__9408\ : Span4Mux_h
    port map (
            O => \N__42562\,
            I => \N__42551\
        );

    \I__9407\ : Odrv4
    port map (
            O => \N__42559\,
            I => comm_buf_1_7
        );

    \I__9406\ : Odrv4
    port map (
            O => \N__42556\,
            I => comm_buf_1_7
        );

    \I__9405\ : Odrv4
    port map (
            O => \N__42551\,
            I => comm_buf_1_7
        );

    \I__9404\ : InMux
    port map (
            O => \N__42544\,
            I => \N__42540\
        );

    \I__9403\ : InMux
    port map (
            O => \N__42543\,
            I => \N__42537\
        );

    \I__9402\ : LocalMux
    port map (
            O => \N__42540\,
            I => \N__42534\
        );

    \I__9401\ : LocalMux
    port map (
            O => \N__42537\,
            I => \N__42531\
        );

    \I__9400\ : Span4Mux_v
    port map (
            O => \N__42534\,
            I => \N__42527\
        );

    \I__9399\ : Span4Mux_v
    port map (
            O => \N__42531\,
            I => \N__42524\
        );

    \I__9398\ : InMux
    port map (
            O => \N__42530\,
            I => \N__42521\
        );

    \I__9397\ : Span4Mux_h
    port map (
            O => \N__42527\,
            I => \N__42518\
        );

    \I__9396\ : Span4Mux_h
    port map (
            O => \N__42524\,
            I => \N__42515\
        );

    \I__9395\ : LocalMux
    port map (
            O => \N__42521\,
            I => buf_dds1_7
        );

    \I__9394\ : Odrv4
    port map (
            O => \N__42518\,
            I => buf_dds1_7
        );

    \I__9393\ : Odrv4
    port map (
            O => \N__42515\,
            I => buf_dds1_7
        );

    \I__9392\ : InMux
    port map (
            O => \N__42508\,
            I => \N__42503\
        );

    \I__9391\ : InMux
    port map (
            O => \N__42507\,
            I => \N__42500\
        );

    \I__9390\ : InMux
    port map (
            O => \N__42506\,
            I => \N__42497\
        );

    \I__9389\ : LocalMux
    port map (
            O => \N__42503\,
            I => data_index_4
        );

    \I__9388\ : LocalMux
    port map (
            O => \N__42500\,
            I => data_index_4
        );

    \I__9387\ : LocalMux
    port map (
            O => \N__42497\,
            I => data_index_4
        );

    \I__9386\ : InMux
    port map (
            O => \N__42490\,
            I => \N__42484\
        );

    \I__9385\ : InMux
    port map (
            O => \N__42489\,
            I => \N__42484\
        );

    \I__9384\ : LocalMux
    port map (
            O => \N__42484\,
            I => n7_adj_1540
        );

    \I__9383\ : InMux
    port map (
            O => \N__42481\,
            I => n19329
        );

    \I__9382\ : InMux
    port map (
            O => \N__42478\,
            I => n19330
        );

    \I__9381\ : InMux
    port map (
            O => \N__42475\,
            I => n19331
        );

    \I__9380\ : InMux
    port map (
            O => \N__42472\,
            I => \N__42468\
        );

    \I__9379\ : InMux
    port map (
            O => \N__42471\,
            I => \N__42465\
        );

    \I__9378\ : LocalMux
    port map (
            O => \N__42468\,
            I => \N__42460\
        );

    \I__9377\ : LocalMux
    port map (
            O => \N__42465\,
            I => \N__42460\
        );

    \I__9376\ : Span4Mux_h
    port map (
            O => \N__42460\,
            I => \N__42456\
        );

    \I__9375\ : InMux
    port map (
            O => \N__42459\,
            I => \N__42453\
        );

    \I__9374\ : Span4Mux_h
    port map (
            O => \N__42456\,
            I => \N__42450\
        );

    \I__9373\ : LocalMux
    port map (
            O => \N__42453\,
            I => \N__42447\
        );

    \I__9372\ : Span4Mux_h
    port map (
            O => \N__42450\,
            I => \N__42444\
        );

    \I__9371\ : Odrv12
    port map (
            O => \N__42447\,
            I => data_index_7
        );

    \I__9370\ : Odrv4
    port map (
            O => \N__42444\,
            I => data_index_7
        );

    \I__9369\ : InMux
    port map (
            O => \N__42439\,
            I => \N__42436\
        );

    \I__9368\ : LocalMux
    port map (
            O => \N__42436\,
            I => \N__42432\
        );

    \I__9367\ : InMux
    port map (
            O => \N__42435\,
            I => \N__42429\
        );

    \I__9366\ : Span4Mux_h
    port map (
            O => \N__42432\,
            I => \N__42426\
        );

    \I__9365\ : LocalMux
    port map (
            O => \N__42429\,
            I => \N__42423\
        );

    \I__9364\ : Span4Mux_h
    port map (
            O => \N__42426\,
            I => \N__42420\
        );

    \I__9363\ : Span12Mux_s11_v
    port map (
            O => \N__42423\,
            I => \N__42417\
        );

    \I__9362\ : Odrv4
    port map (
            O => \N__42420\,
            I => n7_adj_1535
        );

    \I__9361\ : Odrv12
    port map (
            O => \N__42417\,
            I => n7_adj_1535
        );

    \I__9360\ : InMux
    port map (
            O => \N__42412\,
            I => n19332
        );

    \I__9359\ : InMux
    port map (
            O => \N__42409\,
            I => \N__42405\
        );

    \I__9358\ : InMux
    port map (
            O => \N__42408\,
            I => \N__42402\
        );

    \I__9357\ : LocalMux
    port map (
            O => \N__42405\,
            I => \N__42397\
        );

    \I__9356\ : LocalMux
    port map (
            O => \N__42402\,
            I => \N__42397\
        );

    \I__9355\ : Span4Mux_v
    port map (
            O => \N__42397\,
            I => \N__42393\
        );

    \I__9354\ : InMux
    port map (
            O => \N__42396\,
            I => \N__42390\
        );

    \I__9353\ : Span4Mux_h
    port map (
            O => \N__42393\,
            I => \N__42387\
        );

    \I__9352\ : LocalMux
    port map (
            O => \N__42390\,
            I => data_index_8
        );

    \I__9351\ : Odrv4
    port map (
            O => \N__42387\,
            I => data_index_8
        );

    \I__9350\ : InMux
    port map (
            O => \N__42382\,
            I => \N__42376\
        );

    \I__9349\ : InMux
    port map (
            O => \N__42381\,
            I => \N__42376\
        );

    \I__9348\ : LocalMux
    port map (
            O => \N__42376\,
            I => \N__42373\
        );

    \I__9347\ : Span4Mux_v
    port map (
            O => \N__42373\,
            I => \N__42370\
        );

    \I__9346\ : Span4Mux_h
    port map (
            O => \N__42370\,
            I => \N__42367\
        );

    \I__9345\ : Span4Mux_h
    port map (
            O => \N__42367\,
            I => \N__42364\
        );

    \I__9344\ : Odrv4
    port map (
            O => \N__42364\,
            I => n7_adj_1533
        );

    \I__9343\ : InMux
    port map (
            O => \N__42361\,
            I => \bfn_16_16_0_\
        );

    \I__9342\ : CascadeMux
    port map (
            O => \N__42358\,
            I => \N__42354\
        );

    \I__9341\ : CascadeMux
    port map (
            O => \N__42357\,
            I => \N__42350\
        );

    \I__9340\ : InMux
    port map (
            O => \N__42354\,
            I => \N__42347\
        );

    \I__9339\ : CascadeMux
    port map (
            O => \N__42353\,
            I => \N__42336\
        );

    \I__9338\ : InMux
    port map (
            O => \N__42350\,
            I => \N__42333\
        );

    \I__9337\ : LocalMux
    port map (
            O => \N__42347\,
            I => \N__42330\
        );

    \I__9336\ : CascadeMux
    port map (
            O => \N__42346\,
            I => \N__42327\
        );

    \I__9335\ : CascadeMux
    port map (
            O => \N__42345\,
            I => \N__42324\
        );

    \I__9334\ : CascadeMux
    port map (
            O => \N__42344\,
            I => \N__42321\
        );

    \I__9333\ : CascadeMux
    port map (
            O => \N__42343\,
            I => \N__42318\
        );

    \I__9332\ : CascadeMux
    port map (
            O => \N__42342\,
            I => \N__42315\
        );

    \I__9331\ : CascadeMux
    port map (
            O => \N__42341\,
            I => \N__42312\
        );

    \I__9330\ : CascadeMux
    port map (
            O => \N__42340\,
            I => \N__42309\
        );

    \I__9329\ : CascadeMux
    port map (
            O => \N__42339\,
            I => \N__42306\
        );

    \I__9328\ : InMux
    port map (
            O => \N__42336\,
            I => \N__42303\
        );

    \I__9327\ : LocalMux
    port map (
            O => \N__42333\,
            I => \N__42300\
        );

    \I__9326\ : Span4Mux_v
    port map (
            O => \N__42330\,
            I => \N__42297\
        );

    \I__9325\ : InMux
    port map (
            O => \N__42327\,
            I => \N__42288\
        );

    \I__9324\ : InMux
    port map (
            O => \N__42324\,
            I => \N__42288\
        );

    \I__9323\ : InMux
    port map (
            O => \N__42321\,
            I => \N__42288\
        );

    \I__9322\ : InMux
    port map (
            O => \N__42318\,
            I => \N__42288\
        );

    \I__9321\ : InMux
    port map (
            O => \N__42315\,
            I => \N__42279\
        );

    \I__9320\ : InMux
    port map (
            O => \N__42312\,
            I => \N__42279\
        );

    \I__9319\ : InMux
    port map (
            O => \N__42309\,
            I => \N__42279\
        );

    \I__9318\ : InMux
    port map (
            O => \N__42306\,
            I => \N__42279\
        );

    \I__9317\ : LocalMux
    port map (
            O => \N__42303\,
            I => n10579
        );

    \I__9316\ : Odrv4
    port map (
            O => \N__42300\,
            I => n10579
        );

    \I__9315\ : Odrv4
    port map (
            O => \N__42297\,
            I => n10579
        );

    \I__9314\ : LocalMux
    port map (
            O => \N__42288\,
            I => n10579
        );

    \I__9313\ : LocalMux
    port map (
            O => \N__42279\,
            I => n10579
        );

    \I__9312\ : InMux
    port map (
            O => \N__42268\,
            I => n19334
        );

    \I__9311\ : CascadeMux
    port map (
            O => \N__42265\,
            I => \n17338_cascade_\
        );

    \I__9310\ : CascadeMux
    port map (
            O => \N__42262\,
            I => \N__42259\
        );

    \I__9309\ : CascadeBuf
    port map (
            O => \N__42259\,
            I => \N__42256\
        );

    \I__9308\ : CascadeMux
    port map (
            O => \N__42256\,
            I => \N__42253\
        );

    \I__9307\ : CascadeBuf
    port map (
            O => \N__42253\,
            I => \N__42250\
        );

    \I__9306\ : CascadeMux
    port map (
            O => \N__42250\,
            I => \N__42247\
        );

    \I__9305\ : CascadeBuf
    port map (
            O => \N__42247\,
            I => \N__42244\
        );

    \I__9304\ : CascadeMux
    port map (
            O => \N__42244\,
            I => \N__42241\
        );

    \I__9303\ : CascadeBuf
    port map (
            O => \N__42241\,
            I => \N__42238\
        );

    \I__9302\ : CascadeMux
    port map (
            O => \N__42238\,
            I => \N__42235\
        );

    \I__9301\ : CascadeBuf
    port map (
            O => \N__42235\,
            I => \N__42232\
        );

    \I__9300\ : CascadeMux
    port map (
            O => \N__42232\,
            I => \N__42229\
        );

    \I__9299\ : CascadeBuf
    port map (
            O => \N__42229\,
            I => \N__42226\
        );

    \I__9298\ : CascadeMux
    port map (
            O => \N__42226\,
            I => \N__42223\
        );

    \I__9297\ : CascadeBuf
    port map (
            O => \N__42223\,
            I => \N__42220\
        );

    \I__9296\ : CascadeMux
    port map (
            O => \N__42220\,
            I => \N__42217\
        );

    \I__9295\ : CascadeBuf
    port map (
            O => \N__42217\,
            I => \N__42213\
        );

    \I__9294\ : CascadeMux
    port map (
            O => \N__42216\,
            I => \N__42210\
        );

    \I__9293\ : CascadeMux
    port map (
            O => \N__42213\,
            I => \N__42207\
        );

    \I__9292\ : CascadeBuf
    port map (
            O => \N__42210\,
            I => \N__42204\
        );

    \I__9291\ : CascadeBuf
    port map (
            O => \N__42207\,
            I => \N__42201\
        );

    \I__9290\ : CascadeMux
    port map (
            O => \N__42204\,
            I => \N__42198\
        );

    \I__9289\ : CascadeMux
    port map (
            O => \N__42201\,
            I => \N__42195\
        );

    \I__9288\ : InMux
    port map (
            O => \N__42198\,
            I => \N__42192\
        );

    \I__9287\ : InMux
    port map (
            O => \N__42195\,
            I => \N__42189\
        );

    \I__9286\ : LocalMux
    port map (
            O => \N__42192\,
            I => \N__42186\
        );

    \I__9285\ : LocalMux
    port map (
            O => \N__42189\,
            I => \N__42183\
        );

    \I__9284\ : Span4Mux_v
    port map (
            O => \N__42186\,
            I => \N__42180\
        );

    \I__9283\ : Span12Mux_s10_v
    port map (
            O => \N__42183\,
            I => \N__42177\
        );

    \I__9282\ : Sp12to4
    port map (
            O => \N__42180\,
            I => \N__42172\
        );

    \I__9281\ : Span12Mux_h
    port map (
            O => \N__42177\,
            I => \N__42172\
        );

    \I__9280\ : Odrv12
    port map (
            O => \N__42172\,
            I => \data_index_9_N_212_5\
        );

    \I__9279\ : InMux
    port map (
            O => \N__42169\,
            I => \N__42166\
        );

    \I__9278\ : LocalMux
    port map (
            O => \N__42166\,
            I => \N__42163\
        );

    \I__9277\ : Odrv4
    port map (
            O => \N__42163\,
            I => n22_adj_1492
        );

    \I__9276\ : CascadeMux
    port map (
            O => \N__42160\,
            I => \n21_adj_1494_cascade_\
        );

    \I__9275\ : InMux
    port map (
            O => \N__42157\,
            I => \N__42154\
        );

    \I__9274\ : LocalMux
    port map (
            O => \N__42154\,
            I => n24_adj_1530
        );

    \I__9273\ : InMux
    port map (
            O => \N__42151\,
            I => \N__42148\
        );

    \I__9272\ : LocalMux
    port map (
            O => \N__42148\,
            I => n30_adj_1597
        );

    \I__9271\ : CascadeMux
    port map (
            O => \N__42145\,
            I => \N__42140\
        );

    \I__9270\ : InMux
    port map (
            O => \N__42144\,
            I => \N__42136\
        );

    \I__9269\ : InMux
    port map (
            O => \N__42143\,
            I => \N__42132\
        );

    \I__9268\ : InMux
    port map (
            O => \N__42140\,
            I => \N__42127\
        );

    \I__9267\ : InMux
    port map (
            O => \N__42139\,
            I => \N__42127\
        );

    \I__9266\ : LocalMux
    port map (
            O => \N__42136\,
            I => \N__42123\
        );

    \I__9265\ : InMux
    port map (
            O => \N__42135\,
            I => \N__42120\
        );

    \I__9264\ : LocalMux
    port map (
            O => \N__42132\,
            I => \N__42116\
        );

    \I__9263\ : LocalMux
    port map (
            O => \N__42127\,
            I => \N__42113\
        );

    \I__9262\ : InMux
    port map (
            O => \N__42126\,
            I => \N__42110\
        );

    \I__9261\ : Span4Mux_h
    port map (
            O => \N__42123\,
            I => \N__42105\
        );

    \I__9260\ : LocalMux
    port map (
            O => \N__42120\,
            I => \N__42105\
        );

    \I__9259\ : InMux
    port map (
            O => \N__42119\,
            I => \N__42102\
        );

    \I__9258\ : Span4Mux_v
    port map (
            O => \N__42116\,
            I => \N__42095\
        );

    \I__9257\ : Span4Mux_v
    port map (
            O => \N__42113\,
            I => \N__42095\
        );

    \I__9256\ : LocalMux
    port map (
            O => \N__42110\,
            I => \N__42095\
        );

    \I__9255\ : Span4Mux_h
    port map (
            O => \N__42105\,
            I => \N__42090\
        );

    \I__9254\ : LocalMux
    port map (
            O => \N__42102\,
            I => \N__42090\
        );

    \I__9253\ : Span4Mux_h
    port map (
            O => \N__42095\,
            I => \N__42087\
        );

    \I__9252\ : Span4Mux_v
    port map (
            O => \N__42090\,
            I => \N__42084\
        );

    \I__9251\ : Span4Mux_v
    port map (
            O => \N__42087\,
            I => \N__42081\
        );

    \I__9250\ : Odrv4
    port map (
            O => \N__42084\,
            I => n14_adj_1549
        );

    \I__9249\ : Odrv4
    port map (
            O => \N__42081\,
            I => n14_adj_1549
        );

    \I__9248\ : CascadeMux
    port map (
            O => \N__42076\,
            I => \N__42071\
        );

    \I__9247\ : CascadeMux
    port map (
            O => \N__42075\,
            I => \N__42068\
        );

    \I__9246\ : CascadeMux
    port map (
            O => \N__42074\,
            I => \N__42065\
        );

    \I__9245\ : InMux
    port map (
            O => \N__42071\,
            I => \N__42062\
        );

    \I__9244\ : InMux
    port map (
            O => \N__42068\,
            I => \N__42057\
        );

    \I__9243\ : InMux
    port map (
            O => \N__42065\,
            I => \N__42057\
        );

    \I__9242\ : LocalMux
    port map (
            O => \N__42062\,
            I => \N__42054\
        );

    \I__9241\ : LocalMux
    port map (
            O => \N__42057\,
            I => \N__42051\
        );

    \I__9240\ : Span4Mux_v
    port map (
            O => \N__42054\,
            I => \N__42046\
        );

    \I__9239\ : Span4Mux_h
    port map (
            O => \N__42051\,
            I => \N__42046\
        );

    \I__9238\ : Span4Mux_v
    port map (
            O => \N__42046\,
            I => \N__42041\
        );

    \I__9237\ : InMux
    port map (
            O => \N__42045\,
            I => \N__42038\
        );

    \I__9236\ : InMux
    port map (
            O => \N__42044\,
            I => \N__42035\
        );

    \I__9235\ : Sp12to4
    port map (
            O => \N__42041\,
            I => \N__42030\
        );

    \I__9234\ : LocalMux
    port map (
            O => \N__42038\,
            I => \N__42030\
        );

    \I__9233\ : LocalMux
    port map (
            O => \N__42035\,
            I => \buf_cfgRTD_4\
        );

    \I__9232\ : Odrv12
    port map (
            O => \N__42030\,
            I => \buf_cfgRTD_4\
        );

    \I__9231\ : CascadeMux
    port map (
            O => \N__42025\,
            I => \N__42021\
        );

    \I__9230\ : InMux
    port map (
            O => \N__42024\,
            I => \N__42016\
        );

    \I__9229\ : InMux
    port map (
            O => \N__42021\,
            I => \N__42009\
        );

    \I__9228\ : InMux
    port map (
            O => \N__42020\,
            I => \N__42009\
        );

    \I__9227\ : InMux
    port map (
            O => \N__42019\,
            I => \N__42009\
        );

    \I__9226\ : LocalMux
    port map (
            O => \N__42016\,
            I => \N__42001\
        );

    \I__9225\ : LocalMux
    port map (
            O => \N__42009\,
            I => \N__41998\
        );

    \I__9224\ : InMux
    port map (
            O => \N__42008\,
            I => \N__41993\
        );

    \I__9223\ : InMux
    port map (
            O => \N__42007\,
            I => \N__41993\
        );

    \I__9222\ : InMux
    port map (
            O => \N__42006\,
            I => \N__41980\
        );

    \I__9221\ : InMux
    port map (
            O => \N__42005\,
            I => \N__41980\
        );

    \I__9220\ : InMux
    port map (
            O => \N__42004\,
            I => \N__41980\
        );

    \I__9219\ : Span4Mux_v
    port map (
            O => \N__42001\,
            I => \N__41973\
        );

    \I__9218\ : Span4Mux_h
    port map (
            O => \N__41998\,
            I => \N__41973\
        );

    \I__9217\ : LocalMux
    port map (
            O => \N__41993\,
            I => \N__41973\
        );

    \I__9216\ : InMux
    port map (
            O => \N__41992\,
            I => \N__41968\
        );

    \I__9215\ : InMux
    port map (
            O => \N__41991\,
            I => \N__41968\
        );

    \I__9214\ : InMux
    port map (
            O => \N__41990\,
            I => \N__41959\
        );

    \I__9213\ : InMux
    port map (
            O => \N__41989\,
            I => \N__41959\
        );

    \I__9212\ : InMux
    port map (
            O => \N__41988\,
            I => \N__41959\
        );

    \I__9211\ : InMux
    port map (
            O => \N__41987\,
            I => \N__41959\
        );

    \I__9210\ : LocalMux
    port map (
            O => \N__41980\,
            I => n12415
        );

    \I__9209\ : Odrv4
    port map (
            O => \N__41973\,
            I => n12415
        );

    \I__9208\ : LocalMux
    port map (
            O => \N__41968\,
            I => n12415
        );

    \I__9207\ : LocalMux
    port map (
            O => \N__41959\,
            I => n12415
        );

    \I__9206\ : InMux
    port map (
            O => \N__41950\,
            I => \N__41947\
        );

    \I__9205\ : LocalMux
    port map (
            O => \N__41947\,
            I => \N__41944\
        );

    \I__9204\ : Span4Mux_v
    port map (
            O => \N__41944\,
            I => \N__41940\
        );

    \I__9203\ : InMux
    port map (
            O => \N__41943\,
            I => \N__41937\
        );

    \I__9202\ : Span4Mux_h
    port map (
            O => \N__41940\,
            I => \N__41932\
        );

    \I__9201\ : LocalMux
    port map (
            O => \N__41937\,
            I => \N__41932\
        );

    \I__9200\ : Span4Mux_h
    port map (
            O => \N__41932\,
            I => \N__41929\
        );

    \I__9199\ : Odrv4
    port map (
            O => \N__41929\,
            I => n14_adj_1551
        );

    \I__9198\ : CascadeMux
    port map (
            O => \N__41926\,
            I => \N__41923\
        );

    \I__9197\ : InMux
    port map (
            O => \N__41923\,
            I => \N__41920\
        );

    \I__9196\ : LocalMux
    port map (
            O => \N__41920\,
            I => \N__41917\
        );

    \I__9195\ : Span4Mux_v
    port map (
            O => \N__41917\,
            I => \N__41914\
        );

    \I__9194\ : Span4Mux_h
    port map (
            O => \N__41914\,
            I => \N__41909\
        );

    \I__9193\ : InMux
    port map (
            O => \N__41913\,
            I => \N__41904\
        );

    \I__9192\ : InMux
    port map (
            O => \N__41912\,
            I => \N__41904\
        );

    \I__9191\ : Odrv4
    port map (
            O => \N__41909\,
            I => req_data_cnt_10
        );

    \I__9190\ : LocalMux
    port map (
            O => \N__41904\,
            I => req_data_cnt_10
        );

    \I__9189\ : InMux
    port map (
            O => \N__41899\,
            I => \N__41896\
        );

    \I__9188\ : LocalMux
    port map (
            O => \N__41896\,
            I => \N__41892\
        );

    \I__9187\ : InMux
    port map (
            O => \N__41895\,
            I => \N__41888\
        );

    \I__9186\ : Span12Mux_h
    port map (
            O => \N__41892\,
            I => \N__41885\
        );

    \I__9185\ : InMux
    port map (
            O => \N__41891\,
            I => \N__41882\
        );

    \I__9184\ : LocalMux
    port map (
            O => \N__41888\,
            I => req_data_cnt_8
        );

    \I__9183\ : Odrv12
    port map (
            O => \N__41885\,
            I => req_data_cnt_8
        );

    \I__9182\ : LocalMux
    port map (
            O => \N__41882\,
            I => req_data_cnt_8
        );

    \I__9181\ : InMux
    port map (
            O => \N__41875\,
            I => \N__41872\
        );

    \I__9180\ : LocalMux
    port map (
            O => \N__41872\,
            I => n19_adj_1499
        );

    \I__9179\ : InMux
    port map (
            O => \N__41869\,
            I => \bfn_16_15_0_\
        );

    \I__9178\ : InMux
    port map (
            O => \N__41866\,
            I => n19326
        );

    \I__9177\ : InMux
    port map (
            O => \N__41863\,
            I => \N__41858\
        );

    \I__9176\ : InMux
    port map (
            O => \N__41862\,
            I => \N__41855\
        );

    \I__9175\ : InMux
    port map (
            O => \N__41861\,
            I => \N__41852\
        );

    \I__9174\ : LocalMux
    port map (
            O => \N__41858\,
            I => \N__41847\
        );

    \I__9173\ : LocalMux
    port map (
            O => \N__41855\,
            I => \N__41847\
        );

    \I__9172\ : LocalMux
    port map (
            O => \N__41852\,
            I => data_index_2
        );

    \I__9171\ : Odrv12
    port map (
            O => \N__41847\,
            I => data_index_2
        );

    \I__9170\ : InMux
    port map (
            O => \N__41842\,
            I => \N__41836\
        );

    \I__9169\ : InMux
    port map (
            O => \N__41841\,
            I => \N__41836\
        );

    \I__9168\ : LocalMux
    port map (
            O => \N__41836\,
            I => \N__41833\
        );

    \I__9167\ : Odrv4
    port map (
            O => \N__41833\,
            I => n7_adj_1544
        );

    \I__9166\ : InMux
    port map (
            O => \N__41830\,
            I => n19327
        );

    \I__9165\ : InMux
    port map (
            O => \N__41827\,
            I => \N__41822\
        );

    \I__9164\ : InMux
    port map (
            O => \N__41826\,
            I => \N__41819\
        );

    \I__9163\ : InMux
    port map (
            O => \N__41825\,
            I => \N__41816\
        );

    \I__9162\ : LocalMux
    port map (
            O => \N__41822\,
            I => \N__41813\
        );

    \I__9161\ : LocalMux
    port map (
            O => \N__41819\,
            I => \N__41808\
        );

    \I__9160\ : LocalMux
    port map (
            O => \N__41816\,
            I => \N__41808\
        );

    \I__9159\ : Span4Mux_v
    port map (
            O => \N__41813\,
            I => \N__41805\
        );

    \I__9158\ : Span4Mux_h
    port map (
            O => \N__41808\,
            I => \N__41802\
        );

    \I__9157\ : Odrv4
    port map (
            O => \N__41805\,
            I => data_index_3
        );

    \I__9156\ : Odrv4
    port map (
            O => \N__41802\,
            I => data_index_3
        );

    \I__9155\ : InMux
    port map (
            O => \N__41797\,
            I => \N__41791\
        );

    \I__9154\ : InMux
    port map (
            O => \N__41796\,
            I => \N__41791\
        );

    \I__9153\ : LocalMux
    port map (
            O => \N__41791\,
            I => \N__41788\
        );

    \I__9152\ : Odrv12
    port map (
            O => \N__41788\,
            I => n7_adj_1542
        );

    \I__9151\ : InMux
    port map (
            O => \N__41785\,
            I => n19328
        );

    \I__9150\ : InMux
    port map (
            O => \N__41782\,
            I => \N__41778\
        );

    \I__9149\ : InMux
    port map (
            O => \N__41781\,
            I => \N__41775\
        );

    \I__9148\ : LocalMux
    port map (
            O => \N__41778\,
            I => \N__41772\
        );

    \I__9147\ : LocalMux
    port map (
            O => \N__41775\,
            I => \N__41769\
        );

    \I__9146\ : Span4Mux_v
    port map (
            O => \N__41772\,
            I => \N__41766\
        );

    \I__9145\ : Span4Mux_v
    port map (
            O => \N__41769\,
            I => \N__41763\
        );

    \I__9144\ : Span4Mux_h
    port map (
            O => \N__41766\,
            I => \N__41760\
        );

    \I__9143\ : Span4Mux_v
    port map (
            O => \N__41763\,
            I => \N__41757\
        );

    \I__9142\ : Odrv4
    port map (
            O => \N__41760\,
            I => n14_adj_1524
        );

    \I__9141\ : Odrv4
    port map (
            O => \N__41757\,
            I => n14_adj_1524
        );

    \I__9140\ : InMux
    port map (
            O => \N__41752\,
            I => \N__41748\
        );

    \I__9139\ : CascadeMux
    port map (
            O => \N__41751\,
            I => \N__41745\
        );

    \I__9138\ : LocalMux
    port map (
            O => \N__41748\,
            I => \N__41741\
        );

    \I__9137\ : InMux
    port map (
            O => \N__41745\,
            I => \N__41738\
        );

    \I__9136\ : InMux
    port map (
            O => \N__41744\,
            I => \N__41735\
        );

    \I__9135\ : Span4Mux_v
    port map (
            O => \N__41741\,
            I => \N__41732\
        );

    \I__9134\ : LocalMux
    port map (
            O => \N__41738\,
            I => \N__41729\
        );

    \I__9133\ : LocalMux
    port map (
            O => \N__41735\,
            I => req_data_cnt_0
        );

    \I__9132\ : Odrv4
    port map (
            O => \N__41732\,
            I => req_data_cnt_0
        );

    \I__9131\ : Odrv4
    port map (
            O => \N__41729\,
            I => req_data_cnt_0
        );

    \I__9130\ : InMux
    port map (
            O => \N__41722\,
            I => \N__41719\
        );

    \I__9129\ : LocalMux
    port map (
            O => \N__41719\,
            I => \N__41715\
        );

    \I__9128\ : InMux
    port map (
            O => \N__41718\,
            I => \N__41711\
        );

    \I__9127\ : Span12Mux_v
    port map (
            O => \N__41715\,
            I => \N__41708\
        );

    \I__9126\ : InMux
    port map (
            O => \N__41714\,
            I => \N__41705\
        );

    \I__9125\ : LocalMux
    port map (
            O => \N__41711\,
            I => req_data_cnt_6
        );

    \I__9124\ : Odrv12
    port map (
            O => \N__41708\,
            I => req_data_cnt_6
        );

    \I__9123\ : LocalMux
    port map (
            O => \N__41705\,
            I => req_data_cnt_6
        );

    \I__9122\ : InMux
    port map (
            O => \N__41698\,
            I => \N__41695\
        );

    \I__9121\ : LocalMux
    port map (
            O => \N__41695\,
            I => n17_adj_1554
        );

    \I__9120\ : InMux
    port map (
            O => \N__41692\,
            I => \N__41688\
        );

    \I__9119\ : CascadeMux
    port map (
            O => \N__41691\,
            I => \N__41685\
        );

    \I__9118\ : LocalMux
    port map (
            O => \N__41688\,
            I => \N__41681\
        );

    \I__9117\ : InMux
    port map (
            O => \N__41685\,
            I => \N__41678\
        );

    \I__9116\ : InMux
    port map (
            O => \N__41684\,
            I => \N__41675\
        );

    \I__9115\ : Span4Mux_h
    port map (
            O => \N__41681\,
            I => \N__41672\
        );

    \I__9114\ : LocalMux
    port map (
            O => \N__41678\,
            I => \N__41669\
        );

    \I__9113\ : LocalMux
    port map (
            O => \N__41675\,
            I => \N__41664\
        );

    \I__9112\ : Span4Mux_v
    port map (
            O => \N__41672\,
            I => \N__41664\
        );

    \I__9111\ : Span4Mux_v
    port map (
            O => \N__41669\,
            I => \N__41661\
        );

    \I__9110\ : Odrv4
    port map (
            O => \N__41664\,
            I => req_data_cnt_15
        );

    \I__9109\ : Odrv4
    port map (
            O => \N__41661\,
            I => req_data_cnt_15
        );

    \I__9108\ : CascadeMux
    port map (
            O => \N__41656\,
            I => \N__41653\
        );

    \I__9107\ : InMux
    port map (
            O => \N__41653\,
            I => \N__41650\
        );

    \I__9106\ : LocalMux
    port map (
            O => \N__41650\,
            I => \N__41647\
        );

    \I__9105\ : Span4Mux_h
    port map (
            O => \N__41647\,
            I => \N__41643\
        );

    \I__9104\ : InMux
    port map (
            O => \N__41646\,
            I => \N__41639\
        );

    \I__9103\ : Span4Mux_h
    port map (
            O => \N__41643\,
            I => \N__41636\
        );

    \I__9102\ : InMux
    port map (
            O => \N__41642\,
            I => \N__41633\
        );

    \I__9101\ : LocalMux
    port map (
            O => \N__41639\,
            I => req_data_cnt_9
        );

    \I__9100\ : Odrv4
    port map (
            O => \N__41636\,
            I => req_data_cnt_9
        );

    \I__9099\ : LocalMux
    port map (
            O => \N__41633\,
            I => req_data_cnt_9
        );

    \I__9098\ : InMux
    port map (
            O => \N__41626\,
            I => \N__41623\
        );

    \I__9097\ : LocalMux
    port map (
            O => \N__41623\,
            I => \N__41619\
        );

    \I__9096\ : InMux
    port map (
            O => \N__41622\,
            I => \N__41616\
        );

    \I__9095\ : Span4Mux_v
    port map (
            O => \N__41619\,
            I => \N__41609\
        );

    \I__9094\ : LocalMux
    port map (
            O => \N__41616\,
            I => \N__41609\
        );

    \I__9093\ : InMux
    port map (
            O => \N__41615\,
            I => \N__41606\
        );

    \I__9092\ : InMux
    port map (
            O => \N__41614\,
            I => \N__41603\
        );

    \I__9091\ : Odrv4
    port map (
            O => \N__41609\,
            I => n20613
        );

    \I__9090\ : LocalMux
    port map (
            O => \N__41606\,
            I => n20613
        );

    \I__9089\ : LocalMux
    port map (
            O => \N__41603\,
            I => n20613
        );

    \I__9088\ : InMux
    port map (
            O => \N__41596\,
            I => \N__41593\
        );

    \I__9087\ : LocalMux
    port map (
            O => \N__41593\,
            I => \N__41588\
        );

    \I__9086\ : CascadeMux
    port map (
            O => \N__41592\,
            I => \N__41585\
        );

    \I__9085\ : InMux
    port map (
            O => \N__41591\,
            I => \N__41582\
        );

    \I__9084\ : Span4Mux_v
    port map (
            O => \N__41588\,
            I => \N__41579\
        );

    \I__9083\ : InMux
    port map (
            O => \N__41585\,
            I => \N__41576\
        );

    \I__9082\ : LocalMux
    port map (
            O => \N__41582\,
            I => req_data_cnt_2
        );

    \I__9081\ : Odrv4
    port map (
            O => \N__41579\,
            I => req_data_cnt_2
        );

    \I__9080\ : LocalMux
    port map (
            O => \N__41576\,
            I => req_data_cnt_2
        );

    \I__9079\ : InMux
    port map (
            O => \N__41569\,
            I => \N__41566\
        );

    \I__9078\ : LocalMux
    port map (
            O => \N__41566\,
            I => \N__41562\
        );

    \I__9077\ : InMux
    port map (
            O => \N__41565\,
            I => \N__41558\
        );

    \I__9076\ : Span12Mux_v
    port map (
            O => \N__41562\,
            I => \N__41555\
        );

    \I__9075\ : InMux
    port map (
            O => \N__41561\,
            I => \N__41552\
        );

    \I__9074\ : LocalMux
    port map (
            O => \N__41558\,
            I => req_data_cnt_7
        );

    \I__9073\ : Odrv12
    port map (
            O => \N__41555\,
            I => req_data_cnt_7
        );

    \I__9072\ : LocalMux
    port map (
            O => \N__41552\,
            I => req_data_cnt_7
        );

    \I__9071\ : CascadeMux
    port map (
            O => \N__41545\,
            I => \N__41541\
        );

    \I__9070\ : InMux
    port map (
            O => \N__41544\,
            I => \N__41536\
        );

    \I__9069\ : InMux
    port map (
            O => \N__41541\,
            I => \N__41536\
        );

    \I__9068\ : LocalMux
    port map (
            O => \N__41536\,
            I => \N__41532\
        );

    \I__9067\ : CascadeMux
    port map (
            O => \N__41535\,
            I => \N__41529\
        );

    \I__9066\ : Span4Mux_v
    port map (
            O => \N__41532\,
            I => \N__41523\
        );

    \I__9065\ : InMux
    port map (
            O => \N__41529\,
            I => \N__41518\
        );

    \I__9064\ : InMux
    port map (
            O => \N__41528\,
            I => \N__41518\
        );

    \I__9063\ : InMux
    port map (
            O => \N__41527\,
            I => \N__41515\
        );

    \I__9062\ : InMux
    port map (
            O => \N__41526\,
            I => \N__41512\
        );

    \I__9061\ : Span4Mux_h
    port map (
            O => \N__41523\,
            I => \N__41507\
        );

    \I__9060\ : LocalMux
    port map (
            O => \N__41518\,
            I => \N__41507\
        );

    \I__9059\ : LocalMux
    port map (
            O => \N__41515\,
            I => \N__41503\
        );

    \I__9058\ : LocalMux
    port map (
            O => \N__41512\,
            I => \N__41500\
        );

    \I__9057\ : Span4Mux_v
    port map (
            O => \N__41507\,
            I => \N__41497\
        );

    \I__9056\ : InMux
    port map (
            O => \N__41506\,
            I => \N__41494\
        );

    \I__9055\ : Span4Mux_v
    port map (
            O => \N__41503\,
            I => \N__41491\
        );

    \I__9054\ : Span4Mux_h
    port map (
            O => \N__41500\,
            I => \N__41488\
        );

    \I__9053\ : Span4Mux_v
    port map (
            O => \N__41497\,
            I => \N__41485\
        );

    \I__9052\ : LocalMux
    port map (
            O => \N__41494\,
            I => \N__41482\
        );

    \I__9051\ : Span4Mux_h
    port map (
            O => \N__41491\,
            I => \N__41477\
        );

    \I__9050\ : Span4Mux_v
    port map (
            O => \N__41488\,
            I => \N__41477\
        );

    \I__9049\ : Odrv4
    port map (
            O => \N__41485\,
            I => n14_adj_1548
        );

    \I__9048\ : Odrv12
    port map (
            O => \N__41482\,
            I => n14_adj_1548
        );

    \I__9047\ : Odrv4
    port map (
            O => \N__41477\,
            I => n14_adj_1548
        );

    \I__9046\ : CascadeMux
    port map (
            O => \N__41470\,
            I => \N__41466\
        );

    \I__9045\ : InMux
    port map (
            O => \N__41469\,
            I => \N__41463\
        );

    \I__9044\ : InMux
    port map (
            O => \N__41466\,
            I => \N__41460\
        );

    \I__9043\ : LocalMux
    port map (
            O => \N__41463\,
            I => \N__41457\
        );

    \I__9042\ : LocalMux
    port map (
            O => \N__41460\,
            I => \N__41452\
        );

    \I__9041\ : Span4Mux_h
    port map (
            O => \N__41457\,
            I => \N__41452\
        );

    \I__9040\ : Odrv4
    port map (
            O => \N__41452\,
            I => data_idxvec_8
        );

    \I__9039\ : InMux
    port map (
            O => \N__41449\,
            I => \N__41446\
        );

    \I__9038\ : LocalMux
    port map (
            O => \N__41446\,
            I => \N__41443\
        );

    \I__9037\ : Odrv12
    port map (
            O => \N__41443\,
            I => n20779
        );

    \I__9036\ : CascadeMux
    port map (
            O => \N__41440\,
            I => \n12415_cascade_\
        );

    \I__9035\ : CascadeMux
    port map (
            O => \N__41437\,
            I => \N__41433\
        );

    \I__9034\ : CascadeMux
    port map (
            O => \N__41436\,
            I => \N__41430\
        );

    \I__9033\ : InMux
    port map (
            O => \N__41433\,
            I => \N__41427\
        );

    \I__9032\ : InMux
    port map (
            O => \N__41430\,
            I => \N__41422\
        );

    \I__9031\ : LocalMux
    port map (
            O => \N__41427\,
            I => \N__41419\
        );

    \I__9030\ : InMux
    port map (
            O => \N__41426\,
            I => \N__41416\
        );

    \I__9029\ : InMux
    port map (
            O => \N__41425\,
            I => \N__41413\
        );

    \I__9028\ : LocalMux
    port map (
            O => \N__41422\,
            I => \N__41410\
        );

    \I__9027\ : Span4Mux_v
    port map (
            O => \N__41419\,
            I => \N__41405\
        );

    \I__9026\ : LocalMux
    port map (
            O => \N__41416\,
            I => \N__41405\
        );

    \I__9025\ : LocalMux
    port map (
            O => \N__41413\,
            I => \N__41402\
        );

    \I__9024\ : Span4Mux_v
    port map (
            O => \N__41410\,
            I => \N__41399\
        );

    \I__9023\ : Span4Mux_v
    port map (
            O => \N__41405\,
            I => \N__41396\
        );

    \I__9022\ : Span4Mux_h
    port map (
            O => \N__41402\,
            I => \N__41393\
        );

    \I__9021\ : Span4Mux_h
    port map (
            O => \N__41399\,
            I => \N__41390\
        );

    \I__9020\ : Span4Mux_h
    port map (
            O => \N__41396\,
            I => \N__41387\
        );

    \I__9019\ : Span4Mux_h
    port map (
            O => \N__41393\,
            I => \N__41383\
        );

    \I__9018\ : Sp12to4
    port map (
            O => \N__41390\,
            I => \N__41378\
        );

    \I__9017\ : Sp12to4
    port map (
            O => \N__41387\,
            I => \N__41378\
        );

    \I__9016\ : InMux
    port map (
            O => \N__41386\,
            I => \N__41375\
        );

    \I__9015\ : Span4Mux_h
    port map (
            O => \N__41383\,
            I => \N__41372\
        );

    \I__9014\ : Odrv12
    port map (
            O => \N__41378\,
            I => \buf_cfgRTD_5\
        );

    \I__9013\ : LocalMux
    port map (
            O => \N__41375\,
            I => \buf_cfgRTD_5\
        );

    \I__9012\ : Odrv4
    port map (
            O => \N__41372\,
            I => \buf_cfgRTD_5\
        );

    \I__9011\ : InMux
    port map (
            O => \N__41365\,
            I => \N__41360\
        );

    \I__9010\ : CascadeMux
    port map (
            O => \N__41364\,
            I => \N__41357\
        );

    \I__9009\ : CascadeMux
    port map (
            O => \N__41363\,
            I => \N__41351\
        );

    \I__9008\ : LocalMux
    port map (
            O => \N__41360\,
            I => \N__41348\
        );

    \I__9007\ : InMux
    port map (
            O => \N__41357\,
            I => \N__41342\
        );

    \I__9006\ : InMux
    port map (
            O => \N__41356\,
            I => \N__41342\
        );

    \I__9005\ : InMux
    port map (
            O => \N__41355\,
            I => \N__41339\
        );

    \I__9004\ : InMux
    port map (
            O => \N__41354\,
            I => \N__41336\
        );

    \I__9003\ : InMux
    port map (
            O => \N__41351\,
            I => \N__41333\
        );

    \I__9002\ : Span4Mux_h
    port map (
            O => \N__41348\,
            I => \N__41330\
        );

    \I__9001\ : InMux
    port map (
            O => \N__41347\,
            I => \N__41327\
        );

    \I__9000\ : LocalMux
    port map (
            O => \N__41342\,
            I => \N__41324\
        );

    \I__8999\ : LocalMux
    port map (
            O => \N__41339\,
            I => \N__41321\
        );

    \I__8998\ : LocalMux
    port map (
            O => \N__41336\,
            I => \N__41318\
        );

    \I__8997\ : LocalMux
    port map (
            O => \N__41333\,
            I => \N__41315\
        );

    \I__8996\ : Span4Mux_v
    port map (
            O => \N__41330\,
            I => \N__41312\
        );

    \I__8995\ : LocalMux
    port map (
            O => \N__41327\,
            I => \N__41309\
        );

    \I__8994\ : Span4Mux_h
    port map (
            O => \N__41324\,
            I => \N__41306\
        );

    \I__8993\ : Span12Mux_v
    port map (
            O => \N__41321\,
            I => \N__41303\
        );

    \I__8992\ : Span4Mux_v
    port map (
            O => \N__41318\,
            I => \N__41300\
        );

    \I__8991\ : Span4Mux_v
    port map (
            O => \N__41315\,
            I => \N__41293\
        );

    \I__8990\ : Span4Mux_h
    port map (
            O => \N__41312\,
            I => \N__41293\
        );

    \I__8989\ : Span4Mux_v
    port map (
            O => \N__41309\,
            I => \N__41293\
        );

    \I__8988\ : Odrv4
    port map (
            O => \N__41306\,
            I => comm_buf_1_0
        );

    \I__8987\ : Odrv12
    port map (
            O => \N__41303\,
            I => comm_buf_1_0
        );

    \I__8986\ : Odrv4
    port map (
            O => \N__41300\,
            I => comm_buf_1_0
        );

    \I__8985\ : Odrv4
    port map (
            O => \N__41293\,
            I => comm_buf_1_0
        );

    \I__8984\ : InMux
    port map (
            O => \N__41284\,
            I => \N__41280\
        );

    \I__8983\ : InMux
    port map (
            O => \N__41283\,
            I => \N__41277\
        );

    \I__8982\ : LocalMux
    port map (
            O => \N__41280\,
            I => \N__41274\
        );

    \I__8981\ : LocalMux
    port map (
            O => \N__41277\,
            I => \N__41269\
        );

    \I__8980\ : Span4Mux_h
    port map (
            O => \N__41274\,
            I => \N__41269\
        );

    \I__8979\ : Span4Mux_h
    port map (
            O => \N__41269\,
            I => \N__41266\
        );

    \I__8978\ : Odrv4
    port map (
            O => \N__41266\,
            I => n14_adj_1528
        );

    \I__8977\ : InMux
    port map (
            O => \N__41263\,
            I => \N__41260\
        );

    \I__8976\ : LocalMux
    port map (
            O => \N__41260\,
            I => \N__41256\
        );

    \I__8975\ : InMux
    port map (
            O => \N__41259\,
            I => \N__41253\
        );

    \I__8974\ : Span4Mux_h
    port map (
            O => \N__41256\,
            I => \N__41248\
        );

    \I__8973\ : LocalMux
    port map (
            O => \N__41253\,
            I => \N__41248\
        );

    \I__8972\ : Span4Mux_h
    port map (
            O => \N__41248\,
            I => \N__41245\
        );

    \I__8971\ : Odrv4
    port map (
            O => \N__41245\,
            I => n14_adj_1525
        );

    \I__8970\ : InMux
    port map (
            O => \N__41242\,
            I => \N__41239\
        );

    \I__8969\ : LocalMux
    port map (
            O => \N__41239\,
            I => \N__41236\
        );

    \I__8968\ : Span12Mux_v
    port map (
            O => \N__41236\,
            I => \N__41233\
        );

    \I__8967\ : Odrv12
    port map (
            O => \N__41233\,
            I => n20850
        );

    \I__8966\ : InMux
    port map (
            O => \N__41230\,
            I => \N__41227\
        );

    \I__8965\ : LocalMux
    port map (
            O => \N__41227\,
            I => \N__41224\
        );

    \I__8964\ : Span4Mux_h
    port map (
            O => \N__41224\,
            I => \N__41221\
        );

    \I__8963\ : Span4Mux_h
    port map (
            O => \N__41221\,
            I => \N__41218\
        );

    \I__8962\ : Odrv4
    port map (
            O => \N__41218\,
            I => n30_adj_1520
        );

    \I__8961\ : InMux
    port map (
            O => \N__41215\,
            I => \N__41212\
        );

    \I__8960\ : LocalMux
    port map (
            O => \N__41212\,
            I => \N__41209\
        );

    \I__8959\ : Span4Mux_v
    port map (
            O => \N__41209\,
            I => \N__41206\
        );

    \I__8958\ : Odrv4
    port map (
            O => \N__41206\,
            I => n22_adj_1594
        );

    \I__8957\ : InMux
    port map (
            O => \N__41203\,
            I => \N__41200\
        );

    \I__8956\ : LocalMux
    port map (
            O => \N__41200\,
            I => n10_adj_1582
        );

    \I__8955\ : CascadeMux
    port map (
            O => \N__41197\,
            I => \N__41193\
        );

    \I__8954\ : InMux
    port map (
            O => \N__41196\,
            I => \N__41190\
        );

    \I__8953\ : InMux
    port map (
            O => \N__41193\,
            I => \N__41186\
        );

    \I__8952\ : LocalMux
    port map (
            O => \N__41190\,
            I => \N__41183\
        );

    \I__8951\ : InMux
    port map (
            O => \N__41189\,
            I => \N__41180\
        );

    \I__8950\ : LocalMux
    port map (
            O => \N__41186\,
            I => \N__41177\
        );

    \I__8949\ : Odrv12
    port map (
            O => \N__41183\,
            I => clk_cnt_1
        );

    \I__8948\ : LocalMux
    port map (
            O => \N__41180\,
            I => clk_cnt_1
        );

    \I__8947\ : Odrv4
    port map (
            O => \N__41177\,
            I => clk_cnt_1
        );

    \I__8946\ : InMux
    port map (
            O => \N__41170\,
            I => \N__41166\
        );

    \I__8945\ : InMux
    port map (
            O => \N__41169\,
            I => \N__41161\
        );

    \I__8944\ : LocalMux
    port map (
            O => \N__41166\,
            I => \N__41158\
        );

    \I__8943\ : InMux
    port map (
            O => \N__41165\,
            I => \N__41153\
        );

    \I__8942\ : InMux
    port map (
            O => \N__41164\,
            I => \N__41153\
        );

    \I__8941\ : LocalMux
    port map (
            O => \N__41161\,
            I => \N__41150\
        );

    \I__8940\ : Odrv12
    port map (
            O => \N__41158\,
            I => clk_cnt_0
        );

    \I__8939\ : LocalMux
    port map (
            O => \N__41153\,
            I => clk_cnt_0
        );

    \I__8938\ : Odrv4
    port map (
            O => \N__41150\,
            I => clk_cnt_0
        );

    \I__8937\ : ClkMux
    port map (
            O => \N__41143\,
            I => \N__41138\
        );

    \I__8936\ : ClkMux
    port map (
            O => \N__41142\,
            I => \N__41135\
        );

    \I__8935\ : ClkMux
    port map (
            O => \N__41141\,
            I => \N__41126\
        );

    \I__8934\ : LocalMux
    port map (
            O => \N__41138\,
            I => \N__41123\
        );

    \I__8933\ : LocalMux
    port map (
            O => \N__41135\,
            I => \N__41120\
        );

    \I__8932\ : ClkMux
    port map (
            O => \N__41134\,
            I => \N__41117\
        );

    \I__8931\ : ClkMux
    port map (
            O => \N__41133\,
            I => \N__41112\
        );

    \I__8930\ : ClkMux
    port map (
            O => \N__41132\,
            I => \N__41109\
        );

    \I__8929\ : ClkMux
    port map (
            O => \N__41131\,
            I => \N__41106\
        );

    \I__8928\ : ClkMux
    port map (
            O => \N__41130\,
            I => \N__41103\
        );

    \I__8927\ : ClkMux
    port map (
            O => \N__41129\,
            I => \N__41100\
        );

    \I__8926\ : LocalMux
    port map (
            O => \N__41126\,
            I => \N__41094\
        );

    \I__8925\ : Span4Mux_h
    port map (
            O => \N__41123\,
            I => \N__41087\
        );

    \I__8924\ : Span4Mux_v
    port map (
            O => \N__41120\,
            I => \N__41087\
        );

    \I__8923\ : LocalMux
    port map (
            O => \N__41117\,
            I => \N__41087\
        );

    \I__8922\ : ClkMux
    port map (
            O => \N__41116\,
            I => \N__41084\
        );

    \I__8921\ : ClkMux
    port map (
            O => \N__41115\,
            I => \N__41076\
        );

    \I__8920\ : LocalMux
    port map (
            O => \N__41112\,
            I => \N__41073\
        );

    \I__8919\ : LocalMux
    port map (
            O => \N__41109\,
            I => \N__41070\
        );

    \I__8918\ : LocalMux
    port map (
            O => \N__41106\,
            I => \N__41067\
        );

    \I__8917\ : LocalMux
    port map (
            O => \N__41103\,
            I => \N__41062\
        );

    \I__8916\ : LocalMux
    port map (
            O => \N__41100\,
            I => \N__41062\
        );

    \I__8915\ : ClkMux
    port map (
            O => \N__41099\,
            I => \N__41059\
        );

    \I__8914\ : ClkMux
    port map (
            O => \N__41098\,
            I => \N__41056\
        );

    \I__8913\ : ClkMux
    port map (
            O => \N__41097\,
            I => \N__41053\
        );

    \I__8912\ : Span4Mux_h
    port map (
            O => \N__41094\,
            I => \N__41046\
        );

    \I__8911\ : Span4Mux_h
    port map (
            O => \N__41087\,
            I => \N__41046\
        );

    \I__8910\ : LocalMux
    port map (
            O => \N__41084\,
            I => \N__41046\
        );

    \I__8909\ : ClkMux
    port map (
            O => \N__41083\,
            I => \N__41043\
        );

    \I__8908\ : ClkMux
    port map (
            O => \N__41082\,
            I => \N__41040\
        );

    \I__8907\ : ClkMux
    port map (
            O => \N__41081\,
            I => \N__41037\
        );

    \I__8906\ : ClkMux
    port map (
            O => \N__41080\,
            I => \N__41034\
        );

    \I__8905\ : ClkMux
    port map (
            O => \N__41079\,
            I => \N__41031\
        );

    \I__8904\ : LocalMux
    port map (
            O => \N__41076\,
            I => \N__41026\
        );

    \I__8903\ : Span4Mux_v
    port map (
            O => \N__41073\,
            I => \N__41026\
        );

    \I__8902\ : Span4Mux_v
    port map (
            O => \N__41070\,
            I => \N__41017\
        );

    \I__8901\ : Span4Mux_h
    port map (
            O => \N__41067\,
            I => \N__41017\
        );

    \I__8900\ : Span4Mux_v
    port map (
            O => \N__41062\,
            I => \N__41017\
        );

    \I__8899\ : LocalMux
    port map (
            O => \N__41059\,
            I => \N__41017\
        );

    \I__8898\ : LocalMux
    port map (
            O => \N__41056\,
            I => \N__41012\
        );

    \I__8897\ : LocalMux
    port map (
            O => \N__41053\,
            I => \N__41012\
        );

    \I__8896\ : Span4Mux_v
    port map (
            O => \N__41046\,
            I => \N__41009\
        );

    \I__8895\ : LocalMux
    port map (
            O => \N__41043\,
            I => \N__41006\
        );

    \I__8894\ : LocalMux
    port map (
            O => \N__41040\,
            I => \N__41003\
        );

    \I__8893\ : LocalMux
    port map (
            O => \N__41037\,
            I => \N__41000\
        );

    \I__8892\ : LocalMux
    port map (
            O => \N__41034\,
            I => \N__40997\
        );

    \I__8891\ : LocalMux
    port map (
            O => \N__41031\,
            I => \N__40994\
        );

    \I__8890\ : Span4Mux_h
    port map (
            O => \N__41026\,
            I => \N__40987\
        );

    \I__8889\ : Span4Mux_h
    port map (
            O => \N__41017\,
            I => \N__40987\
        );

    \I__8888\ : Span4Mux_v
    port map (
            O => \N__41012\,
            I => \N__40987\
        );

    \I__8887\ : Span4Mux_h
    port map (
            O => \N__41009\,
            I => \N__40984\
        );

    \I__8886\ : Span4Mux_v
    port map (
            O => \N__41006\,
            I => \N__40979\
        );

    \I__8885\ : Span4Mux_v
    port map (
            O => \N__41003\,
            I => \N__40979\
        );

    \I__8884\ : Span4Mux_v
    port map (
            O => \N__41000\,
            I => \N__40970\
        );

    \I__8883\ : Span4Mux_v
    port map (
            O => \N__40997\,
            I => \N__40970\
        );

    \I__8882\ : Span4Mux_v
    port map (
            O => \N__40994\,
            I => \N__40970\
        );

    \I__8881\ : Span4Mux_h
    port map (
            O => \N__40987\,
            I => \N__40970\
        );

    \I__8880\ : Span4Mux_h
    port map (
            O => \N__40984\,
            I => \N__40967\
        );

    \I__8879\ : Sp12to4
    port map (
            O => \N__40979\,
            I => \N__40962\
        );

    \I__8878\ : Sp12to4
    port map (
            O => \N__40970\,
            I => \N__40962\
        );

    \I__8877\ : Span4Mux_h
    port map (
            O => \N__40967\,
            I => \N__40958\
        );

    \I__8876\ : Span12Mux_h
    port map (
            O => \N__40962\,
            I => \N__40955\
        );

    \I__8875\ : InMux
    port map (
            O => \N__40961\,
            I => \N__40952\
        );

    \I__8874\ : Odrv4
    port map (
            O => \N__40958\,
            I => \clk_RTD\
        );

    \I__8873\ : Odrv12
    port map (
            O => \N__40955\,
            I => \clk_RTD\
        );

    \I__8872\ : LocalMux
    port map (
            O => \N__40952\,
            I => \clk_RTD\
        );

    \I__8871\ : IoInMux
    port map (
            O => \N__40945\,
            I => \N__40942\
        );

    \I__8870\ : LocalMux
    port map (
            O => \N__40942\,
            I => \N__40939\
        );

    \I__8869\ : IoSpan4Mux
    port map (
            O => \N__40939\,
            I => \N__40935\
        );

    \I__8868\ : ClkMux
    port map (
            O => \N__40938\,
            I => \N__40932\
        );

    \I__8867\ : Span4Mux_s1_v
    port map (
            O => \N__40935\,
            I => \N__40929\
        );

    \I__8866\ : LocalMux
    port map (
            O => \N__40932\,
            I => \N__40925\
        );

    \I__8865\ : Sp12to4
    port map (
            O => \N__40929\,
            I => \N__40922\
        );

    \I__8864\ : ClkMux
    port map (
            O => \N__40928\,
            I => \N__40919\
        );

    \I__8863\ : Span4Mux_h
    port map (
            O => \N__40925\,
            I => \N__40916\
        );

    \I__8862\ : Span12Mux_h
    port map (
            O => \N__40922\,
            I => \N__40913\
        );

    \I__8861\ : LocalMux
    port map (
            O => \N__40919\,
            I => \N__40910\
        );

    \I__8860\ : Span4Mux_v
    port map (
            O => \N__40916\,
            I => \N__40907\
        );

    \I__8859\ : Span12Mux_v
    port map (
            O => \N__40913\,
            I => \N__40901\
        );

    \I__8858\ : Span12Mux_h
    port map (
            O => \N__40910\,
            I => \N__40901\
        );

    \I__8857\ : Span4Mux_h
    port map (
            O => \N__40907\,
            I => \N__40898\
        );

    \I__8856\ : InMux
    port map (
            O => \N__40906\,
            I => \N__40895\
        );

    \I__8855\ : Odrv12
    port map (
            O => \N__40901\,
            I => \TEST_LED\
        );

    \I__8854\ : Odrv4
    port map (
            O => \N__40898\,
            I => \TEST_LED\
        );

    \I__8853\ : LocalMux
    port map (
            O => \N__40895\,
            I => \TEST_LED\
        );

    \I__8852\ : InMux
    port map (
            O => \N__40888\,
            I => \N__40885\
        );

    \I__8851\ : LocalMux
    port map (
            O => \N__40885\,
            I => \N__40882\
        );

    \I__8850\ : Span4Mux_h
    port map (
            O => \N__40882\,
            I => \N__40878\
        );

    \I__8849\ : CascadeMux
    port map (
            O => \N__40881\,
            I => \N__40875\
        );

    \I__8848\ : Span4Mux_v
    port map (
            O => \N__40878\,
            I => \N__40872\
        );

    \I__8847\ : InMux
    port map (
            O => \N__40875\,
            I => \N__40869\
        );

    \I__8846\ : Odrv4
    port map (
            O => \N__40872\,
            I => buf_adcdata_vdc_6
        );

    \I__8845\ : LocalMux
    port map (
            O => \N__40869\,
            I => buf_adcdata_vdc_6
        );

    \I__8844\ : InMux
    port map (
            O => \N__40864\,
            I => \N__40861\
        );

    \I__8843\ : LocalMux
    port map (
            O => \N__40861\,
            I => \N__40857\
        );

    \I__8842\ : InMux
    port map (
            O => \N__40860\,
            I => \N__40854\
        );

    \I__8841\ : Span4Mux_v
    port map (
            O => \N__40857\,
            I => \N__40850\
        );

    \I__8840\ : LocalMux
    port map (
            O => \N__40854\,
            I => \N__40847\
        );

    \I__8839\ : InMux
    port map (
            O => \N__40853\,
            I => \N__40844\
        );

    \I__8838\ : Sp12to4
    port map (
            O => \N__40850\,
            I => \N__40841\
        );

    \I__8837\ : Span4Mux_v
    port map (
            O => \N__40847\,
            I => \N__40838\
        );

    \I__8836\ : LocalMux
    port map (
            O => \N__40844\,
            I => buf_adcdata_vac_6
        );

    \I__8835\ : Odrv12
    port map (
            O => \N__40841\,
            I => buf_adcdata_vac_6
        );

    \I__8834\ : Odrv4
    port map (
            O => \N__40838\,
            I => buf_adcdata_vac_6
        );

    \I__8833\ : InMux
    port map (
            O => \N__40831\,
            I => \N__40828\
        );

    \I__8832\ : LocalMux
    port map (
            O => \N__40828\,
            I => n19_adj_1593
        );

    \I__8831\ : CascadeMux
    port map (
            O => \N__40825\,
            I => \N__40822\
        );

    \I__8830\ : InMux
    port map (
            O => \N__40822\,
            I => \N__40819\
        );

    \I__8829\ : LocalMux
    port map (
            O => \N__40819\,
            I => \N__40816\
        );

    \I__8828\ : Odrv12
    port map (
            O => \N__40816\,
            I => n21071
        );

    \I__8827\ : InMux
    port map (
            O => \N__40813\,
            I => \N__40810\
        );

    \I__8826\ : LocalMux
    port map (
            O => \N__40810\,
            I => \N__40807\
        );

    \I__8825\ : Odrv4
    port map (
            O => \N__40807\,
            I => n20_adj_1607
        );

    \I__8824\ : InMux
    port map (
            O => \N__40804\,
            I => \N__40801\
        );

    \I__8823\ : LocalMux
    port map (
            O => \N__40801\,
            I => \N__40798\
        );

    \I__8822\ : Odrv12
    port map (
            O => \N__40798\,
            I => comm_buf_5_4
        );

    \I__8821\ : InMux
    port map (
            O => \N__40795\,
            I => \N__40792\
        );

    \I__8820\ : LocalMux
    port map (
            O => \N__40792\,
            I => \N__40789\
        );

    \I__8819\ : Odrv12
    port map (
            O => \N__40789\,
            I => comm_buf_4_4
        );

    \I__8818\ : InMux
    port map (
            O => \N__40786\,
            I => \N__40781\
        );

    \I__8817\ : InMux
    port map (
            O => \N__40785\,
            I => \N__40778\
        );

    \I__8816\ : InMux
    port map (
            O => \N__40784\,
            I => \N__40775\
        );

    \I__8815\ : LocalMux
    port map (
            O => \N__40781\,
            I => \N__40772\
        );

    \I__8814\ : LocalMux
    port map (
            O => \N__40778\,
            I => \N__40769\
        );

    \I__8813\ : LocalMux
    port map (
            O => \N__40775\,
            I => \N__40766\
        );

    \I__8812\ : Span4Mux_v
    port map (
            O => \N__40772\,
            I => \N__40763\
        );

    \I__8811\ : Span4Mux_v
    port map (
            O => \N__40769\,
            I => \N__40760\
        );

    \I__8810\ : Sp12to4
    port map (
            O => \N__40766\,
            I => \N__40757\
        );

    \I__8809\ : Sp12to4
    port map (
            O => \N__40763\,
            I => \N__40750\
        );

    \I__8808\ : Sp12to4
    port map (
            O => \N__40760\,
            I => \N__40750\
        );

    \I__8807\ : Span12Mux_v
    port map (
            O => \N__40757\,
            I => \N__40750\
        );

    \I__8806\ : Odrv12
    port map (
            O => \N__40750\,
            I => comm_buf_0_6
        );

    \I__8805\ : InMux
    port map (
            O => \N__40747\,
            I => \N__40744\
        );

    \I__8804\ : LocalMux
    port map (
            O => \N__40744\,
            I => n28
        );

    \I__8803\ : InMux
    port map (
            O => \N__40741\,
            I => \N__40738\
        );

    \I__8802\ : LocalMux
    port map (
            O => \N__40738\,
            I => n27
        );

    \I__8801\ : CascadeMux
    port map (
            O => \N__40735\,
            I => \n26_adj_1625_cascade_\
        );

    \I__8800\ : InMux
    port map (
            O => \N__40732\,
            I => \N__40729\
        );

    \I__8799\ : LocalMux
    port map (
            O => \N__40729\,
            I => n25_adj_1616
        );

    \I__8798\ : CascadeMux
    port map (
            O => \N__40726\,
            I => \n19553_cascade_\
        );

    \I__8797\ : SRMux
    port map (
            O => \N__40723\,
            I => \N__40720\
        );

    \I__8796\ : LocalMux
    port map (
            O => \N__40720\,
            I => \N__40717\
        );

    \I__8795\ : Span4Mux_v
    port map (
            O => \N__40717\,
            I => \N__40714\
        );

    \I__8794\ : Odrv4
    port map (
            O => \N__40714\,
            I => n17393
        );

    \I__8793\ : CascadeMux
    port map (
            O => \N__40711\,
            I => \N__40708\
        );

    \I__8792\ : InMux
    port map (
            O => \N__40708\,
            I => \N__40705\
        );

    \I__8791\ : LocalMux
    port map (
            O => \N__40705\,
            I => \N__40702\
        );

    \I__8790\ : Span4Mux_h
    port map (
            O => \N__40702\,
            I => \N__40699\
        );

    \I__8789\ : Span4Mux_v
    port map (
            O => \N__40699\,
            I => \N__40696\
        );

    \I__8788\ : Span4Mux_h
    port map (
            O => \N__40696\,
            I => \N__40693\
        );

    \I__8787\ : Odrv4
    port map (
            O => \N__40693\,
            I => n30
        );

    \I__8786\ : CascadeMux
    port map (
            O => \N__40690\,
            I => \comm_state_3_N_412_3_cascade_\
        );

    \I__8785\ : CascadeMux
    port map (
            O => \N__40687\,
            I => \n20700_cascade_\
        );

    \I__8784\ : SRMux
    port map (
            O => \N__40684\,
            I => \N__40680\
        );

    \I__8783\ : SRMux
    port map (
            O => \N__40683\,
            I => \N__40677\
        );

    \I__8782\ : LocalMux
    port map (
            O => \N__40680\,
            I => \N__40674\
        );

    \I__8781\ : LocalMux
    port map (
            O => \N__40677\,
            I => \N__40671\
        );

    \I__8780\ : Span4Mux_v
    port map (
            O => \N__40674\,
            I => \N__40668\
        );

    \I__8779\ : Span4Mux_h
    port map (
            O => \N__40671\,
            I => \N__40665\
        );

    \I__8778\ : Odrv4
    port map (
            O => \N__40668\,
            I => flagcntwd
        );

    \I__8777\ : Odrv4
    port map (
            O => \N__40665\,
            I => flagcntwd
        );

    \I__8776\ : CEMux
    port map (
            O => \N__40660\,
            I => \N__40657\
        );

    \I__8775\ : LocalMux
    port map (
            O => \N__40657\,
            I => \N__40654\
        );

    \I__8774\ : Span4Mux_h
    port map (
            O => \N__40654\,
            I => \N__40651\
        );

    \I__8773\ : Odrv4
    port map (
            O => \N__40651\,
            I => n11411
        );

    \I__8772\ : SRMux
    port map (
            O => \N__40648\,
            I => \N__40645\
        );

    \I__8771\ : LocalMux
    port map (
            O => \N__40645\,
            I => \N__40642\
        );

    \I__8770\ : Span4Mux_v
    port map (
            O => \N__40642\,
            I => \N__40638\
        );

    \I__8769\ : SRMux
    port map (
            O => \N__40641\,
            I => \N__40635\
        );

    \I__8768\ : Span4Mux_v
    port map (
            O => \N__40638\,
            I => \N__40632\
        );

    \I__8767\ : LocalMux
    port map (
            O => \N__40635\,
            I => \N__40629\
        );

    \I__8766\ : Span4Mux_h
    port map (
            O => \N__40632\,
            I => \N__40626\
        );

    \I__8765\ : Odrv4
    port map (
            O => \N__40629\,
            I => n20081
        );

    \I__8764\ : Odrv4
    port map (
            O => \N__40626\,
            I => n20081
        );

    \I__8763\ : CascadeMux
    port map (
            O => \N__40621\,
            I => \N__40618\
        );

    \I__8762\ : InMux
    port map (
            O => \N__40618\,
            I => \N__40615\
        );

    \I__8761\ : LocalMux
    port map (
            O => \N__40615\,
            I => \N__40612\
        );

    \I__8760\ : Span4Mux_h
    port map (
            O => \N__40612\,
            I => \N__40609\
        );

    \I__8759\ : Span4Mux_h
    port map (
            O => \N__40609\,
            I => \N__40606\
        );

    \I__8758\ : Odrv4
    port map (
            O => \N__40606\,
            I => n11333
        );

    \I__8757\ : CascadeMux
    port map (
            O => \N__40603\,
            I => \N__40600\
        );

    \I__8756\ : CascadeBuf
    port map (
            O => \N__40600\,
            I => \N__40597\
        );

    \I__8755\ : CascadeMux
    port map (
            O => \N__40597\,
            I => \N__40594\
        );

    \I__8754\ : CascadeBuf
    port map (
            O => \N__40594\,
            I => \N__40591\
        );

    \I__8753\ : CascadeMux
    port map (
            O => \N__40591\,
            I => \N__40588\
        );

    \I__8752\ : CascadeBuf
    port map (
            O => \N__40588\,
            I => \N__40585\
        );

    \I__8751\ : CascadeMux
    port map (
            O => \N__40585\,
            I => \N__40582\
        );

    \I__8750\ : CascadeBuf
    port map (
            O => \N__40582\,
            I => \N__40579\
        );

    \I__8749\ : CascadeMux
    port map (
            O => \N__40579\,
            I => \N__40576\
        );

    \I__8748\ : CascadeBuf
    port map (
            O => \N__40576\,
            I => \N__40573\
        );

    \I__8747\ : CascadeMux
    port map (
            O => \N__40573\,
            I => \N__40570\
        );

    \I__8746\ : CascadeBuf
    port map (
            O => \N__40570\,
            I => \N__40567\
        );

    \I__8745\ : CascadeMux
    port map (
            O => \N__40567\,
            I => \N__40564\
        );

    \I__8744\ : CascadeBuf
    port map (
            O => \N__40564\,
            I => \N__40561\
        );

    \I__8743\ : CascadeMux
    port map (
            O => \N__40561\,
            I => \N__40558\
        );

    \I__8742\ : CascadeBuf
    port map (
            O => \N__40558\,
            I => \N__40555\
        );

    \I__8741\ : CascadeMux
    port map (
            O => \N__40555\,
            I => \N__40552\
        );

    \I__8740\ : CascadeBuf
    port map (
            O => \N__40552\,
            I => \N__40548\
        );

    \I__8739\ : CascadeMux
    port map (
            O => \N__40551\,
            I => \N__40545\
        );

    \I__8738\ : CascadeMux
    port map (
            O => \N__40548\,
            I => \N__40542\
        );

    \I__8737\ : CascadeBuf
    port map (
            O => \N__40545\,
            I => \N__40539\
        );

    \I__8736\ : InMux
    port map (
            O => \N__40542\,
            I => \N__40536\
        );

    \I__8735\ : CascadeMux
    port map (
            O => \N__40539\,
            I => \N__40533\
        );

    \I__8734\ : LocalMux
    port map (
            O => \N__40536\,
            I => \N__40530\
        );

    \I__8733\ : InMux
    port map (
            O => \N__40533\,
            I => \N__40527\
        );

    \I__8732\ : Span4Mux_h
    port map (
            O => \N__40530\,
            I => \N__40524\
        );

    \I__8731\ : LocalMux
    port map (
            O => \N__40527\,
            I => \N__40520\
        );

    \I__8730\ : Span4Mux_h
    port map (
            O => \N__40524\,
            I => \N__40517\
        );

    \I__8729\ : InMux
    port map (
            O => \N__40523\,
            I => \N__40514\
        );

    \I__8728\ : Span12Mux_h
    port map (
            O => \N__40520\,
            I => \N__40511\
        );

    \I__8727\ : Span4Mux_h
    port map (
            O => \N__40517\,
            I => \N__40508\
        );

    \I__8726\ : LocalMux
    port map (
            O => \N__40514\,
            I => data_count_8
        );

    \I__8725\ : Odrv12
    port map (
            O => \N__40511\,
            I => data_count_8
        );

    \I__8724\ : Odrv4
    port map (
            O => \N__40508\,
            I => data_count_8
        );

    \I__8723\ : InMux
    port map (
            O => \N__40501\,
            I => \bfn_15_18_0_\
        );

    \I__8722\ : InMux
    port map (
            O => \N__40498\,
            I => n19295
        );

    \I__8721\ : CascadeMux
    port map (
            O => \N__40495\,
            I => \N__40492\
        );

    \I__8720\ : CascadeBuf
    port map (
            O => \N__40492\,
            I => \N__40489\
        );

    \I__8719\ : CascadeMux
    port map (
            O => \N__40489\,
            I => \N__40486\
        );

    \I__8718\ : CascadeBuf
    port map (
            O => \N__40486\,
            I => \N__40483\
        );

    \I__8717\ : CascadeMux
    port map (
            O => \N__40483\,
            I => \N__40480\
        );

    \I__8716\ : CascadeBuf
    port map (
            O => \N__40480\,
            I => \N__40477\
        );

    \I__8715\ : CascadeMux
    port map (
            O => \N__40477\,
            I => \N__40474\
        );

    \I__8714\ : CascadeBuf
    port map (
            O => \N__40474\,
            I => \N__40471\
        );

    \I__8713\ : CascadeMux
    port map (
            O => \N__40471\,
            I => \N__40468\
        );

    \I__8712\ : CascadeBuf
    port map (
            O => \N__40468\,
            I => \N__40465\
        );

    \I__8711\ : CascadeMux
    port map (
            O => \N__40465\,
            I => \N__40462\
        );

    \I__8710\ : CascadeBuf
    port map (
            O => \N__40462\,
            I => \N__40459\
        );

    \I__8709\ : CascadeMux
    port map (
            O => \N__40459\,
            I => \N__40456\
        );

    \I__8708\ : CascadeBuf
    port map (
            O => \N__40456\,
            I => \N__40453\
        );

    \I__8707\ : CascadeMux
    port map (
            O => \N__40453\,
            I => \N__40450\
        );

    \I__8706\ : CascadeBuf
    port map (
            O => \N__40450\,
            I => \N__40447\
        );

    \I__8705\ : CascadeMux
    port map (
            O => \N__40447\,
            I => \N__40443\
        );

    \I__8704\ : CascadeMux
    port map (
            O => \N__40446\,
            I => \N__40440\
        );

    \I__8703\ : CascadeBuf
    port map (
            O => \N__40443\,
            I => \N__40437\
        );

    \I__8702\ : CascadeBuf
    port map (
            O => \N__40440\,
            I => \N__40434\
        );

    \I__8701\ : CascadeMux
    port map (
            O => \N__40437\,
            I => \N__40431\
        );

    \I__8700\ : CascadeMux
    port map (
            O => \N__40434\,
            I => \N__40428\
        );

    \I__8699\ : InMux
    port map (
            O => \N__40431\,
            I => \N__40425\
        );

    \I__8698\ : InMux
    port map (
            O => \N__40428\,
            I => \N__40422\
        );

    \I__8697\ : LocalMux
    port map (
            O => \N__40425\,
            I => \N__40419\
        );

    \I__8696\ : LocalMux
    port map (
            O => \N__40422\,
            I => \N__40416\
        );

    \I__8695\ : Span4Mux_h
    port map (
            O => \N__40419\,
            I => \N__40413\
        );

    \I__8694\ : Span4Mux_h
    port map (
            O => \N__40416\,
            I => \N__40409\
        );

    \I__8693\ : Span4Mux_h
    port map (
            O => \N__40413\,
            I => \N__40406\
        );

    \I__8692\ : InMux
    port map (
            O => \N__40412\,
            I => \N__40403\
        );

    \I__8691\ : Span4Mux_v
    port map (
            O => \N__40409\,
            I => \N__40400\
        );

    \I__8690\ : Span4Mux_h
    port map (
            O => \N__40406\,
            I => \N__40397\
        );

    \I__8689\ : LocalMux
    port map (
            O => \N__40403\,
            I => data_count_9
        );

    \I__8688\ : Odrv4
    port map (
            O => \N__40400\,
            I => data_count_9
        );

    \I__8687\ : Odrv4
    port map (
            O => \N__40397\,
            I => data_count_9
        );

    \I__8686\ : CascadeMux
    port map (
            O => \N__40390\,
            I => \N__40387\
        );

    \I__8685\ : InMux
    port map (
            O => \N__40387\,
            I => \N__40384\
        );

    \I__8684\ : LocalMux
    port map (
            O => \N__40384\,
            I => \N__40381\
        );

    \I__8683\ : Span4Mux_h
    port map (
            O => \N__40381\,
            I => \N__40378\
        );

    \I__8682\ : Odrv4
    port map (
            O => \N__40378\,
            I => \SIG_DDS.tmp_buf_14\
        );

    \I__8681\ : InMux
    port map (
            O => \N__40375\,
            I => \N__40370\
        );

    \I__8680\ : InMux
    port map (
            O => \N__40374\,
            I => \N__40367\
        );

    \I__8679\ : CascadeMux
    port map (
            O => \N__40373\,
            I => \N__40364\
        );

    \I__8678\ : LocalMux
    port map (
            O => \N__40370\,
            I => \N__40361\
        );

    \I__8677\ : LocalMux
    port map (
            O => \N__40367\,
            I => \N__40358\
        );

    \I__8676\ : InMux
    port map (
            O => \N__40364\,
            I => \N__40355\
        );

    \I__8675\ : Span4Mux_h
    port map (
            O => \N__40361\,
            I => \N__40352\
        );

    \I__8674\ : Span4Mux_h
    port map (
            O => \N__40358\,
            I => \N__40349\
        );

    \I__8673\ : LocalMux
    port map (
            O => \N__40355\,
            I => buf_dds0_0
        );

    \I__8672\ : Odrv4
    port map (
            O => \N__40352\,
            I => buf_dds0_0
        );

    \I__8671\ : Odrv4
    port map (
            O => \N__40349\,
            I => buf_dds0_0
        );

    \I__8670\ : CascadeMux
    port map (
            O => \N__40342\,
            I => \N__40339\
        );

    \I__8669\ : InMux
    port map (
            O => \N__40339\,
            I => \N__40336\
        );

    \I__8668\ : LocalMux
    port map (
            O => \N__40336\,
            I => \N__40333\
        );

    \I__8667\ : Odrv4
    port map (
            O => \N__40333\,
            I => \SIG_DDS.tmp_buf_0\
        );

    \I__8666\ : CEMux
    port map (
            O => \N__40330\,
            I => \N__40326\
        );

    \I__8665\ : CEMux
    port map (
            O => \N__40329\,
            I => \N__40323\
        );

    \I__8664\ : LocalMux
    port map (
            O => \N__40326\,
            I => \N__40320\
        );

    \I__8663\ : LocalMux
    port map (
            O => \N__40323\,
            I => \N__40317\
        );

    \I__8662\ : Span4Mux_h
    port map (
            O => \N__40320\,
            I => \N__40311\
        );

    \I__8661\ : Span4Mux_h
    port map (
            O => \N__40317\,
            I => \N__40308\
        );

    \I__8660\ : CEMux
    port map (
            O => \N__40316\,
            I => \N__40305\
        );

    \I__8659\ : CEMux
    port map (
            O => \N__40315\,
            I => \N__40302\
        );

    \I__8658\ : CEMux
    port map (
            O => \N__40314\,
            I => \N__40299\
        );

    \I__8657\ : Odrv4
    port map (
            O => \N__40311\,
            I => \SIG_DDS.n12700\
        );

    \I__8656\ : Odrv4
    port map (
            O => \N__40308\,
            I => \SIG_DDS.n12700\
        );

    \I__8655\ : LocalMux
    port map (
            O => \N__40305\,
            I => \SIG_DDS.n12700\
        );

    \I__8654\ : LocalMux
    port map (
            O => \N__40302\,
            I => \SIG_DDS.n12700\
        );

    \I__8653\ : LocalMux
    port map (
            O => \N__40299\,
            I => \SIG_DDS.n12700\
        );

    \I__8652\ : InMux
    port map (
            O => \N__40288\,
            I => \N__40285\
        );

    \I__8651\ : LocalMux
    port map (
            O => \N__40285\,
            I => \N__40282\
        );

    \I__8650\ : Span4Mux_v
    port map (
            O => \N__40282\,
            I => \N__40279\
        );

    \I__8649\ : Span4Mux_v
    port map (
            O => \N__40279\,
            I => \N__40276\
        );

    \I__8648\ : Span4Mux_h
    port map (
            O => \N__40276\,
            I => \N__40271\
        );

    \I__8647\ : InMux
    port map (
            O => \N__40275\,
            I => \N__40266\
        );

    \I__8646\ : InMux
    port map (
            O => \N__40274\,
            I => \N__40266\
        );

    \I__8645\ : Odrv4
    port map (
            O => \N__40271\,
            I => comm_tx_buf_6
        );

    \I__8644\ : LocalMux
    port map (
            O => \N__40266\,
            I => comm_tx_buf_6
        );

    \I__8643\ : SRMux
    port map (
            O => \N__40261\,
            I => \N__40257\
        );

    \I__8642\ : SRMux
    port map (
            O => \N__40260\,
            I => \N__40253\
        );

    \I__8641\ : LocalMux
    port map (
            O => \N__40257\,
            I => \N__40250\
        );

    \I__8640\ : SRMux
    port map (
            O => \N__40256\,
            I => \N__40247\
        );

    \I__8639\ : LocalMux
    port map (
            O => \N__40253\,
            I => \N__40242\
        );

    \I__8638\ : Span4Mux_h
    port map (
            O => \N__40250\,
            I => \N__40242\
        );

    \I__8637\ : LocalMux
    port map (
            O => \N__40247\,
            I => \N__40239\
        );

    \I__8636\ : Odrv4
    port map (
            O => \N__40242\,
            I => \comm_spi.data_tx_7__N_758\
        );

    \I__8635\ : Odrv4
    port map (
            O => \N__40239\,
            I => \comm_spi.data_tx_7__N_758\
        );

    \I__8634\ : InMux
    port map (
            O => \N__40234\,
            I => \N__40231\
        );

    \I__8633\ : LocalMux
    port map (
            O => \N__40231\,
            I => \N__40226\
        );

    \I__8632\ : InMux
    port map (
            O => \N__40230\,
            I => \N__40223\
        );

    \I__8631\ : InMux
    port map (
            O => \N__40229\,
            I => \N__40220\
        );

    \I__8630\ : Odrv4
    port map (
            O => \N__40226\,
            I => \comm_spi.n22623\
        );

    \I__8629\ : LocalMux
    port map (
            O => \N__40223\,
            I => \comm_spi.n22623\
        );

    \I__8628\ : LocalMux
    port map (
            O => \N__40220\,
            I => \comm_spi.n22623\
        );

    \I__8627\ : InMux
    port map (
            O => \N__40213\,
            I => \N__40210\
        );

    \I__8626\ : LocalMux
    port map (
            O => \N__40210\,
            I => \N__40206\
        );

    \I__8625\ : InMux
    port map (
            O => \N__40209\,
            I => \N__40203\
        );

    \I__8624\ : Span4Mux_v
    port map (
            O => \N__40206\,
            I => \N__40200\
        );

    \I__8623\ : LocalMux
    port map (
            O => \N__40203\,
            I => \N__40197\
        );

    \I__8622\ : Odrv4
    port map (
            O => \N__40200\,
            I => \comm_spi.n14592\
        );

    \I__8621\ : Odrv4
    port map (
            O => \N__40197\,
            I => \comm_spi.n14592\
        );

    \I__8620\ : InMux
    port map (
            O => \N__40192\,
            I => \N__40189\
        );

    \I__8619\ : LocalMux
    port map (
            O => \N__40189\,
            I => \N__40186\
        );

    \I__8618\ : Span4Mux_v
    port map (
            O => \N__40186\,
            I => \N__40182\
        );

    \I__8617\ : InMux
    port map (
            O => \N__40185\,
            I => \N__40179\
        );

    \I__8616\ : Odrv4
    port map (
            O => \N__40182\,
            I => \comm_spi.n14593\
        );

    \I__8615\ : LocalMux
    port map (
            O => \N__40179\,
            I => \comm_spi.n14593\
        );

    \I__8614\ : CascadeMux
    port map (
            O => \N__40174\,
            I => \N__40171\
        );

    \I__8613\ : CascadeBuf
    port map (
            O => \N__40171\,
            I => \N__40168\
        );

    \I__8612\ : CascadeMux
    port map (
            O => \N__40168\,
            I => \N__40165\
        );

    \I__8611\ : CascadeBuf
    port map (
            O => \N__40165\,
            I => \N__40162\
        );

    \I__8610\ : CascadeMux
    port map (
            O => \N__40162\,
            I => \N__40159\
        );

    \I__8609\ : CascadeBuf
    port map (
            O => \N__40159\,
            I => \N__40156\
        );

    \I__8608\ : CascadeMux
    port map (
            O => \N__40156\,
            I => \N__40153\
        );

    \I__8607\ : CascadeBuf
    port map (
            O => \N__40153\,
            I => \N__40150\
        );

    \I__8606\ : CascadeMux
    port map (
            O => \N__40150\,
            I => \N__40147\
        );

    \I__8605\ : CascadeBuf
    port map (
            O => \N__40147\,
            I => \N__40144\
        );

    \I__8604\ : CascadeMux
    port map (
            O => \N__40144\,
            I => \N__40141\
        );

    \I__8603\ : CascadeBuf
    port map (
            O => \N__40141\,
            I => \N__40138\
        );

    \I__8602\ : CascadeMux
    port map (
            O => \N__40138\,
            I => \N__40135\
        );

    \I__8601\ : CascadeBuf
    port map (
            O => \N__40135\,
            I => \N__40132\
        );

    \I__8600\ : CascadeMux
    port map (
            O => \N__40132\,
            I => \N__40129\
        );

    \I__8599\ : CascadeBuf
    port map (
            O => \N__40129\,
            I => \N__40126\
        );

    \I__8598\ : CascadeMux
    port map (
            O => \N__40126\,
            I => \N__40122\
        );

    \I__8597\ : CascadeMux
    port map (
            O => \N__40125\,
            I => \N__40119\
        );

    \I__8596\ : CascadeBuf
    port map (
            O => \N__40122\,
            I => \N__40116\
        );

    \I__8595\ : CascadeBuf
    port map (
            O => \N__40119\,
            I => \N__40113\
        );

    \I__8594\ : CascadeMux
    port map (
            O => \N__40116\,
            I => \N__40110\
        );

    \I__8593\ : CascadeMux
    port map (
            O => \N__40113\,
            I => \N__40107\
        );

    \I__8592\ : InMux
    port map (
            O => \N__40110\,
            I => \N__40104\
        );

    \I__8591\ : InMux
    port map (
            O => \N__40107\,
            I => \N__40101\
        );

    \I__8590\ : LocalMux
    port map (
            O => \N__40104\,
            I => \N__40098\
        );

    \I__8589\ : LocalMux
    port map (
            O => \N__40101\,
            I => \N__40094\
        );

    \I__8588\ : Span4Mux_v
    port map (
            O => \N__40098\,
            I => \N__40091\
        );

    \I__8587\ : CascadeMux
    port map (
            O => \N__40097\,
            I => \N__40088\
        );

    \I__8586\ : Span4Mux_v
    port map (
            O => \N__40094\,
            I => \N__40085\
        );

    \I__8585\ : Span4Mux_h
    port map (
            O => \N__40091\,
            I => \N__40082\
        );

    \I__8584\ : InMux
    port map (
            O => \N__40088\,
            I => \N__40079\
        );

    \I__8583\ : Span4Mux_h
    port map (
            O => \N__40085\,
            I => \N__40074\
        );

    \I__8582\ : Span4Mux_h
    port map (
            O => \N__40082\,
            I => \N__40074\
        );

    \I__8581\ : LocalMux
    port map (
            O => \N__40079\,
            I => data_count_0
        );

    \I__8580\ : Odrv4
    port map (
            O => \N__40074\,
            I => data_count_0
        );

    \I__8579\ : CascadeMux
    port map (
            O => \N__40069\,
            I => \N__40066\
        );

    \I__8578\ : CascadeBuf
    port map (
            O => \N__40066\,
            I => \N__40063\
        );

    \I__8577\ : CascadeMux
    port map (
            O => \N__40063\,
            I => \N__40060\
        );

    \I__8576\ : CascadeBuf
    port map (
            O => \N__40060\,
            I => \N__40057\
        );

    \I__8575\ : CascadeMux
    port map (
            O => \N__40057\,
            I => \N__40054\
        );

    \I__8574\ : CascadeBuf
    port map (
            O => \N__40054\,
            I => \N__40051\
        );

    \I__8573\ : CascadeMux
    port map (
            O => \N__40051\,
            I => \N__40048\
        );

    \I__8572\ : CascadeBuf
    port map (
            O => \N__40048\,
            I => \N__40045\
        );

    \I__8571\ : CascadeMux
    port map (
            O => \N__40045\,
            I => \N__40042\
        );

    \I__8570\ : CascadeBuf
    port map (
            O => \N__40042\,
            I => \N__40039\
        );

    \I__8569\ : CascadeMux
    port map (
            O => \N__40039\,
            I => \N__40036\
        );

    \I__8568\ : CascadeBuf
    port map (
            O => \N__40036\,
            I => \N__40033\
        );

    \I__8567\ : CascadeMux
    port map (
            O => \N__40033\,
            I => \N__40030\
        );

    \I__8566\ : CascadeBuf
    port map (
            O => \N__40030\,
            I => \N__40027\
        );

    \I__8565\ : CascadeMux
    port map (
            O => \N__40027\,
            I => \N__40024\
        );

    \I__8564\ : CascadeBuf
    port map (
            O => \N__40024\,
            I => \N__40021\
        );

    \I__8563\ : CascadeMux
    port map (
            O => \N__40021\,
            I => \N__40017\
        );

    \I__8562\ : CascadeMux
    port map (
            O => \N__40020\,
            I => \N__40014\
        );

    \I__8561\ : CascadeBuf
    port map (
            O => \N__40017\,
            I => \N__40011\
        );

    \I__8560\ : CascadeBuf
    port map (
            O => \N__40014\,
            I => \N__40008\
        );

    \I__8559\ : CascadeMux
    port map (
            O => \N__40011\,
            I => \N__40005\
        );

    \I__8558\ : CascadeMux
    port map (
            O => \N__40008\,
            I => \N__40002\
        );

    \I__8557\ : InMux
    port map (
            O => \N__40005\,
            I => \N__39999\
        );

    \I__8556\ : InMux
    port map (
            O => \N__40002\,
            I => \N__39996\
        );

    \I__8555\ : LocalMux
    port map (
            O => \N__39999\,
            I => \N__39993\
        );

    \I__8554\ : LocalMux
    port map (
            O => \N__39996\,
            I => \N__39990\
        );

    \I__8553\ : Span4Mux_v
    port map (
            O => \N__39993\,
            I => \N__39987\
        );

    \I__8552\ : Span4Mux_v
    port map (
            O => \N__39990\,
            I => \N__39983\
        );

    \I__8551\ : Span4Mux_h
    port map (
            O => \N__39987\,
            I => \N__39980\
        );

    \I__8550\ : InMux
    port map (
            O => \N__39986\,
            I => \N__39977\
        );

    \I__8549\ : Span4Mux_h
    port map (
            O => \N__39983\,
            I => \N__39972\
        );

    \I__8548\ : Span4Mux_h
    port map (
            O => \N__39980\,
            I => \N__39972\
        );

    \I__8547\ : LocalMux
    port map (
            O => \N__39977\,
            I => data_count_1
        );

    \I__8546\ : Odrv4
    port map (
            O => \N__39972\,
            I => data_count_1
        );

    \I__8545\ : InMux
    port map (
            O => \N__39967\,
            I => n19287
        );

    \I__8544\ : CascadeMux
    port map (
            O => \N__39964\,
            I => \N__39961\
        );

    \I__8543\ : CascadeBuf
    port map (
            O => \N__39961\,
            I => \N__39958\
        );

    \I__8542\ : CascadeMux
    port map (
            O => \N__39958\,
            I => \N__39955\
        );

    \I__8541\ : CascadeBuf
    port map (
            O => \N__39955\,
            I => \N__39952\
        );

    \I__8540\ : CascadeMux
    port map (
            O => \N__39952\,
            I => \N__39949\
        );

    \I__8539\ : CascadeBuf
    port map (
            O => \N__39949\,
            I => \N__39946\
        );

    \I__8538\ : CascadeMux
    port map (
            O => \N__39946\,
            I => \N__39943\
        );

    \I__8537\ : CascadeBuf
    port map (
            O => \N__39943\,
            I => \N__39940\
        );

    \I__8536\ : CascadeMux
    port map (
            O => \N__39940\,
            I => \N__39937\
        );

    \I__8535\ : CascadeBuf
    port map (
            O => \N__39937\,
            I => \N__39934\
        );

    \I__8534\ : CascadeMux
    port map (
            O => \N__39934\,
            I => \N__39931\
        );

    \I__8533\ : CascadeBuf
    port map (
            O => \N__39931\,
            I => \N__39928\
        );

    \I__8532\ : CascadeMux
    port map (
            O => \N__39928\,
            I => \N__39925\
        );

    \I__8531\ : CascadeBuf
    port map (
            O => \N__39925\,
            I => \N__39922\
        );

    \I__8530\ : CascadeMux
    port map (
            O => \N__39922\,
            I => \N__39919\
        );

    \I__8529\ : CascadeBuf
    port map (
            O => \N__39919\,
            I => \N__39916\
        );

    \I__8528\ : CascadeMux
    port map (
            O => \N__39916\,
            I => \N__39912\
        );

    \I__8527\ : CascadeMux
    port map (
            O => \N__39915\,
            I => \N__39909\
        );

    \I__8526\ : CascadeBuf
    port map (
            O => \N__39912\,
            I => \N__39906\
        );

    \I__8525\ : CascadeBuf
    port map (
            O => \N__39909\,
            I => \N__39903\
        );

    \I__8524\ : CascadeMux
    port map (
            O => \N__39906\,
            I => \N__39900\
        );

    \I__8523\ : CascadeMux
    port map (
            O => \N__39903\,
            I => \N__39897\
        );

    \I__8522\ : InMux
    port map (
            O => \N__39900\,
            I => \N__39894\
        );

    \I__8521\ : InMux
    port map (
            O => \N__39897\,
            I => \N__39891\
        );

    \I__8520\ : LocalMux
    port map (
            O => \N__39894\,
            I => \N__39888\
        );

    \I__8519\ : LocalMux
    port map (
            O => \N__39891\,
            I => \N__39885\
        );

    \I__8518\ : Span4Mux_h
    port map (
            O => \N__39888\,
            I => \N__39882\
        );

    \I__8517\ : Span4Mux_h
    port map (
            O => \N__39885\,
            I => \N__39878\
        );

    \I__8516\ : Span4Mux_h
    port map (
            O => \N__39882\,
            I => \N__39875\
        );

    \I__8515\ : InMux
    port map (
            O => \N__39881\,
            I => \N__39872\
        );

    \I__8514\ : Span4Mux_h
    port map (
            O => \N__39878\,
            I => \N__39869\
        );

    \I__8513\ : Span4Mux_h
    port map (
            O => \N__39875\,
            I => \N__39866\
        );

    \I__8512\ : LocalMux
    port map (
            O => \N__39872\,
            I => data_count_2
        );

    \I__8511\ : Odrv4
    port map (
            O => \N__39869\,
            I => data_count_2
        );

    \I__8510\ : Odrv4
    port map (
            O => \N__39866\,
            I => data_count_2
        );

    \I__8509\ : InMux
    port map (
            O => \N__39859\,
            I => n19288
        );

    \I__8508\ : CascadeMux
    port map (
            O => \N__39856\,
            I => \N__39853\
        );

    \I__8507\ : CascadeBuf
    port map (
            O => \N__39853\,
            I => \N__39850\
        );

    \I__8506\ : CascadeMux
    port map (
            O => \N__39850\,
            I => \N__39847\
        );

    \I__8505\ : CascadeBuf
    port map (
            O => \N__39847\,
            I => \N__39844\
        );

    \I__8504\ : CascadeMux
    port map (
            O => \N__39844\,
            I => \N__39841\
        );

    \I__8503\ : CascadeBuf
    port map (
            O => \N__39841\,
            I => \N__39838\
        );

    \I__8502\ : CascadeMux
    port map (
            O => \N__39838\,
            I => \N__39835\
        );

    \I__8501\ : CascadeBuf
    port map (
            O => \N__39835\,
            I => \N__39832\
        );

    \I__8500\ : CascadeMux
    port map (
            O => \N__39832\,
            I => \N__39829\
        );

    \I__8499\ : CascadeBuf
    port map (
            O => \N__39829\,
            I => \N__39826\
        );

    \I__8498\ : CascadeMux
    port map (
            O => \N__39826\,
            I => \N__39823\
        );

    \I__8497\ : CascadeBuf
    port map (
            O => \N__39823\,
            I => \N__39820\
        );

    \I__8496\ : CascadeMux
    port map (
            O => \N__39820\,
            I => \N__39817\
        );

    \I__8495\ : CascadeBuf
    port map (
            O => \N__39817\,
            I => \N__39814\
        );

    \I__8494\ : CascadeMux
    port map (
            O => \N__39814\,
            I => \N__39810\
        );

    \I__8493\ : CascadeMux
    port map (
            O => \N__39813\,
            I => \N__39807\
        );

    \I__8492\ : CascadeBuf
    port map (
            O => \N__39810\,
            I => \N__39804\
        );

    \I__8491\ : CascadeBuf
    port map (
            O => \N__39807\,
            I => \N__39801\
        );

    \I__8490\ : CascadeMux
    port map (
            O => \N__39804\,
            I => \N__39798\
        );

    \I__8489\ : CascadeMux
    port map (
            O => \N__39801\,
            I => \N__39795\
        );

    \I__8488\ : CascadeBuf
    port map (
            O => \N__39798\,
            I => \N__39792\
        );

    \I__8487\ : InMux
    port map (
            O => \N__39795\,
            I => \N__39789\
        );

    \I__8486\ : CascadeMux
    port map (
            O => \N__39792\,
            I => \N__39786\
        );

    \I__8485\ : LocalMux
    port map (
            O => \N__39789\,
            I => \N__39783\
        );

    \I__8484\ : InMux
    port map (
            O => \N__39786\,
            I => \N__39780\
        );

    \I__8483\ : Span4Mux_h
    port map (
            O => \N__39783\,
            I => \N__39776\
        );

    \I__8482\ : LocalMux
    port map (
            O => \N__39780\,
            I => \N__39773\
        );

    \I__8481\ : InMux
    port map (
            O => \N__39779\,
            I => \N__39770\
        );

    \I__8480\ : Span4Mux_h
    port map (
            O => \N__39776\,
            I => \N__39767\
        );

    \I__8479\ : Span12Mux_h
    port map (
            O => \N__39773\,
            I => \N__39764\
        );

    \I__8478\ : LocalMux
    port map (
            O => \N__39770\,
            I => data_count_3
        );

    \I__8477\ : Odrv4
    port map (
            O => \N__39767\,
            I => data_count_3
        );

    \I__8476\ : Odrv12
    port map (
            O => \N__39764\,
            I => data_count_3
        );

    \I__8475\ : InMux
    port map (
            O => \N__39757\,
            I => n19289
        );

    \I__8474\ : CascadeMux
    port map (
            O => \N__39754\,
            I => \N__39751\
        );

    \I__8473\ : CascadeBuf
    port map (
            O => \N__39751\,
            I => \N__39748\
        );

    \I__8472\ : CascadeMux
    port map (
            O => \N__39748\,
            I => \N__39745\
        );

    \I__8471\ : CascadeBuf
    port map (
            O => \N__39745\,
            I => \N__39742\
        );

    \I__8470\ : CascadeMux
    port map (
            O => \N__39742\,
            I => \N__39739\
        );

    \I__8469\ : CascadeBuf
    port map (
            O => \N__39739\,
            I => \N__39736\
        );

    \I__8468\ : CascadeMux
    port map (
            O => \N__39736\,
            I => \N__39733\
        );

    \I__8467\ : CascadeBuf
    port map (
            O => \N__39733\,
            I => \N__39730\
        );

    \I__8466\ : CascadeMux
    port map (
            O => \N__39730\,
            I => \N__39727\
        );

    \I__8465\ : CascadeBuf
    port map (
            O => \N__39727\,
            I => \N__39724\
        );

    \I__8464\ : CascadeMux
    port map (
            O => \N__39724\,
            I => \N__39721\
        );

    \I__8463\ : CascadeBuf
    port map (
            O => \N__39721\,
            I => \N__39718\
        );

    \I__8462\ : CascadeMux
    port map (
            O => \N__39718\,
            I => \N__39715\
        );

    \I__8461\ : CascadeBuf
    port map (
            O => \N__39715\,
            I => \N__39712\
        );

    \I__8460\ : CascadeMux
    port map (
            O => \N__39712\,
            I => \N__39709\
        );

    \I__8459\ : CascadeBuf
    port map (
            O => \N__39709\,
            I => \N__39706\
        );

    \I__8458\ : CascadeMux
    port map (
            O => \N__39706\,
            I => \N__39702\
        );

    \I__8457\ : CascadeMux
    port map (
            O => \N__39705\,
            I => \N__39699\
        );

    \I__8456\ : CascadeBuf
    port map (
            O => \N__39702\,
            I => \N__39696\
        );

    \I__8455\ : CascadeBuf
    port map (
            O => \N__39699\,
            I => \N__39693\
        );

    \I__8454\ : CascadeMux
    port map (
            O => \N__39696\,
            I => \N__39690\
        );

    \I__8453\ : CascadeMux
    port map (
            O => \N__39693\,
            I => \N__39687\
        );

    \I__8452\ : InMux
    port map (
            O => \N__39690\,
            I => \N__39684\
        );

    \I__8451\ : InMux
    port map (
            O => \N__39687\,
            I => \N__39681\
        );

    \I__8450\ : LocalMux
    port map (
            O => \N__39684\,
            I => \N__39678\
        );

    \I__8449\ : LocalMux
    port map (
            O => \N__39681\,
            I => \N__39675\
        );

    \I__8448\ : Span4Mux_h
    port map (
            O => \N__39678\,
            I => \N__39672\
        );

    \I__8447\ : Span4Mux_v
    port map (
            O => \N__39675\,
            I => \N__39668\
        );

    \I__8446\ : Span4Mux_h
    port map (
            O => \N__39672\,
            I => \N__39665\
        );

    \I__8445\ : InMux
    port map (
            O => \N__39671\,
            I => \N__39662\
        );

    \I__8444\ : Span4Mux_h
    port map (
            O => \N__39668\,
            I => \N__39659\
        );

    \I__8443\ : Span4Mux_h
    port map (
            O => \N__39665\,
            I => \N__39656\
        );

    \I__8442\ : LocalMux
    port map (
            O => \N__39662\,
            I => data_count_4
        );

    \I__8441\ : Odrv4
    port map (
            O => \N__39659\,
            I => data_count_4
        );

    \I__8440\ : Odrv4
    port map (
            O => \N__39656\,
            I => data_count_4
        );

    \I__8439\ : InMux
    port map (
            O => \N__39649\,
            I => n19290
        );

    \I__8438\ : CascadeMux
    port map (
            O => \N__39646\,
            I => \N__39643\
        );

    \I__8437\ : CascadeBuf
    port map (
            O => \N__39643\,
            I => \N__39640\
        );

    \I__8436\ : CascadeMux
    port map (
            O => \N__39640\,
            I => \N__39637\
        );

    \I__8435\ : CascadeBuf
    port map (
            O => \N__39637\,
            I => \N__39634\
        );

    \I__8434\ : CascadeMux
    port map (
            O => \N__39634\,
            I => \N__39631\
        );

    \I__8433\ : CascadeBuf
    port map (
            O => \N__39631\,
            I => \N__39628\
        );

    \I__8432\ : CascadeMux
    port map (
            O => \N__39628\,
            I => \N__39625\
        );

    \I__8431\ : CascadeBuf
    port map (
            O => \N__39625\,
            I => \N__39622\
        );

    \I__8430\ : CascadeMux
    port map (
            O => \N__39622\,
            I => \N__39619\
        );

    \I__8429\ : CascadeBuf
    port map (
            O => \N__39619\,
            I => \N__39616\
        );

    \I__8428\ : CascadeMux
    port map (
            O => \N__39616\,
            I => \N__39613\
        );

    \I__8427\ : CascadeBuf
    port map (
            O => \N__39613\,
            I => \N__39610\
        );

    \I__8426\ : CascadeMux
    port map (
            O => \N__39610\,
            I => \N__39607\
        );

    \I__8425\ : CascadeBuf
    port map (
            O => \N__39607\,
            I => \N__39604\
        );

    \I__8424\ : CascadeMux
    port map (
            O => \N__39604\,
            I => \N__39601\
        );

    \I__8423\ : CascadeBuf
    port map (
            O => \N__39601\,
            I => \N__39598\
        );

    \I__8422\ : CascadeMux
    port map (
            O => \N__39598\,
            I => \N__39594\
        );

    \I__8421\ : CascadeMux
    port map (
            O => \N__39597\,
            I => \N__39591\
        );

    \I__8420\ : CascadeBuf
    port map (
            O => \N__39594\,
            I => \N__39588\
        );

    \I__8419\ : CascadeBuf
    port map (
            O => \N__39591\,
            I => \N__39585\
        );

    \I__8418\ : CascadeMux
    port map (
            O => \N__39588\,
            I => \N__39582\
        );

    \I__8417\ : CascadeMux
    port map (
            O => \N__39585\,
            I => \N__39579\
        );

    \I__8416\ : InMux
    port map (
            O => \N__39582\,
            I => \N__39576\
        );

    \I__8415\ : InMux
    port map (
            O => \N__39579\,
            I => \N__39573\
        );

    \I__8414\ : LocalMux
    port map (
            O => \N__39576\,
            I => \N__39570\
        );

    \I__8413\ : LocalMux
    port map (
            O => \N__39573\,
            I => \N__39567\
        );

    \I__8412\ : Span4Mux_h
    port map (
            O => \N__39570\,
            I => \N__39564\
        );

    \I__8411\ : Span4Mux_v
    port map (
            O => \N__39567\,
            I => \N__39560\
        );

    \I__8410\ : Span4Mux_h
    port map (
            O => \N__39564\,
            I => \N__39557\
        );

    \I__8409\ : InMux
    port map (
            O => \N__39563\,
            I => \N__39554\
        );

    \I__8408\ : Span4Mux_h
    port map (
            O => \N__39560\,
            I => \N__39551\
        );

    \I__8407\ : Span4Mux_h
    port map (
            O => \N__39557\,
            I => \N__39548\
        );

    \I__8406\ : LocalMux
    port map (
            O => \N__39554\,
            I => data_count_5
        );

    \I__8405\ : Odrv4
    port map (
            O => \N__39551\,
            I => data_count_5
        );

    \I__8404\ : Odrv4
    port map (
            O => \N__39548\,
            I => data_count_5
        );

    \I__8403\ : InMux
    port map (
            O => \N__39541\,
            I => n19291
        );

    \I__8402\ : CascadeMux
    port map (
            O => \N__39538\,
            I => \N__39535\
        );

    \I__8401\ : CascadeBuf
    port map (
            O => \N__39535\,
            I => \N__39532\
        );

    \I__8400\ : CascadeMux
    port map (
            O => \N__39532\,
            I => \N__39529\
        );

    \I__8399\ : CascadeBuf
    port map (
            O => \N__39529\,
            I => \N__39526\
        );

    \I__8398\ : CascadeMux
    port map (
            O => \N__39526\,
            I => \N__39523\
        );

    \I__8397\ : CascadeBuf
    port map (
            O => \N__39523\,
            I => \N__39520\
        );

    \I__8396\ : CascadeMux
    port map (
            O => \N__39520\,
            I => \N__39517\
        );

    \I__8395\ : CascadeBuf
    port map (
            O => \N__39517\,
            I => \N__39514\
        );

    \I__8394\ : CascadeMux
    port map (
            O => \N__39514\,
            I => \N__39511\
        );

    \I__8393\ : CascadeBuf
    port map (
            O => \N__39511\,
            I => \N__39508\
        );

    \I__8392\ : CascadeMux
    port map (
            O => \N__39508\,
            I => \N__39505\
        );

    \I__8391\ : CascadeBuf
    port map (
            O => \N__39505\,
            I => \N__39502\
        );

    \I__8390\ : CascadeMux
    port map (
            O => \N__39502\,
            I => \N__39499\
        );

    \I__8389\ : CascadeBuf
    port map (
            O => \N__39499\,
            I => \N__39496\
        );

    \I__8388\ : CascadeMux
    port map (
            O => \N__39496\,
            I => \N__39493\
        );

    \I__8387\ : CascadeBuf
    port map (
            O => \N__39493\,
            I => \N__39489\
        );

    \I__8386\ : CascadeMux
    port map (
            O => \N__39492\,
            I => \N__39486\
        );

    \I__8385\ : CascadeMux
    port map (
            O => \N__39489\,
            I => \N__39483\
        );

    \I__8384\ : CascadeBuf
    port map (
            O => \N__39486\,
            I => \N__39480\
        );

    \I__8383\ : CascadeBuf
    port map (
            O => \N__39483\,
            I => \N__39477\
        );

    \I__8382\ : CascadeMux
    port map (
            O => \N__39480\,
            I => \N__39474\
        );

    \I__8381\ : CascadeMux
    port map (
            O => \N__39477\,
            I => \N__39471\
        );

    \I__8380\ : InMux
    port map (
            O => \N__39474\,
            I => \N__39468\
        );

    \I__8379\ : InMux
    port map (
            O => \N__39471\,
            I => \N__39465\
        );

    \I__8378\ : LocalMux
    port map (
            O => \N__39468\,
            I => \N__39462\
        );

    \I__8377\ : LocalMux
    port map (
            O => \N__39465\,
            I => \N__39459\
        );

    \I__8376\ : Span4Mux_h
    port map (
            O => \N__39462\,
            I => \N__39455\
        );

    \I__8375\ : Span4Mux_v
    port map (
            O => \N__39459\,
            I => \N__39452\
        );

    \I__8374\ : InMux
    port map (
            O => \N__39458\,
            I => \N__39449\
        );

    \I__8373\ : Span4Mux_h
    port map (
            O => \N__39455\,
            I => \N__39446\
        );

    \I__8372\ : Sp12to4
    port map (
            O => \N__39452\,
            I => \N__39443\
        );

    \I__8371\ : LocalMux
    port map (
            O => \N__39449\,
            I => data_count_6
        );

    \I__8370\ : Odrv4
    port map (
            O => \N__39446\,
            I => data_count_6
        );

    \I__8369\ : Odrv12
    port map (
            O => \N__39443\,
            I => data_count_6
        );

    \I__8368\ : InMux
    port map (
            O => \N__39436\,
            I => n19292
        );

    \I__8367\ : CascadeMux
    port map (
            O => \N__39433\,
            I => \N__39430\
        );

    \I__8366\ : CascadeBuf
    port map (
            O => \N__39430\,
            I => \N__39427\
        );

    \I__8365\ : CascadeMux
    port map (
            O => \N__39427\,
            I => \N__39424\
        );

    \I__8364\ : CascadeBuf
    port map (
            O => \N__39424\,
            I => \N__39421\
        );

    \I__8363\ : CascadeMux
    port map (
            O => \N__39421\,
            I => \N__39418\
        );

    \I__8362\ : CascadeBuf
    port map (
            O => \N__39418\,
            I => \N__39415\
        );

    \I__8361\ : CascadeMux
    port map (
            O => \N__39415\,
            I => \N__39412\
        );

    \I__8360\ : CascadeBuf
    port map (
            O => \N__39412\,
            I => \N__39409\
        );

    \I__8359\ : CascadeMux
    port map (
            O => \N__39409\,
            I => \N__39406\
        );

    \I__8358\ : CascadeBuf
    port map (
            O => \N__39406\,
            I => \N__39403\
        );

    \I__8357\ : CascadeMux
    port map (
            O => \N__39403\,
            I => \N__39400\
        );

    \I__8356\ : CascadeBuf
    port map (
            O => \N__39400\,
            I => \N__39397\
        );

    \I__8355\ : CascadeMux
    port map (
            O => \N__39397\,
            I => \N__39394\
        );

    \I__8354\ : CascadeBuf
    port map (
            O => \N__39394\,
            I => \N__39391\
        );

    \I__8353\ : CascadeMux
    port map (
            O => \N__39391\,
            I => \N__39387\
        );

    \I__8352\ : CascadeMux
    port map (
            O => \N__39390\,
            I => \N__39384\
        );

    \I__8351\ : CascadeBuf
    port map (
            O => \N__39387\,
            I => \N__39381\
        );

    \I__8350\ : CascadeBuf
    port map (
            O => \N__39384\,
            I => \N__39378\
        );

    \I__8349\ : CascadeMux
    port map (
            O => \N__39381\,
            I => \N__39375\
        );

    \I__8348\ : CascadeMux
    port map (
            O => \N__39378\,
            I => \N__39372\
        );

    \I__8347\ : CascadeBuf
    port map (
            O => \N__39375\,
            I => \N__39369\
        );

    \I__8346\ : InMux
    port map (
            O => \N__39372\,
            I => \N__39366\
        );

    \I__8345\ : CascadeMux
    port map (
            O => \N__39369\,
            I => \N__39363\
        );

    \I__8344\ : LocalMux
    port map (
            O => \N__39366\,
            I => \N__39360\
        );

    \I__8343\ : InMux
    port map (
            O => \N__39363\,
            I => \N__39357\
        );

    \I__8342\ : Span4Mux_v
    port map (
            O => \N__39360\,
            I => \N__39353\
        );

    \I__8341\ : LocalMux
    port map (
            O => \N__39357\,
            I => \N__39350\
        );

    \I__8340\ : InMux
    port map (
            O => \N__39356\,
            I => \N__39347\
        );

    \I__8339\ : Span4Mux_h
    port map (
            O => \N__39353\,
            I => \N__39344\
        );

    \I__8338\ : Span12Mux_s9_v
    port map (
            O => \N__39350\,
            I => \N__39341\
        );

    \I__8337\ : LocalMux
    port map (
            O => \N__39347\,
            I => data_count_7
        );

    \I__8336\ : Odrv4
    port map (
            O => \N__39344\,
            I => data_count_7
        );

    \I__8335\ : Odrv12
    port map (
            O => \N__39341\,
            I => data_count_7
        );

    \I__8334\ : InMux
    port map (
            O => \N__39334\,
            I => n19293
        );

    \I__8333\ : CascadeMux
    port map (
            O => \N__39331\,
            I => \N__39324\
        );

    \I__8332\ : InMux
    port map (
            O => \N__39330\,
            I => \N__39318\
        );

    \I__8331\ : InMux
    port map (
            O => \N__39329\,
            I => \N__39318\
        );

    \I__8330\ : InMux
    port map (
            O => \N__39328\,
            I => \N__39308\
        );

    \I__8329\ : InMux
    port map (
            O => \N__39327\,
            I => \N__39308\
        );

    \I__8328\ : InMux
    port map (
            O => \N__39324\,
            I => \N__39303\
        );

    \I__8327\ : InMux
    port map (
            O => \N__39323\,
            I => \N__39303\
        );

    \I__8326\ : LocalMux
    port map (
            O => \N__39318\,
            I => \N__39300\
        );

    \I__8325\ : InMux
    port map (
            O => \N__39317\,
            I => \N__39293\
        );

    \I__8324\ : InMux
    port map (
            O => \N__39316\,
            I => \N__39293\
        );

    \I__8323\ : InMux
    port map (
            O => \N__39315\,
            I => \N__39293\
        );

    \I__8322\ : InMux
    port map (
            O => \N__39314\,
            I => \N__39288\
        );

    \I__8321\ : InMux
    port map (
            O => \N__39313\,
            I => \N__39288\
        );

    \I__8320\ : LocalMux
    port map (
            O => \N__39308\,
            I => \N__39280\
        );

    \I__8319\ : LocalMux
    port map (
            O => \N__39303\,
            I => \N__39280\
        );

    \I__8318\ : Span4Mux_v
    port map (
            O => \N__39300\,
            I => \N__39277\
        );

    \I__8317\ : LocalMux
    port map (
            O => \N__39293\,
            I => \N__39274\
        );

    \I__8316\ : LocalMux
    port map (
            O => \N__39288\,
            I => \N__39269\
        );

    \I__8315\ : InMux
    port map (
            O => \N__39287\,
            I => \N__39262\
        );

    \I__8314\ : InMux
    port map (
            O => \N__39286\,
            I => \N__39262\
        );

    \I__8313\ : InMux
    port map (
            O => \N__39285\,
            I => \N__39262\
        );

    \I__8312\ : Span4Mux_h
    port map (
            O => \N__39280\,
            I => \N__39255\
        );

    \I__8311\ : Span4Mux_h
    port map (
            O => \N__39277\,
            I => \N__39255\
        );

    \I__8310\ : Span4Mux_h
    port map (
            O => \N__39274\,
            I => \N__39255\
        );

    \I__8309\ : InMux
    port map (
            O => \N__39273\,
            I => \N__39250\
        );

    \I__8308\ : InMux
    port map (
            O => \N__39272\,
            I => \N__39250\
        );

    \I__8307\ : Odrv4
    port map (
            O => \N__39269\,
            I => n12391
        );

    \I__8306\ : LocalMux
    port map (
            O => \N__39262\,
            I => n12391
        );

    \I__8305\ : Odrv4
    port map (
            O => \N__39255\,
            I => n12391
        );

    \I__8304\ : LocalMux
    port map (
            O => \N__39250\,
            I => n12391
        );

    \I__8303\ : InMux
    port map (
            O => \N__39241\,
            I => \N__39233\
        );

    \I__8302\ : InMux
    port map (
            O => \N__39240\,
            I => \N__39226\
        );

    \I__8301\ : InMux
    port map (
            O => \N__39239\,
            I => \N__39226\
        );

    \I__8300\ : InMux
    port map (
            O => \N__39238\,
            I => \N__39226\
        );

    \I__8299\ : InMux
    port map (
            O => \N__39237\,
            I => \N__39223\
        );

    \I__8298\ : InMux
    port map (
            O => \N__39236\,
            I => \N__39220\
        );

    \I__8297\ : LocalMux
    port map (
            O => \N__39233\,
            I => \N__39212\
        );

    \I__8296\ : LocalMux
    port map (
            O => \N__39226\,
            I => \N__39212\
        );

    \I__8295\ : LocalMux
    port map (
            O => \N__39223\,
            I => \N__39212\
        );

    \I__8294\ : LocalMux
    port map (
            O => \N__39220\,
            I => \N__39209\
        );

    \I__8293\ : InMux
    port map (
            O => \N__39219\,
            I => \N__39206\
        );

    \I__8292\ : Span4Mux_v
    port map (
            O => \N__39212\,
            I => \N__39198\
        );

    \I__8291\ : Span4Mux_h
    port map (
            O => \N__39209\,
            I => \N__39198\
        );

    \I__8290\ : LocalMux
    port map (
            O => \N__39206\,
            I => \N__39198\
        );

    \I__8289\ : InMux
    port map (
            O => \N__39205\,
            I => \N__39195\
        );

    \I__8288\ : Sp12to4
    port map (
            O => \N__39198\,
            I => \N__39190\
        );

    \I__8287\ : LocalMux
    port map (
            O => \N__39195\,
            I => \N__39190\
        );

    \I__8286\ : Odrv12
    port map (
            O => \N__39190\,
            I => n12367
        );

    \I__8285\ : InMux
    port map (
            O => \N__39187\,
            I => \N__39184\
        );

    \I__8284\ : LocalMux
    port map (
            O => \N__39184\,
            I => \N__39180\
        );

    \I__8283\ : CascadeMux
    port map (
            O => \N__39183\,
            I => \N__39177\
        );

    \I__8282\ : Span4Mux_v
    port map (
            O => \N__39180\,
            I => \N__39174\
        );

    \I__8281\ : InMux
    port map (
            O => \N__39177\,
            I => \N__39171\
        );

    \I__8280\ : Span4Mux_h
    port map (
            O => \N__39174\,
            I => \N__39168\
        );

    \I__8279\ : LocalMux
    port map (
            O => \N__39171\,
            I => \N__39165\
        );

    \I__8278\ : Odrv4
    port map (
            O => \N__39168\,
            I => n11324
        );

    \I__8277\ : Odrv12
    port map (
            O => \N__39165\,
            I => n11324
        );

    \I__8276\ : CascadeMux
    port map (
            O => \N__39160\,
            I => \n8780_cascade_\
        );

    \I__8275\ : CascadeMux
    port map (
            O => \N__39157\,
            I => \N__39153\
        );

    \I__8274\ : InMux
    port map (
            O => \N__39156\,
            I => \N__39143\
        );

    \I__8273\ : InMux
    port map (
            O => \N__39153\,
            I => \N__39143\
        );

    \I__8272\ : InMux
    port map (
            O => \N__39152\,
            I => \N__39143\
        );

    \I__8271\ : CascadeMux
    port map (
            O => \N__39151\,
            I => \N__39138\
        );

    \I__8270\ : InMux
    port map (
            O => \N__39150\,
            I => \N__39134\
        );

    \I__8269\ : LocalMux
    port map (
            O => \N__39143\,
            I => \N__39131\
        );

    \I__8268\ : InMux
    port map (
            O => \N__39142\,
            I => \N__39128\
        );

    \I__8267\ : InMux
    port map (
            O => \N__39141\,
            I => \N__39123\
        );

    \I__8266\ : InMux
    port map (
            O => \N__39138\,
            I => \N__39123\
        );

    \I__8265\ : InMux
    port map (
            O => \N__39137\,
            I => \N__39119\
        );

    \I__8264\ : LocalMux
    port map (
            O => \N__39134\,
            I => \N__39116\
        );

    \I__8263\ : Span4Mux_v
    port map (
            O => \N__39131\,
            I => \N__39109\
        );

    \I__8262\ : LocalMux
    port map (
            O => \N__39128\,
            I => \N__39109\
        );

    \I__8261\ : LocalMux
    port map (
            O => \N__39123\,
            I => \N__39109\
        );

    \I__8260\ : CascadeMux
    port map (
            O => \N__39122\,
            I => \N__39102\
        );

    \I__8259\ : LocalMux
    port map (
            O => \N__39119\,
            I => \N__39099\
        );

    \I__8258\ : Span4Mux_v
    port map (
            O => \N__39116\,
            I => \N__39094\
        );

    \I__8257\ : Span4Mux_v
    port map (
            O => \N__39109\,
            I => \N__39094\
        );

    \I__8256\ : InMux
    port map (
            O => \N__39108\,
            I => \N__39089\
        );

    \I__8255\ : InMux
    port map (
            O => \N__39107\,
            I => \N__39089\
        );

    \I__8254\ : InMux
    port map (
            O => \N__39106\,
            I => \N__39086\
        );

    \I__8253\ : InMux
    port map (
            O => \N__39105\,
            I => \N__39081\
        );

    \I__8252\ : InMux
    port map (
            O => \N__39102\,
            I => \N__39081\
        );

    \I__8251\ : Span4Mux_v
    port map (
            O => \N__39099\,
            I => \N__39076\
        );

    \I__8250\ : Span4Mux_h
    port map (
            O => \N__39094\,
            I => \N__39076\
        );

    \I__8249\ : LocalMux
    port map (
            O => \N__39089\,
            I => \N__39073\
        );

    \I__8248\ : LocalMux
    port map (
            O => \N__39086\,
            I => eis_state_1
        );

    \I__8247\ : LocalMux
    port map (
            O => \N__39081\,
            I => eis_state_1
        );

    \I__8246\ : Odrv4
    port map (
            O => \N__39076\,
            I => eis_state_1
        );

    \I__8245\ : Odrv12
    port map (
            O => \N__39073\,
            I => eis_state_1
        );

    \I__8244\ : InMux
    port map (
            O => \N__39064\,
            I => \N__39058\
        );

    \I__8243\ : InMux
    port map (
            O => \N__39063\,
            I => \N__39058\
        );

    \I__8242\ : LocalMux
    port map (
            O => \N__39058\,
            I => \N__39054\
        );

    \I__8241\ : InMux
    port map (
            O => \N__39057\,
            I => \N__39051\
        );

    \I__8240\ : Span4Mux_h
    port map (
            O => \N__39054\,
            I => \N__39048\
        );

    \I__8239\ : LocalMux
    port map (
            O => \N__39051\,
            I => buf_dds0_7
        );

    \I__8238\ : Odrv4
    port map (
            O => \N__39048\,
            I => buf_dds0_7
        );

    \I__8237\ : InMux
    port map (
            O => \N__39043\,
            I => \N__39040\
        );

    \I__8236\ : LocalMux
    port map (
            O => \N__39040\,
            I => n8_adj_1541
        );

    \I__8235\ : CascadeMux
    port map (
            O => \N__39037\,
            I => \n8_adj_1541_cascade_\
        );

    \I__8234\ : CascadeMux
    port map (
            O => \N__39034\,
            I => \N__39031\
        );

    \I__8233\ : CascadeBuf
    port map (
            O => \N__39031\,
            I => \N__39028\
        );

    \I__8232\ : CascadeMux
    port map (
            O => \N__39028\,
            I => \N__39025\
        );

    \I__8231\ : CascadeBuf
    port map (
            O => \N__39025\,
            I => \N__39022\
        );

    \I__8230\ : CascadeMux
    port map (
            O => \N__39022\,
            I => \N__39019\
        );

    \I__8229\ : CascadeBuf
    port map (
            O => \N__39019\,
            I => \N__39016\
        );

    \I__8228\ : CascadeMux
    port map (
            O => \N__39016\,
            I => \N__39013\
        );

    \I__8227\ : CascadeBuf
    port map (
            O => \N__39013\,
            I => \N__39010\
        );

    \I__8226\ : CascadeMux
    port map (
            O => \N__39010\,
            I => \N__39007\
        );

    \I__8225\ : CascadeBuf
    port map (
            O => \N__39007\,
            I => \N__39004\
        );

    \I__8224\ : CascadeMux
    port map (
            O => \N__39004\,
            I => \N__39001\
        );

    \I__8223\ : CascadeBuf
    port map (
            O => \N__39001\,
            I => \N__38998\
        );

    \I__8222\ : CascadeMux
    port map (
            O => \N__38998\,
            I => \N__38995\
        );

    \I__8221\ : CascadeBuf
    port map (
            O => \N__38995\,
            I => \N__38992\
        );

    \I__8220\ : CascadeMux
    port map (
            O => \N__38992\,
            I => \N__38988\
        );

    \I__8219\ : CascadeMux
    port map (
            O => \N__38991\,
            I => \N__38985\
        );

    \I__8218\ : CascadeBuf
    port map (
            O => \N__38988\,
            I => \N__38982\
        );

    \I__8217\ : CascadeBuf
    port map (
            O => \N__38985\,
            I => \N__38979\
        );

    \I__8216\ : CascadeMux
    port map (
            O => \N__38982\,
            I => \N__38976\
        );

    \I__8215\ : CascadeMux
    port map (
            O => \N__38979\,
            I => \N__38973\
        );

    \I__8214\ : CascadeBuf
    port map (
            O => \N__38976\,
            I => \N__38970\
        );

    \I__8213\ : InMux
    port map (
            O => \N__38973\,
            I => \N__38967\
        );

    \I__8212\ : CascadeMux
    port map (
            O => \N__38970\,
            I => \N__38964\
        );

    \I__8211\ : LocalMux
    port map (
            O => \N__38967\,
            I => \N__38961\
        );

    \I__8210\ : InMux
    port map (
            O => \N__38964\,
            I => \N__38958\
        );

    \I__8209\ : Span4Mux_h
    port map (
            O => \N__38961\,
            I => \N__38955\
        );

    \I__8208\ : LocalMux
    port map (
            O => \N__38958\,
            I => \N__38952\
        );

    \I__8207\ : Span4Mux_h
    port map (
            O => \N__38955\,
            I => \N__38949\
        );

    \I__8206\ : Span12Mux_s10_v
    port map (
            O => \N__38952\,
            I => \N__38946\
        );

    \I__8205\ : Odrv4
    port map (
            O => \N__38949\,
            I => \data_index_9_N_212_4\
        );

    \I__8204\ : Odrv12
    port map (
            O => \N__38946\,
            I => \data_index_9_N_212_4\
        );

    \I__8203\ : InMux
    port map (
            O => \N__38941\,
            I => \N__38938\
        );

    \I__8202\ : LocalMux
    port map (
            O => \N__38938\,
            I => \N__38932\
        );

    \I__8201\ : InMux
    port map (
            O => \N__38937\,
            I => \N__38929\
        );

    \I__8200\ : InMux
    port map (
            O => \N__38936\,
            I => \N__38926\
        );

    \I__8199\ : InMux
    port map (
            O => \N__38935\,
            I => \N__38923\
        );

    \I__8198\ : Span4Mux_h
    port map (
            O => \N__38932\,
            I => \N__38920\
        );

    \I__8197\ : LocalMux
    port map (
            O => \N__38929\,
            I => \N__38917\
        );

    \I__8196\ : LocalMux
    port map (
            O => \N__38926\,
            I => \N__38914\
        );

    \I__8195\ : LocalMux
    port map (
            O => \N__38923\,
            I => \N__38907\
        );

    \I__8194\ : Span4Mux_v
    port map (
            O => \N__38920\,
            I => \N__38907\
        );

    \I__8193\ : Span4Mux_h
    port map (
            O => \N__38917\,
            I => \N__38907\
        );

    \I__8192\ : Odrv4
    port map (
            O => \N__38914\,
            I => eis_stop
        );

    \I__8191\ : Odrv4
    port map (
            O => \N__38907\,
            I => eis_stop
        );

    \I__8190\ : CascadeMux
    port map (
            O => \N__38902\,
            I => \n29_cascade_\
        );

    \I__8189\ : InMux
    port map (
            O => \N__38899\,
            I => \N__38894\
        );

    \I__8188\ : InMux
    port map (
            O => \N__38898\,
            I => \N__38891\
        );

    \I__8187\ : InMux
    port map (
            O => \N__38897\,
            I => \N__38888\
        );

    \I__8186\ : LocalMux
    port map (
            O => \N__38894\,
            I => \N__38885\
        );

    \I__8185\ : LocalMux
    port map (
            O => \N__38891\,
            I => \N__38882\
        );

    \I__8184\ : LocalMux
    port map (
            O => \N__38888\,
            I => \N__38879\
        );

    \I__8183\ : Span4Mux_h
    port map (
            O => \N__38885\,
            I => \N__38874\
        );

    \I__8182\ : Span4Mux_h
    port map (
            O => \N__38882\,
            I => \N__38874\
        );

    \I__8181\ : Odrv12
    port map (
            O => \N__38879\,
            I => n16_adj_1609
        );

    \I__8180\ : Odrv4
    port map (
            O => \N__38874\,
            I => n16_adj_1609
        );

    \I__8179\ : CascadeMux
    port map (
            O => \N__38869\,
            I => \N__38866\
        );

    \I__8178\ : InMux
    port map (
            O => \N__38866\,
            I => \N__38862\
        );

    \I__8177\ : InMux
    port map (
            O => \N__38865\,
            I => \N__38859\
        );

    \I__8176\ : LocalMux
    port map (
            O => \N__38862\,
            I => \N__38856\
        );

    \I__8175\ : LocalMux
    port map (
            O => \N__38859\,
            I => \N__38852\
        );

    \I__8174\ : Span4Mux_h
    port map (
            O => \N__38856\,
            I => \N__38849\
        );

    \I__8173\ : InMux
    port map (
            O => \N__38855\,
            I => \N__38846\
        );

    \I__8172\ : Span4Mux_v
    port map (
            O => \N__38852\,
            I => \N__38843\
        );

    \I__8171\ : Span4Mux_v
    port map (
            O => \N__38849\,
            I => \N__38838\
        );

    \I__8170\ : LocalMux
    port map (
            O => \N__38846\,
            I => \N__38838\
        );

    \I__8169\ : Odrv4
    port map (
            O => \N__38843\,
            I => n14_adj_1558
        );

    \I__8168\ : Odrv4
    port map (
            O => \N__38838\,
            I => n14_adj_1558
        );

    \I__8167\ : InMux
    port map (
            O => \N__38833\,
            I => \N__38830\
        );

    \I__8166\ : LocalMux
    port map (
            O => \N__38830\,
            I => \N__38827\
        );

    \I__8165\ : Span4Mux_h
    port map (
            O => \N__38827\,
            I => \N__38822\
        );

    \I__8164\ : InMux
    port map (
            O => \N__38826\,
            I => \N__38817\
        );

    \I__8163\ : InMux
    port map (
            O => \N__38825\,
            I => \N__38817\
        );

    \I__8162\ : Odrv4
    port map (
            O => \N__38822\,
            I => req_data_cnt_3
        );

    \I__8161\ : LocalMux
    port map (
            O => \N__38817\,
            I => req_data_cnt_3
        );

    \I__8160\ : InMux
    port map (
            O => \N__38812\,
            I => \N__38809\
        );

    \I__8159\ : LocalMux
    port map (
            O => \N__38809\,
            I => \N__38805\
        );

    \I__8158\ : InMux
    port map (
            O => \N__38808\,
            I => \N__38802\
        );

    \I__8157\ : Span4Mux_h
    port map (
            O => \N__38805\,
            I => \N__38799\
        );

    \I__8156\ : LocalMux
    port map (
            O => \N__38802\,
            I => acadc_skipcnt_12
        );

    \I__8155\ : Odrv4
    port map (
            O => \N__38799\,
            I => acadc_skipcnt_12
        );

    \I__8154\ : InMux
    port map (
            O => \N__38794\,
            I => \N__38791\
        );

    \I__8153\ : LocalMux
    port map (
            O => \N__38791\,
            I => \N__38787\
        );

    \I__8152\ : InMux
    port map (
            O => \N__38790\,
            I => \N__38784\
        );

    \I__8151\ : Span4Mux_h
    port map (
            O => \N__38787\,
            I => \N__38781\
        );

    \I__8150\ : LocalMux
    port map (
            O => \N__38784\,
            I => acadc_skipcnt_10
        );

    \I__8149\ : Odrv4
    port map (
            O => \N__38781\,
            I => acadc_skipcnt_10
        );

    \I__8148\ : InMux
    port map (
            O => \N__38776\,
            I => \N__38773\
        );

    \I__8147\ : LocalMux
    port map (
            O => \N__38773\,
            I => n21
        );

    \I__8146\ : CascadeMux
    port map (
            O => \N__38770\,
            I => \n9_adj_1408_cascade_\
        );

    \I__8145\ : InMux
    port map (
            O => \N__38767\,
            I => \N__38764\
        );

    \I__8144\ : LocalMux
    port map (
            O => \N__38764\,
            I => \N__38760\
        );

    \I__8143\ : CascadeMux
    port map (
            O => \N__38763\,
            I => \N__38756\
        );

    \I__8142\ : Span4Mux_v
    port map (
            O => \N__38760\,
            I => \N__38753\
        );

    \I__8141\ : CascadeMux
    port map (
            O => \N__38759\,
            I => \N__38750\
        );

    \I__8140\ : InMux
    port map (
            O => \N__38756\,
            I => \N__38747\
        );

    \I__8139\ : Span4Mux_h
    port map (
            O => \N__38753\,
            I => \N__38744\
        );

    \I__8138\ : InMux
    port map (
            O => \N__38750\,
            I => \N__38741\
        );

    \I__8137\ : LocalMux
    port map (
            O => \N__38747\,
            I => cmd_rdadctmp_14_adj_1429
        );

    \I__8136\ : Odrv4
    port map (
            O => \N__38744\,
            I => cmd_rdadctmp_14_adj_1429
        );

    \I__8135\ : LocalMux
    port map (
            O => \N__38741\,
            I => cmd_rdadctmp_14_adj_1429
        );

    \I__8134\ : CascadeMux
    port map (
            O => \N__38734\,
            I => \N__38726\
        );

    \I__8133\ : CascadeMux
    port map (
            O => \N__38733\,
            I => \N__38723\
        );

    \I__8132\ : CascadeMux
    port map (
            O => \N__38732\,
            I => \N__38720\
        );

    \I__8131\ : CascadeMux
    port map (
            O => \N__38731\,
            I => \N__38716\
        );

    \I__8130\ : CascadeMux
    port map (
            O => \N__38730\,
            I => \N__38713\
        );

    \I__8129\ : CascadeMux
    port map (
            O => \N__38729\,
            I => \N__38709\
        );

    \I__8128\ : InMux
    port map (
            O => \N__38726\,
            I => \N__38706\
        );

    \I__8127\ : InMux
    port map (
            O => \N__38723\,
            I => \N__38703\
        );

    \I__8126\ : InMux
    port map (
            O => \N__38720\,
            I => \N__38700\
        );

    \I__8125\ : InMux
    port map (
            O => \N__38719\,
            I => \N__38697\
        );

    \I__8124\ : InMux
    port map (
            O => \N__38716\,
            I => \N__38694\
        );

    \I__8123\ : InMux
    port map (
            O => \N__38713\,
            I => \N__38691\
        );

    \I__8122\ : InMux
    port map (
            O => \N__38712\,
            I => \N__38688\
        );

    \I__8121\ : InMux
    port map (
            O => \N__38709\,
            I => \N__38685\
        );

    \I__8120\ : LocalMux
    port map (
            O => \N__38706\,
            I => \N__38682\
        );

    \I__8119\ : LocalMux
    port map (
            O => \N__38703\,
            I => \N__38679\
        );

    \I__8118\ : LocalMux
    port map (
            O => \N__38700\,
            I => \N__38676\
        );

    \I__8117\ : LocalMux
    port map (
            O => \N__38697\,
            I => \N__38673\
        );

    \I__8116\ : LocalMux
    port map (
            O => \N__38694\,
            I => \N__38668\
        );

    \I__8115\ : LocalMux
    port map (
            O => \N__38691\,
            I => \N__38668\
        );

    \I__8114\ : LocalMux
    port map (
            O => \N__38688\,
            I => \N__38665\
        );

    \I__8113\ : LocalMux
    port map (
            O => \N__38685\,
            I => \N__38662\
        );

    \I__8112\ : Span4Mux_v
    port map (
            O => \N__38682\,
            I => \N__38659\
        );

    \I__8111\ : Span4Mux_v
    port map (
            O => \N__38679\,
            I => \N__38654\
        );

    \I__8110\ : Span4Mux_h
    port map (
            O => \N__38676\,
            I => \N__38654\
        );

    \I__8109\ : Span4Mux_h
    port map (
            O => \N__38673\,
            I => \N__38651\
        );

    \I__8108\ : Span4Mux_v
    port map (
            O => \N__38668\,
            I => \N__38645\
        );

    \I__8107\ : Span4Mux_h
    port map (
            O => \N__38665\,
            I => \N__38645\
        );

    \I__8106\ : Span12Mux_v
    port map (
            O => \N__38662\,
            I => \N__38640\
        );

    \I__8105\ : Sp12to4
    port map (
            O => \N__38659\,
            I => \N__38640\
        );

    \I__8104\ : Span4Mux_v
    port map (
            O => \N__38654\,
            I => \N__38635\
        );

    \I__8103\ : Span4Mux_h
    port map (
            O => \N__38651\,
            I => \N__38635\
        );

    \I__8102\ : InMux
    port map (
            O => \N__38650\,
            I => \N__38632\
        );

    \I__8101\ : Odrv4
    port map (
            O => \N__38645\,
            I => comm_buf_0_2
        );

    \I__8100\ : Odrv12
    port map (
            O => \N__38640\,
            I => comm_buf_0_2
        );

    \I__8099\ : Odrv4
    port map (
            O => \N__38635\,
            I => comm_buf_0_2
        );

    \I__8098\ : LocalMux
    port map (
            O => \N__38632\,
            I => comm_buf_0_2
        );

    \I__8097\ : InMux
    port map (
            O => \N__38623\,
            I => \N__38620\
        );

    \I__8096\ : LocalMux
    port map (
            O => \N__38620\,
            I => \N__38617\
        );

    \I__8095\ : Span4Mux_h
    port map (
            O => \N__38617\,
            I => \N__38614\
        );

    \I__8094\ : Span4Mux_h
    port map (
            O => \N__38614\,
            I => \N__38609\
        );

    \I__8093\ : CascadeMux
    port map (
            O => \N__38613\,
            I => \N__38606\
        );

    \I__8092\ : InMux
    port map (
            O => \N__38612\,
            I => \N__38603\
        );

    \I__8091\ : Span4Mux_v
    port map (
            O => \N__38609\,
            I => \N__38600\
        );

    \I__8090\ : InMux
    port map (
            O => \N__38606\,
            I => \N__38597\
        );

    \I__8089\ : LocalMux
    port map (
            O => \N__38603\,
            I => \acadc_skipCount_10\
        );

    \I__8088\ : Odrv4
    port map (
            O => \N__38600\,
            I => \acadc_skipCount_10\
        );

    \I__8087\ : LocalMux
    port map (
            O => \N__38597\,
            I => \acadc_skipCount_10\
        );

    \I__8086\ : InMux
    port map (
            O => \N__38590\,
            I => \N__38587\
        );

    \I__8085\ : LocalMux
    port map (
            O => \N__38587\,
            I => \N__38584\
        );

    \I__8084\ : Odrv4
    port map (
            O => \N__38584\,
            I => n14_adj_1550
        );

    \I__8083\ : CEMux
    port map (
            O => \N__38581\,
            I => \N__38577\
        );

    \I__8082\ : CEMux
    port map (
            O => \N__38580\,
            I => \N__38574\
        );

    \I__8081\ : LocalMux
    port map (
            O => \N__38577\,
            I => \N__38571\
        );

    \I__8080\ : LocalMux
    port map (
            O => \N__38574\,
            I => \N__38568\
        );

    \I__8079\ : Span4Mux_h
    port map (
            O => \N__38571\,
            I => \N__38565\
        );

    \I__8078\ : Span4Mux_h
    port map (
            O => \N__38568\,
            I => \N__38562\
        );

    \I__8077\ : Odrv4
    port map (
            O => \N__38565\,
            I => n12254
        );

    \I__8076\ : Odrv4
    port map (
            O => \N__38562\,
            I => n12254
        );

    \I__8075\ : CEMux
    port map (
            O => \N__38557\,
            I => \N__38554\
        );

    \I__8074\ : LocalMux
    port map (
            O => \N__38554\,
            I => \N__38551\
        );

    \I__8073\ : Span4Mux_v
    port map (
            O => \N__38551\,
            I => \N__38547\
        );

    \I__8072\ : CEMux
    port map (
            O => \N__38550\,
            I => \N__38541\
        );

    \I__8071\ : Span4Mux_h
    port map (
            O => \N__38547\,
            I => \N__38537\
        );

    \I__8070\ : CEMux
    port map (
            O => \N__38546\,
            I => \N__38534\
        );

    \I__8069\ : CEMux
    port map (
            O => \N__38545\,
            I => \N__38530\
        );

    \I__8068\ : CEMux
    port map (
            O => \N__38544\,
            I => \N__38527\
        );

    \I__8067\ : LocalMux
    port map (
            O => \N__38541\,
            I => \N__38524\
        );

    \I__8066\ : CEMux
    port map (
            O => \N__38540\,
            I => \N__38520\
        );

    \I__8065\ : Span4Mux_h
    port map (
            O => \N__38537\,
            I => \N__38515\
        );

    \I__8064\ : LocalMux
    port map (
            O => \N__38534\,
            I => \N__38515\
        );

    \I__8063\ : CEMux
    port map (
            O => \N__38533\,
            I => \N__38512\
        );

    \I__8062\ : LocalMux
    port map (
            O => \N__38530\,
            I => \N__38509\
        );

    \I__8061\ : LocalMux
    port map (
            O => \N__38527\,
            I => \N__38504\
        );

    \I__8060\ : Span4Mux_v
    port map (
            O => \N__38524\,
            I => \N__38504\
        );

    \I__8059\ : CEMux
    port map (
            O => \N__38523\,
            I => \N__38501\
        );

    \I__8058\ : LocalMux
    port map (
            O => \N__38520\,
            I => \N__38498\
        );

    \I__8057\ : Span4Mux_h
    port map (
            O => \N__38515\,
            I => \N__38494\
        );

    \I__8056\ : LocalMux
    port map (
            O => \N__38512\,
            I => \N__38487\
        );

    \I__8055\ : Span4Mux_v
    port map (
            O => \N__38509\,
            I => \N__38487\
        );

    \I__8054\ : Span4Mux_h
    port map (
            O => \N__38504\,
            I => \N__38487\
        );

    \I__8053\ : LocalMux
    port map (
            O => \N__38501\,
            I => \N__38482\
        );

    \I__8052\ : Span4Mux_v
    port map (
            O => \N__38498\,
            I => \N__38482\
        );

    \I__8051\ : InMux
    port map (
            O => \N__38497\,
            I => \N__38479\
        );

    \I__8050\ : Odrv4
    port map (
            O => \N__38494\,
            I => n12007
        );

    \I__8049\ : Odrv4
    port map (
            O => \N__38487\,
            I => n12007
        );

    \I__8048\ : Odrv4
    port map (
            O => \N__38482\,
            I => n12007
        );

    \I__8047\ : LocalMux
    port map (
            O => \N__38479\,
            I => n12007
        );

    \I__8046\ : InMux
    port map (
            O => \N__38470\,
            I => \N__38466\
        );

    \I__8045\ : InMux
    port map (
            O => \N__38469\,
            I => \N__38463\
        );

    \I__8044\ : LocalMux
    port map (
            O => \N__38466\,
            I => \N__38460\
        );

    \I__8043\ : LocalMux
    port map (
            O => \N__38463\,
            I => \N__38457\
        );

    \I__8042\ : Span4Mux_v
    port map (
            O => \N__38460\,
            I => \N__38454\
        );

    \I__8041\ : Span4Mux_h
    port map (
            O => \N__38457\,
            I => \N__38451\
        );

    \I__8040\ : Span4Mux_h
    port map (
            O => \N__38454\,
            I => \N__38446\
        );

    \I__8039\ : Span4Mux_v
    port map (
            O => \N__38451\,
            I => \N__38446\
        );

    \I__8038\ : Odrv4
    port map (
            O => \N__38446\,
            I => n14_adj_1527
        );

    \I__8037\ : InMux
    port map (
            O => \N__38443\,
            I => \N__38439\
        );

    \I__8036\ : InMux
    port map (
            O => \N__38442\,
            I => \N__38436\
        );

    \I__8035\ : LocalMux
    port map (
            O => \N__38439\,
            I => \N__38433\
        );

    \I__8034\ : LocalMux
    port map (
            O => \N__38436\,
            I => \N__38430\
        );

    \I__8033\ : Span4Mux_h
    port map (
            O => \N__38433\,
            I => \N__38427\
        );

    \I__8032\ : Odrv12
    port map (
            O => \N__38430\,
            I => n14_adj_1529
        );

    \I__8031\ : Odrv4
    port map (
            O => \N__38427\,
            I => n14_adj_1529
        );

    \I__8030\ : InMux
    port map (
            O => \N__38422\,
            I => \N__38419\
        );

    \I__8029\ : LocalMux
    port map (
            O => \N__38419\,
            I => \N__38414\
        );

    \I__8028\ : CascadeMux
    port map (
            O => \N__38418\,
            I => \N__38411\
        );

    \I__8027\ : InMux
    port map (
            O => \N__38417\,
            I => \N__38408\
        );

    \I__8026\ : Span4Mux_h
    port map (
            O => \N__38414\,
            I => \N__38405\
        );

    \I__8025\ : InMux
    port map (
            O => \N__38411\,
            I => \N__38402\
        );

    \I__8024\ : LocalMux
    port map (
            O => \N__38408\,
            I => req_data_cnt_5
        );

    \I__8023\ : Odrv4
    port map (
            O => \N__38405\,
            I => req_data_cnt_5
        );

    \I__8022\ : LocalMux
    port map (
            O => \N__38402\,
            I => req_data_cnt_5
        );

    \I__8021\ : InMux
    port map (
            O => \N__38395\,
            I => \N__38391\
        );

    \I__8020\ : CascadeMux
    port map (
            O => \N__38394\,
            I => \N__38387\
        );

    \I__8019\ : LocalMux
    port map (
            O => \N__38391\,
            I => \N__38384\
        );

    \I__8018\ : InMux
    port map (
            O => \N__38390\,
            I => \N__38379\
        );

    \I__8017\ : InMux
    port map (
            O => \N__38387\,
            I => \N__38379\
        );

    \I__8016\ : Odrv4
    port map (
            O => \N__38384\,
            I => req_data_cnt_4
        );

    \I__8015\ : LocalMux
    port map (
            O => \N__38379\,
            I => req_data_cnt_4
        );

    \I__8014\ : InMux
    port map (
            O => \N__38374\,
            I => \N__38369\
        );

    \I__8013\ : InMux
    port map (
            O => \N__38373\,
            I => \N__38364\
        );

    \I__8012\ : InMux
    port map (
            O => \N__38372\,
            I => \N__38364\
        );

    \I__8011\ : LocalMux
    port map (
            O => \N__38369\,
            I => req_data_cnt_1
        );

    \I__8010\ : LocalMux
    port map (
            O => \N__38364\,
            I => req_data_cnt_1
        );

    \I__8009\ : InMux
    port map (
            O => \N__38359\,
            I => \N__38356\
        );

    \I__8008\ : LocalMux
    port map (
            O => \N__38356\,
            I => n20_adj_1496
        );

    \I__8007\ : CascadeMux
    port map (
            O => \N__38353\,
            I => \n18_adj_1553_cascade_\
        );

    \I__8006\ : SRMux
    port map (
            O => \N__38350\,
            I => \N__38347\
        );

    \I__8005\ : LocalMux
    port map (
            O => \N__38347\,
            I => \N__38343\
        );

    \I__8004\ : SRMux
    port map (
            O => \N__38346\,
            I => \N__38340\
        );

    \I__8003\ : Span4Mux_h
    port map (
            O => \N__38343\,
            I => \N__38337\
        );

    \I__8002\ : LocalMux
    port map (
            O => \N__38340\,
            I => \N__38334\
        );

    \I__8001\ : Odrv4
    port map (
            O => \N__38337\,
            I => n14749
        );

    \I__8000\ : Odrv12
    port map (
            O => \N__38334\,
            I => n14749
        );

    \I__7999\ : InMux
    port map (
            O => \N__38329\,
            I => \N__38326\
        );

    \I__7998\ : LocalMux
    port map (
            O => \N__38326\,
            I => \N__38323\
        );

    \I__7997\ : Span4Mux_v
    port map (
            O => \N__38323\,
            I => \N__38320\
        );

    \I__7996\ : Span4Mux_h
    port map (
            O => \N__38320\,
            I => \N__38316\
        );

    \I__7995\ : InMux
    port map (
            O => \N__38319\,
            I => \N__38313\
        );

    \I__7994\ : Odrv4
    port map (
            O => \N__38316\,
            I => buf_adcdata_vdc_5
        );

    \I__7993\ : LocalMux
    port map (
            O => \N__38313\,
            I => buf_adcdata_vdc_5
        );

    \I__7992\ : InMux
    port map (
            O => \N__38308\,
            I => \N__38305\
        );

    \I__7991\ : LocalMux
    port map (
            O => \N__38305\,
            I => \N__38300\
        );

    \I__7990\ : CascadeMux
    port map (
            O => \N__38304\,
            I => \N__38297\
        );

    \I__7989\ : InMux
    port map (
            O => \N__38303\,
            I => \N__38294\
        );

    \I__7988\ : Span4Mux_v
    port map (
            O => \N__38300\,
            I => \N__38291\
        );

    \I__7987\ : InMux
    port map (
            O => \N__38297\,
            I => \N__38288\
        );

    \I__7986\ : LocalMux
    port map (
            O => \N__38294\,
            I => \N__38285\
        );

    \I__7985\ : Span4Mux_h
    port map (
            O => \N__38291\,
            I => \N__38282\
        );

    \I__7984\ : LocalMux
    port map (
            O => \N__38288\,
            I => buf_adcdata_vac_5
        );

    \I__7983\ : Odrv4
    port map (
            O => \N__38285\,
            I => buf_adcdata_vac_5
        );

    \I__7982\ : Odrv4
    port map (
            O => \N__38282\,
            I => buf_adcdata_vac_5
        );

    \I__7981\ : InMux
    port map (
            O => \N__38275\,
            I => \N__38272\
        );

    \I__7980\ : LocalMux
    port map (
            O => \N__38272\,
            I => n19_adj_1598
        );

    \I__7979\ : InMux
    port map (
            O => \N__38269\,
            I => \N__38266\
        );

    \I__7978\ : LocalMux
    port map (
            O => \N__38266\,
            I => comm_buf_2_5
        );

    \I__7977\ : CascadeMux
    port map (
            O => \N__38263\,
            I => \N__38260\
        );

    \I__7976\ : InMux
    port map (
            O => \N__38260\,
            I => \N__38256\
        );

    \I__7975\ : InMux
    port map (
            O => \N__38259\,
            I => \N__38253\
        );

    \I__7974\ : LocalMux
    port map (
            O => \N__38256\,
            I => \N__38250\
        );

    \I__7973\ : LocalMux
    port map (
            O => \N__38253\,
            I => \N__38245\
        );

    \I__7972\ : Span4Mux_h
    port map (
            O => \N__38250\,
            I => \N__38245\
        );

    \I__7971\ : Odrv4
    port map (
            O => \N__38245\,
            I => comm_buf_6_5
        );

    \I__7970\ : InMux
    port map (
            O => \N__38242\,
            I => \N__38239\
        );

    \I__7969\ : LocalMux
    port map (
            O => \N__38239\,
            I => \N__38236\
        );

    \I__7968\ : Span4Mux_h
    port map (
            O => \N__38236\,
            I => \N__38233\
        );

    \I__7967\ : Span4Mux_h
    port map (
            O => \N__38233\,
            I => \N__38230\
        );

    \I__7966\ : Span4Mux_v
    port map (
            O => \N__38230\,
            I => \N__38227\
        );

    \I__7965\ : Odrv4
    port map (
            O => \N__38227\,
            I => comm_buf_4_5
        );

    \I__7964\ : CascadeMux
    port map (
            O => \N__38224\,
            I => \n22123_cascade_\
        );

    \I__7963\ : InMux
    port map (
            O => \N__38221\,
            I => \N__38218\
        );

    \I__7962\ : LocalMux
    port map (
            O => \N__38218\,
            I => \N__38215\
        );

    \I__7961\ : Span4Mux_h
    port map (
            O => \N__38215\,
            I => \N__38212\
        );

    \I__7960\ : Odrv4
    port map (
            O => \N__38212\,
            I => n22126
        );

    \I__7959\ : InMux
    port map (
            O => \N__38209\,
            I => \N__38203\
        );

    \I__7958\ : InMux
    port map (
            O => \N__38208\,
            I => \N__38203\
        );

    \I__7957\ : LocalMux
    port map (
            O => \N__38203\,
            I => \N__38198\
        );

    \I__7956\ : InMux
    port map (
            O => \N__38202\,
            I => \N__38193\
        );

    \I__7955\ : InMux
    port map (
            O => \N__38201\,
            I => \N__38193\
        );

    \I__7954\ : Span4Mux_h
    port map (
            O => \N__38198\,
            I => \N__38190\
        );

    \I__7953\ : LocalMux
    port map (
            O => \N__38193\,
            I => n20602
        );

    \I__7952\ : Odrv4
    port map (
            O => \N__38190\,
            I => n20602
        );

    \I__7951\ : IoInMux
    port map (
            O => \N__38185\,
            I => \N__38182\
        );

    \I__7950\ : LocalMux
    port map (
            O => \N__38182\,
            I => \N__38179\
        );

    \I__7949\ : IoSpan4Mux
    port map (
            O => \N__38179\,
            I => \N__38176\
        );

    \I__7948\ : IoSpan4Mux
    port map (
            O => \N__38176\,
            I => \N__38172\
        );

    \I__7947\ : InMux
    port map (
            O => \N__38175\,
            I => \N__38169\
        );

    \I__7946\ : Span4Mux_s3_v
    port map (
            O => \N__38172\,
            I => \N__38166\
        );

    \I__7945\ : LocalMux
    port map (
            O => \N__38169\,
            I => \N__38163\
        );

    \I__7944\ : Span4Mux_v
    port map (
            O => \N__38166\,
            I => \N__38159\
        );

    \I__7943\ : Span4Mux_h
    port map (
            O => \N__38163\,
            I => \N__38156\
        );

    \I__7942\ : InMux
    port map (
            O => \N__38162\,
            I => \N__38153\
        );

    \I__7941\ : Span4Mux_v
    port map (
            O => \N__38159\,
            I => \N__38148\
        );

    \I__7940\ : Span4Mux_h
    port map (
            O => \N__38156\,
            I => \N__38148\
        );

    \I__7939\ : LocalMux
    port map (
            O => \N__38153\,
            I => \SELIRNG0\
        );

    \I__7938\ : Odrv4
    port map (
            O => \N__38148\,
            I => \SELIRNG0\
        );

    \I__7937\ : InMux
    port map (
            O => \N__38143\,
            I => \N__38140\
        );

    \I__7936\ : LocalMux
    port map (
            O => \N__38140\,
            I => \N__38137\
        );

    \I__7935\ : Odrv12
    port map (
            O => \N__38137\,
            I => n14_adj_1552
        );

    \I__7934\ : CascadeMux
    port map (
            O => \N__38134\,
            I => \n14_adj_1552_cascade_\
        );

    \I__7933\ : InMux
    port map (
            O => \N__38131\,
            I => \N__38128\
        );

    \I__7932\ : LocalMux
    port map (
            O => \N__38128\,
            I => n16_adj_1570
        );

    \I__7931\ : CascadeMux
    port map (
            O => \N__38125\,
            I => \n12080_cascade_\
        );

    \I__7930\ : InMux
    port map (
            O => \N__38122\,
            I => \N__38119\
        );

    \I__7929\ : LocalMux
    port map (
            O => \N__38119\,
            I => \N__38116\
        );

    \I__7928\ : Odrv4
    port map (
            O => \N__38116\,
            I => comm_buf_4_0
        );

    \I__7927\ : InMux
    port map (
            O => \N__38113\,
            I => \N__38110\
        );

    \I__7926\ : LocalMux
    port map (
            O => \N__38110\,
            I => \N__38107\
        );

    \I__7925\ : Odrv4
    port map (
            O => \N__38107\,
            I => n22132
        );

    \I__7924\ : CEMux
    port map (
            O => \N__38104\,
            I => \N__38101\
        );

    \I__7923\ : LocalMux
    port map (
            O => \N__38101\,
            I => \N__38098\
        );

    \I__7922\ : Odrv4
    port map (
            O => \N__38098\,
            I => n12206
        );

    \I__7921\ : CascadeMux
    port map (
            O => \N__38095\,
            I => \n12206_cascade_\
        );

    \I__7920\ : SRMux
    port map (
            O => \N__38092\,
            I => \N__38089\
        );

    \I__7919\ : LocalMux
    port map (
            O => \N__38089\,
            I => \N__38086\
        );

    \I__7918\ : Odrv4
    port map (
            O => \N__38086\,
            I => n14770
        );

    \I__7917\ : InMux
    port map (
            O => \N__38083\,
            I => \N__38080\
        );

    \I__7916\ : LocalMux
    port map (
            O => \N__38080\,
            I => \N__38077\
        );

    \I__7915\ : Span4Mux_v
    port map (
            O => \N__38077\,
            I => \N__38073\
        );

    \I__7914\ : CascadeMux
    port map (
            O => \N__38076\,
            I => \N__38070\
        );

    \I__7913\ : Span4Mux_h
    port map (
            O => \N__38073\,
            I => \N__38067\
        );

    \I__7912\ : InMux
    port map (
            O => \N__38070\,
            I => \N__38064\
        );

    \I__7911\ : Span4Mux_v
    port map (
            O => \N__38067\,
            I => \N__38061\
        );

    \I__7910\ : LocalMux
    port map (
            O => \N__38064\,
            I => comm_buf_6_0
        );

    \I__7909\ : Odrv4
    port map (
            O => \N__38061\,
            I => comm_buf_6_0
        );

    \I__7908\ : CascadeMux
    port map (
            O => \N__38056\,
            I => \N__38053\
        );

    \I__7907\ : InMux
    port map (
            O => \N__38053\,
            I => \N__38050\
        );

    \I__7906\ : LocalMux
    port map (
            O => \N__38050\,
            I => comm_buf_2_0
        );

    \I__7905\ : InMux
    port map (
            O => \N__38047\,
            I => \N__38044\
        );

    \I__7904\ : LocalMux
    port map (
            O => \N__38044\,
            I => n22129
        );

    \I__7903\ : InMux
    port map (
            O => \N__38041\,
            I => \N__38038\
        );

    \I__7902\ : LocalMux
    port map (
            O => \N__38038\,
            I => \N__38035\
        );

    \I__7901\ : Span12Mux_v
    port map (
            O => \N__38035\,
            I => \N__38032\
        );

    \I__7900\ : Odrv12
    port map (
            O => \N__38032\,
            I => buf_data_iac_5
        );

    \I__7899\ : CascadeMux
    port map (
            O => \N__38029\,
            I => \n22_adj_1599_cascade_\
        );

    \I__7898\ : CascadeMux
    port map (
            O => \N__38026\,
            I => \n30_adj_1600_cascade_\
        );

    \I__7897\ : CascadeMux
    port map (
            O => \N__38023\,
            I => \N__38019\
        );

    \I__7896\ : InMux
    port map (
            O => \N__38022\,
            I => \N__38013\
        );

    \I__7895\ : InMux
    port map (
            O => \N__38019\,
            I => \N__38010\
        );

    \I__7894\ : InMux
    port map (
            O => \N__38018\,
            I => \N__38007\
        );

    \I__7893\ : InMux
    port map (
            O => \N__38017\,
            I => \N__38004\
        );

    \I__7892\ : CascadeMux
    port map (
            O => \N__38016\,
            I => \N__38001\
        );

    \I__7891\ : LocalMux
    port map (
            O => \N__38013\,
            I => \N__37996\
        );

    \I__7890\ : LocalMux
    port map (
            O => \N__38010\,
            I => \N__37996\
        );

    \I__7889\ : LocalMux
    port map (
            O => \N__38007\,
            I => \N__37991\
        );

    \I__7888\ : LocalMux
    port map (
            O => \N__38004\,
            I => \N__37988\
        );

    \I__7887\ : InMux
    port map (
            O => \N__38001\,
            I => \N__37985\
        );

    \I__7886\ : Span4Mux_v
    port map (
            O => \N__37996\,
            I => \N__37982\
        );

    \I__7885\ : InMux
    port map (
            O => \N__37995\,
            I => \N__37978\
        );

    \I__7884\ : CascadeMux
    port map (
            O => \N__37994\,
            I => \N__37975\
        );

    \I__7883\ : Span4Mux_v
    port map (
            O => \N__37991\,
            I => \N__37972\
        );

    \I__7882\ : Span4Mux_v
    port map (
            O => \N__37988\,
            I => \N__37969\
        );

    \I__7881\ : LocalMux
    port map (
            O => \N__37985\,
            I => \N__37966\
        );

    \I__7880\ : Span4Mux_h
    port map (
            O => \N__37982\,
            I => \N__37963\
        );

    \I__7879\ : InMux
    port map (
            O => \N__37981\,
            I => \N__37960\
        );

    \I__7878\ : LocalMux
    port map (
            O => \N__37978\,
            I => \N__37957\
        );

    \I__7877\ : InMux
    port map (
            O => \N__37975\,
            I => \N__37954\
        );

    \I__7876\ : Span4Mux_v
    port map (
            O => \N__37972\,
            I => \N__37948\
        );

    \I__7875\ : Span4Mux_v
    port map (
            O => \N__37969\,
            I => \N__37948\
        );

    \I__7874\ : Span4Mux_h
    port map (
            O => \N__37966\,
            I => \N__37941\
        );

    \I__7873\ : Span4Mux_h
    port map (
            O => \N__37963\,
            I => \N__37941\
        );

    \I__7872\ : LocalMux
    port map (
            O => \N__37960\,
            I => \N__37941\
        );

    \I__7871\ : Span4Mux_h
    port map (
            O => \N__37957\,
            I => \N__37938\
        );

    \I__7870\ : LocalMux
    port map (
            O => \N__37954\,
            I => \N__37935\
        );

    \I__7869\ : InMux
    port map (
            O => \N__37953\,
            I => \N__37932\
        );

    \I__7868\ : Odrv4
    port map (
            O => \N__37948\,
            I => comm_rx_buf_5
        );

    \I__7867\ : Odrv4
    port map (
            O => \N__37941\,
            I => comm_rx_buf_5
        );

    \I__7866\ : Odrv4
    port map (
            O => \N__37938\,
            I => comm_rx_buf_5
        );

    \I__7865\ : Odrv4
    port map (
            O => \N__37935\,
            I => comm_rx_buf_5
        );

    \I__7864\ : LocalMux
    port map (
            O => \N__37932\,
            I => comm_rx_buf_5
        );

    \I__7863\ : CEMux
    port map (
            O => \N__37921\,
            I => \N__37917\
        );

    \I__7862\ : CEMux
    port map (
            O => \N__37920\,
            I => \N__37914\
        );

    \I__7861\ : LocalMux
    port map (
            O => \N__37917\,
            I => n12080
        );

    \I__7860\ : LocalMux
    port map (
            O => \N__37914\,
            I => n12080
        );

    \I__7859\ : CascadeMux
    port map (
            O => \N__37909\,
            I => \n11839_cascade_\
        );

    \I__7858\ : InMux
    port map (
            O => \N__37906\,
            I => \N__37902\
        );

    \I__7857\ : InMux
    port map (
            O => \N__37905\,
            I => \N__37899\
        );

    \I__7856\ : LocalMux
    port map (
            O => \N__37902\,
            I => n9222
        );

    \I__7855\ : LocalMux
    port map (
            O => \N__37899\,
            I => n9222
        );

    \I__7854\ : CascadeMux
    port map (
            O => \N__37894\,
            I => \n9222_cascade_\
        );

    \I__7853\ : CascadeMux
    port map (
            O => \N__37891\,
            I => \n24_adj_1579_cascade_\
        );

    \I__7852\ : CascadeMux
    port map (
            O => \N__37888\,
            I => \n21079_cascade_\
        );

    \I__7851\ : InMux
    port map (
            O => \N__37885\,
            I => \N__37879\
        );

    \I__7850\ : InMux
    port map (
            O => \N__37884\,
            I => \N__37879\
        );

    \I__7849\ : LocalMux
    port map (
            O => \N__37879\,
            I => \N__37865\
        );

    \I__7848\ : InMux
    port map (
            O => \N__37878\,
            I => \N__37860\
        );

    \I__7847\ : InMux
    port map (
            O => \N__37877\,
            I => \N__37860\
        );

    \I__7846\ : InMux
    port map (
            O => \N__37876\,
            I => \N__37851\
        );

    \I__7845\ : InMux
    port map (
            O => \N__37875\,
            I => \N__37851\
        );

    \I__7844\ : InMux
    port map (
            O => \N__37874\,
            I => \N__37851\
        );

    \I__7843\ : InMux
    port map (
            O => \N__37873\,
            I => \N__37851\
        );

    \I__7842\ : InMux
    port map (
            O => \N__37872\,
            I => \N__37848\
        );

    \I__7841\ : InMux
    port map (
            O => \N__37871\,
            I => \N__37845\
        );

    \I__7840\ : InMux
    port map (
            O => \N__37870\,
            I => \N__37841\
        );

    \I__7839\ : InMux
    port map (
            O => \N__37869\,
            I => \N__37827\
        );

    \I__7838\ : InMux
    port map (
            O => \N__37868\,
            I => \N__37827\
        );

    \I__7837\ : Span4Mux_v
    port map (
            O => \N__37865\,
            I => \N__37824\
        );

    \I__7836\ : LocalMux
    port map (
            O => \N__37860\,
            I => \N__37817\
        );

    \I__7835\ : LocalMux
    port map (
            O => \N__37851\,
            I => \N__37817\
        );

    \I__7834\ : LocalMux
    port map (
            O => \N__37848\,
            I => \N__37817\
        );

    \I__7833\ : LocalMux
    port map (
            O => \N__37845\,
            I => \N__37814\
        );

    \I__7832\ : InMux
    port map (
            O => \N__37844\,
            I => \N__37811\
        );

    \I__7831\ : LocalMux
    port map (
            O => \N__37841\,
            I => \N__37808\
        );

    \I__7830\ : InMux
    port map (
            O => \N__37840\,
            I => \N__37801\
        );

    \I__7829\ : InMux
    port map (
            O => \N__37839\,
            I => \N__37801\
        );

    \I__7828\ : InMux
    port map (
            O => \N__37838\,
            I => \N__37801\
        );

    \I__7827\ : InMux
    port map (
            O => \N__37837\,
            I => \N__37788\
        );

    \I__7826\ : InMux
    port map (
            O => \N__37836\,
            I => \N__37788\
        );

    \I__7825\ : InMux
    port map (
            O => \N__37835\,
            I => \N__37788\
        );

    \I__7824\ : InMux
    port map (
            O => \N__37834\,
            I => \N__37788\
        );

    \I__7823\ : InMux
    port map (
            O => \N__37833\,
            I => \N__37788\
        );

    \I__7822\ : InMux
    port map (
            O => \N__37832\,
            I => \N__37788\
        );

    \I__7821\ : LocalMux
    port map (
            O => \N__37827\,
            I => \N__37776\
        );

    \I__7820\ : Span4Mux_h
    port map (
            O => \N__37824\,
            I => \N__37771\
        );

    \I__7819\ : Span4Mux_v
    port map (
            O => \N__37817\,
            I => \N__37771\
        );

    \I__7818\ : Span12Mux_h
    port map (
            O => \N__37814\,
            I => \N__37766\
        );

    \I__7817\ : LocalMux
    port map (
            O => \N__37811\,
            I => \N__37766\
        );

    \I__7816\ : Span4Mux_v
    port map (
            O => \N__37808\,
            I => \N__37759\
        );

    \I__7815\ : LocalMux
    port map (
            O => \N__37801\,
            I => \N__37759\
        );

    \I__7814\ : LocalMux
    port map (
            O => \N__37788\,
            I => \N__37759\
        );

    \I__7813\ : InMux
    port map (
            O => \N__37787\,
            I => \N__37752\
        );

    \I__7812\ : InMux
    port map (
            O => \N__37786\,
            I => \N__37752\
        );

    \I__7811\ : InMux
    port map (
            O => \N__37785\,
            I => \N__37752\
        );

    \I__7810\ : InMux
    port map (
            O => \N__37784\,
            I => \N__37739\
        );

    \I__7809\ : InMux
    port map (
            O => \N__37783\,
            I => \N__37739\
        );

    \I__7808\ : InMux
    port map (
            O => \N__37782\,
            I => \N__37739\
        );

    \I__7807\ : InMux
    port map (
            O => \N__37781\,
            I => \N__37739\
        );

    \I__7806\ : InMux
    port map (
            O => \N__37780\,
            I => \N__37739\
        );

    \I__7805\ : InMux
    port map (
            O => \N__37779\,
            I => \N__37739\
        );

    \I__7804\ : Odrv4
    port map (
            O => \N__37776\,
            I => n12643
        );

    \I__7803\ : Odrv4
    port map (
            O => \N__37771\,
            I => n12643
        );

    \I__7802\ : Odrv12
    port map (
            O => \N__37766\,
            I => n12643
        );

    \I__7801\ : Odrv4
    port map (
            O => \N__37759\,
            I => n12643
        );

    \I__7800\ : LocalMux
    port map (
            O => \N__37752\,
            I => n12643
        );

    \I__7799\ : LocalMux
    port map (
            O => \N__37739\,
            I => n12643
        );

    \I__7798\ : InMux
    port map (
            O => \N__37726\,
            I => \N__37723\
        );

    \I__7797\ : LocalMux
    port map (
            O => \N__37723\,
            I => \N__37720\
        );

    \I__7796\ : Span4Mux_v
    port map (
            O => \N__37720\,
            I => \N__37715\
        );

    \I__7795\ : InMux
    port map (
            O => \N__37719\,
            I => \N__37712\
        );

    \I__7794\ : InMux
    port map (
            O => \N__37718\,
            I => \N__37709\
        );

    \I__7793\ : Odrv4
    port map (
            O => \N__37715\,
            I => \comm_spi.n22644\
        );

    \I__7792\ : LocalMux
    port map (
            O => \N__37712\,
            I => \comm_spi.n22644\
        );

    \I__7791\ : LocalMux
    port map (
            O => \N__37709\,
            I => \comm_spi.n22644\
        );

    \I__7790\ : SRMux
    port map (
            O => \N__37702\,
            I => \N__37699\
        );

    \I__7789\ : LocalMux
    port map (
            O => \N__37699\,
            I => \N__37696\
        );

    \I__7788\ : Odrv4
    port map (
            O => \N__37696\,
            I => \comm_spi.data_tx_7__N_778\
        );

    \I__7787\ : InMux
    port map (
            O => \N__37693\,
            I => \N__37690\
        );

    \I__7786\ : LocalMux
    port map (
            O => \N__37690\,
            I => \N__37686\
        );

    \I__7785\ : InMux
    port map (
            O => \N__37689\,
            I => \N__37683\
        );

    \I__7784\ : Odrv4
    port map (
            O => \N__37686\,
            I => \comm_spi.n14608\
        );

    \I__7783\ : LocalMux
    port map (
            O => \N__37683\,
            I => \comm_spi.n14608\
        );

    \I__7782\ : SRMux
    port map (
            O => \N__37678\,
            I => \N__37675\
        );

    \I__7781\ : LocalMux
    port map (
            O => \N__37675\,
            I => \N__37672\
        );

    \I__7780\ : Span4Mux_h
    port map (
            O => \N__37672\,
            I => \N__37669\
        );

    \I__7779\ : Odrv4
    port map (
            O => \N__37669\,
            I => \comm_spi.data_tx_7__N_781\
        );

    \I__7778\ : InMux
    port map (
            O => \N__37666\,
            I => \N__37663\
        );

    \I__7777\ : LocalMux
    port map (
            O => \N__37663\,
            I => \N__37659\
        );

    \I__7776\ : InMux
    port map (
            O => \N__37662\,
            I => \N__37656\
        );

    \I__7775\ : Span4Mux_v
    port map (
            O => \N__37659\,
            I => \N__37653\
        );

    \I__7774\ : LocalMux
    port map (
            O => \N__37656\,
            I => \N__37650\
        );

    \I__7773\ : Odrv4
    port map (
            O => \N__37653\,
            I => \comm_spi.n14607\
        );

    \I__7772\ : Odrv4
    port map (
            O => \N__37650\,
            I => \comm_spi.n14607\
        );

    \I__7771\ : SRMux
    port map (
            O => \N__37645\,
            I => \N__37642\
        );

    \I__7770\ : LocalMux
    port map (
            O => \N__37642\,
            I => \N__37639\
        );

    \I__7769\ : Sp12to4
    port map (
            O => \N__37639\,
            I => \N__37636\
        );

    \I__7768\ : Odrv12
    port map (
            O => \N__37636\,
            I => \comm_spi.data_tx_7__N_763\
        );

    \I__7767\ : InMux
    port map (
            O => \N__37633\,
            I => \N__37630\
        );

    \I__7766\ : LocalMux
    port map (
            O => \N__37630\,
            I => \N__37625\
        );

    \I__7765\ : InMux
    port map (
            O => \N__37629\,
            I => \N__37620\
        );

    \I__7764\ : InMux
    port map (
            O => \N__37628\,
            I => \N__37620\
        );

    \I__7763\ : Span4Mux_h
    port map (
            O => \N__37625\,
            I => \N__37617\
        );

    \I__7762\ : LocalMux
    port map (
            O => \N__37620\,
            I => \N__37614\
        );

    \I__7761\ : Span4Mux_h
    port map (
            O => \N__37617\,
            I => \N__37609\
        );

    \I__7760\ : Span4Mux_v
    port map (
            O => \N__37614\,
            I => \N__37609\
        );

    \I__7759\ : Odrv4
    port map (
            O => \N__37609\,
            I => comm_tx_buf_3
        );

    \I__7758\ : InMux
    port map (
            O => \N__37606\,
            I => \N__37599\
        );

    \I__7757\ : CascadeMux
    port map (
            O => \N__37605\,
            I => \N__37596\
        );

    \I__7756\ : InMux
    port map (
            O => \N__37604\,
            I => \N__37590\
        );

    \I__7755\ : InMux
    port map (
            O => \N__37603\,
            I => \N__37587\
        );

    \I__7754\ : InMux
    port map (
            O => \N__37602\,
            I => \N__37584\
        );

    \I__7753\ : LocalMux
    port map (
            O => \N__37599\,
            I => \N__37577\
        );

    \I__7752\ : InMux
    port map (
            O => \N__37596\,
            I => \N__37574\
        );

    \I__7751\ : InMux
    port map (
            O => \N__37595\,
            I => \N__37569\
        );

    \I__7750\ : InMux
    port map (
            O => \N__37594\,
            I => \N__37569\
        );

    \I__7749\ : InMux
    port map (
            O => \N__37593\,
            I => \N__37566\
        );

    \I__7748\ : LocalMux
    port map (
            O => \N__37590\,
            I => \N__37559\
        );

    \I__7747\ : LocalMux
    port map (
            O => \N__37587\,
            I => \N__37559\
        );

    \I__7746\ : LocalMux
    port map (
            O => \N__37584\,
            I => \N__37559\
        );

    \I__7745\ : InMux
    port map (
            O => \N__37583\,
            I => \N__37550\
        );

    \I__7744\ : InMux
    port map (
            O => \N__37582\,
            I => \N__37550\
        );

    \I__7743\ : InMux
    port map (
            O => \N__37581\,
            I => \N__37550\
        );

    \I__7742\ : InMux
    port map (
            O => \N__37580\,
            I => \N__37550\
        );

    \I__7741\ : Span4Mux_h
    port map (
            O => \N__37577\,
            I => \N__37547\
        );

    \I__7740\ : LocalMux
    port map (
            O => \N__37574\,
            I => \N__37540\
        );

    \I__7739\ : LocalMux
    port map (
            O => \N__37569\,
            I => \N__37540\
        );

    \I__7738\ : LocalMux
    port map (
            O => \N__37566\,
            I => \N__37540\
        );

    \I__7737\ : Span4Mux_v
    port map (
            O => \N__37559\,
            I => \N__37537\
        );

    \I__7736\ : LocalMux
    port map (
            O => \N__37550\,
            I => eis_state_0
        );

    \I__7735\ : Odrv4
    port map (
            O => \N__37547\,
            I => eis_state_0
        );

    \I__7734\ : Odrv12
    port map (
            O => \N__37540\,
            I => eis_state_0
        );

    \I__7733\ : Odrv4
    port map (
            O => \N__37537\,
            I => eis_state_0
        );

    \I__7732\ : InMux
    port map (
            O => \N__37528\,
            I => \N__37525\
        );

    \I__7731\ : LocalMux
    port map (
            O => \N__37525\,
            I => \N__37522\
        );

    \I__7730\ : Span4Mux_v
    port map (
            O => \N__37522\,
            I => \N__37519\
        );

    \I__7729\ : Odrv4
    port map (
            O => \N__37519\,
            I => n21067
        );

    \I__7728\ : InMux
    port map (
            O => \N__37516\,
            I => \N__37512\
        );

    \I__7727\ : InMux
    port map (
            O => \N__37515\,
            I => \N__37509\
        );

    \I__7726\ : LocalMux
    port map (
            O => \N__37512\,
            I => \N__37506\
        );

    \I__7725\ : LocalMux
    port map (
            O => \N__37509\,
            I => n10508
        );

    \I__7724\ : Odrv12
    port map (
            O => \N__37506\,
            I => n10508
        );

    \I__7723\ : InMux
    port map (
            O => \N__37501\,
            I => \ADC_VDC.genclk.n19439\
        );

    \I__7722\ : CascadeMux
    port map (
            O => \N__37498\,
            I => \N__37494\
        );

    \I__7721\ : InMux
    port map (
            O => \N__37497\,
            I => \N__37491\
        );

    \I__7720\ : InMux
    port map (
            O => \N__37494\,
            I => \N__37488\
        );

    \I__7719\ : LocalMux
    port map (
            O => \N__37491\,
            I => \ADC_VDC.genclk.t0on_15\
        );

    \I__7718\ : LocalMux
    port map (
            O => \N__37488\,
            I => \ADC_VDC.genclk.t0on_15\
        );

    \I__7717\ : CEMux
    port map (
            O => \N__37483\,
            I => \N__37479\
        );

    \I__7716\ : CEMux
    port map (
            O => \N__37482\,
            I => \N__37476\
        );

    \I__7715\ : LocalMux
    port map (
            O => \N__37479\,
            I => \N__37473\
        );

    \I__7714\ : LocalMux
    port map (
            O => \N__37476\,
            I => \N__37470\
        );

    \I__7713\ : Span4Mux_v
    port map (
            O => \N__37473\,
            I => \N__37467\
        );

    \I__7712\ : Span4Mux_v
    port map (
            O => \N__37470\,
            I => \N__37464\
        );

    \I__7711\ : Span4Mux_h
    port map (
            O => \N__37467\,
            I => \N__37459\
        );

    \I__7710\ : Span4Mux_h
    port map (
            O => \N__37464\,
            I => \N__37459\
        );

    \I__7709\ : Odrv4
    port map (
            O => \N__37459\,
            I => \ADC_VDC.genclk.div_state_1__N_1266\
        );

    \I__7708\ : SRMux
    port map (
            O => \N__37456\,
            I => \N__37453\
        );

    \I__7707\ : LocalMux
    port map (
            O => \N__37453\,
            I => \N__37449\
        );

    \I__7706\ : SRMux
    port map (
            O => \N__37452\,
            I => \N__37446\
        );

    \I__7705\ : Span4Mux_v
    port map (
            O => \N__37449\,
            I => \N__37439\
        );

    \I__7704\ : LocalMux
    port map (
            O => \N__37446\,
            I => \N__37439\
        );

    \I__7703\ : SRMux
    port map (
            O => \N__37445\,
            I => \N__37436\
        );

    \I__7702\ : SRMux
    port map (
            O => \N__37444\,
            I => \N__37433\
        );

    \I__7701\ : Odrv4
    port map (
            O => \N__37439\,
            I => \ADC_VDC.genclk.n14695\
        );

    \I__7700\ : LocalMux
    port map (
            O => \N__37436\,
            I => \ADC_VDC.genclk.n14695\
        );

    \I__7699\ : LocalMux
    port map (
            O => \N__37433\,
            I => \ADC_VDC.genclk.n14695\
        );

    \I__7698\ : InMux
    port map (
            O => \N__37426\,
            I => \N__37421\
        );

    \I__7697\ : InMux
    port map (
            O => \N__37425\,
            I => \N__37418\
        );

    \I__7696\ : InMux
    port map (
            O => \N__37424\,
            I => \N__37415\
        );

    \I__7695\ : LocalMux
    port map (
            O => \N__37421\,
            I => \N__37412\
        );

    \I__7694\ : LocalMux
    port map (
            O => \N__37418\,
            I => \N__37407\
        );

    \I__7693\ : LocalMux
    port map (
            O => \N__37415\,
            I => \N__37407\
        );

    \I__7692\ : Span4Mux_v
    port map (
            O => \N__37412\,
            I => \N__37404\
        );

    \I__7691\ : Span4Mux_h
    port map (
            O => \N__37407\,
            I => \N__37401\
        );

    \I__7690\ : Odrv4
    port map (
            O => \N__37404\,
            I => \comm_spi.n14585\
        );

    \I__7689\ : Odrv4
    port map (
            O => \N__37401\,
            I => \comm_spi.n14585\
        );

    \I__7688\ : CascadeMux
    port map (
            O => \N__37396\,
            I => \N__37392\
        );

    \I__7687\ : InMux
    port map (
            O => \N__37395\,
            I => \N__37388\
        );

    \I__7686\ : InMux
    port map (
            O => \N__37392\,
            I => \N__37383\
        );

    \I__7685\ : InMux
    port map (
            O => \N__37391\,
            I => \N__37383\
        );

    \I__7684\ : LocalMux
    port map (
            O => \N__37388\,
            I => comm_tx_buf_7
        );

    \I__7683\ : LocalMux
    port map (
            O => \N__37383\,
            I => comm_tx_buf_7
        );

    \I__7682\ : InMux
    port map (
            O => \N__37378\,
            I => \N__37369\
        );

    \I__7681\ : InMux
    port map (
            O => \N__37377\,
            I => \N__37369\
        );

    \I__7680\ : InMux
    port map (
            O => \N__37376\,
            I => \N__37369\
        );

    \I__7679\ : LocalMux
    port map (
            O => \N__37369\,
            I => \N__37366\
        );

    \I__7678\ : Odrv4
    port map (
            O => \N__37366\,
            I => comm_tx_buf_2
        );

    \I__7677\ : SRMux
    port map (
            O => \N__37363\,
            I => \N__37360\
        );

    \I__7676\ : LocalMux
    port map (
            O => \N__37360\,
            I => \comm_spi.imosi_N_744\
        );

    \I__7675\ : InMux
    port map (
            O => \N__37357\,
            I => \N__37350\
        );

    \I__7674\ : InMux
    port map (
            O => \N__37356\,
            I => \N__37350\
        );

    \I__7673\ : InMux
    port map (
            O => \N__37355\,
            I => \N__37347\
        );

    \I__7672\ : LocalMux
    port map (
            O => \N__37350\,
            I => \N__37343\
        );

    \I__7671\ : LocalMux
    port map (
            O => \N__37347\,
            I => \N__37339\
        );

    \I__7670\ : InMux
    port map (
            O => \N__37346\,
            I => \N__37336\
        );

    \I__7669\ : Span4Mux_v
    port map (
            O => \N__37343\,
            I => \N__37333\
        );

    \I__7668\ : InMux
    port map (
            O => \N__37342\,
            I => \N__37330\
        );

    \I__7667\ : Span4Mux_h
    port map (
            O => \N__37339\,
            I => \N__37325\
        );

    \I__7666\ : LocalMux
    port map (
            O => \N__37336\,
            I => \N__37325\
        );

    \I__7665\ : Sp12to4
    port map (
            O => \N__37333\,
            I => \N__37322\
        );

    \I__7664\ : LocalMux
    port map (
            O => \N__37330\,
            I => \N__37317\
        );

    \I__7663\ : Sp12to4
    port map (
            O => \N__37325\,
            I => \N__37317\
        );

    \I__7662\ : Span12Mux_h
    port map (
            O => \N__37322\,
            I => \N__37314\
        );

    \I__7661\ : Span12Mux_v
    port map (
            O => \N__37317\,
            I => \N__37311\
        );

    \I__7660\ : Span12Mux_v
    port map (
            O => \N__37314\,
            I => \N__37308\
        );

    \I__7659\ : Span12Mux_h
    port map (
            O => \N__37311\,
            I => \N__37305\
        );

    \I__7658\ : Odrv12
    port map (
            O => \N__37308\,
            I => \ICE_SPI_MOSI\
        );

    \I__7657\ : Odrv12
    port map (
            O => \N__37305\,
            I => \ICE_SPI_MOSI\
        );

    \I__7656\ : SRMux
    port map (
            O => \N__37300\,
            I => \N__37297\
        );

    \I__7655\ : LocalMux
    port map (
            O => \N__37297\,
            I => \N__37294\
        );

    \I__7654\ : Span4Mux_h
    port map (
            O => \N__37294\,
            I => \N__37291\
        );

    \I__7653\ : Odrv4
    port map (
            O => \N__37291\,
            I => \comm_spi.imosi_N_745\
        );

    \I__7652\ : CascadeMux
    port map (
            O => \N__37288\,
            I => \N__37284\
        );

    \I__7651\ : InMux
    port map (
            O => \N__37287\,
            I => \N__37281\
        );

    \I__7650\ : InMux
    port map (
            O => \N__37284\,
            I => \N__37278\
        );

    \I__7649\ : LocalMux
    port map (
            O => \N__37281\,
            I => \ADC_VDC.genclk.t0on_7\
        );

    \I__7648\ : LocalMux
    port map (
            O => \N__37278\,
            I => \ADC_VDC.genclk.t0on_7\
        );

    \I__7647\ : InMux
    port map (
            O => \N__37273\,
            I => \ADC_VDC.genclk.n19431\
        );

    \I__7646\ : InMux
    port map (
            O => \N__37270\,
            I => \N__37266\
        );

    \I__7645\ : InMux
    port map (
            O => \N__37269\,
            I => \N__37263\
        );

    \I__7644\ : LocalMux
    port map (
            O => \N__37266\,
            I => \ADC_VDC.genclk.t0on_8\
        );

    \I__7643\ : LocalMux
    port map (
            O => \N__37263\,
            I => \ADC_VDC.genclk.t0on_8\
        );

    \I__7642\ : InMux
    port map (
            O => \N__37258\,
            I => \bfn_15_4_0_\
        );

    \I__7641\ : CascadeMux
    port map (
            O => \N__37255\,
            I => \N__37252\
        );

    \I__7640\ : InMux
    port map (
            O => \N__37252\,
            I => \N__37248\
        );

    \I__7639\ : InMux
    port map (
            O => \N__37251\,
            I => \N__37245\
        );

    \I__7638\ : LocalMux
    port map (
            O => \N__37248\,
            I => \ADC_VDC.genclk.t0on_9\
        );

    \I__7637\ : LocalMux
    port map (
            O => \N__37245\,
            I => \ADC_VDC.genclk.t0on_9\
        );

    \I__7636\ : InMux
    port map (
            O => \N__37240\,
            I => \ADC_VDC.genclk.n19433\
        );

    \I__7635\ : InMux
    port map (
            O => \N__37237\,
            I => \N__37233\
        );

    \I__7634\ : InMux
    port map (
            O => \N__37236\,
            I => \N__37230\
        );

    \I__7633\ : LocalMux
    port map (
            O => \N__37233\,
            I => \ADC_VDC.genclk.t0on_10\
        );

    \I__7632\ : LocalMux
    port map (
            O => \N__37230\,
            I => \ADC_VDC.genclk.t0on_10\
        );

    \I__7631\ : InMux
    port map (
            O => \N__37225\,
            I => \ADC_VDC.genclk.n19434\
        );

    \I__7630\ : CascadeMux
    port map (
            O => \N__37222\,
            I => \N__37219\
        );

    \I__7629\ : InMux
    port map (
            O => \N__37219\,
            I => \N__37215\
        );

    \I__7628\ : InMux
    port map (
            O => \N__37218\,
            I => \N__37212\
        );

    \I__7627\ : LocalMux
    port map (
            O => \N__37215\,
            I => \ADC_VDC.genclk.t0on_11\
        );

    \I__7626\ : LocalMux
    port map (
            O => \N__37212\,
            I => \ADC_VDC.genclk.t0on_11\
        );

    \I__7625\ : InMux
    port map (
            O => \N__37207\,
            I => \ADC_VDC.genclk.n19435\
        );

    \I__7624\ : InMux
    port map (
            O => \N__37204\,
            I => \N__37200\
        );

    \I__7623\ : InMux
    port map (
            O => \N__37203\,
            I => \N__37197\
        );

    \I__7622\ : LocalMux
    port map (
            O => \N__37200\,
            I => \ADC_VDC.genclk.t0on_12\
        );

    \I__7621\ : LocalMux
    port map (
            O => \N__37197\,
            I => \ADC_VDC.genclk.t0on_12\
        );

    \I__7620\ : InMux
    port map (
            O => \N__37192\,
            I => \ADC_VDC.genclk.n19436\
        );

    \I__7619\ : CascadeMux
    port map (
            O => \N__37189\,
            I => \N__37186\
        );

    \I__7618\ : InMux
    port map (
            O => \N__37186\,
            I => \N__37182\
        );

    \I__7617\ : InMux
    port map (
            O => \N__37185\,
            I => \N__37179\
        );

    \I__7616\ : LocalMux
    port map (
            O => \N__37182\,
            I => \ADC_VDC.genclk.t0on_13\
        );

    \I__7615\ : LocalMux
    port map (
            O => \N__37179\,
            I => \ADC_VDC.genclk.t0on_13\
        );

    \I__7614\ : InMux
    port map (
            O => \N__37174\,
            I => \ADC_VDC.genclk.n19437\
        );

    \I__7613\ : InMux
    port map (
            O => \N__37171\,
            I => \N__37167\
        );

    \I__7612\ : InMux
    port map (
            O => \N__37170\,
            I => \N__37164\
        );

    \I__7611\ : LocalMux
    port map (
            O => \N__37167\,
            I => \ADC_VDC.genclk.t0on_14\
        );

    \I__7610\ : LocalMux
    port map (
            O => \N__37164\,
            I => \ADC_VDC.genclk.t0on_14\
        );

    \I__7609\ : InMux
    port map (
            O => \N__37159\,
            I => \ADC_VDC.genclk.n19438\
        );

    \I__7608\ : CascadeMux
    port map (
            O => \N__37156\,
            I => \N__37153\
        );

    \I__7607\ : InMux
    port map (
            O => \N__37153\,
            I => \N__37150\
        );

    \I__7606\ : LocalMux
    port map (
            O => \N__37150\,
            I => \SIG_DDS.tmp_buf_4\
        );

    \I__7605\ : CascadeMux
    port map (
            O => \N__37147\,
            I => \N__37144\
        );

    \I__7604\ : InMux
    port map (
            O => \N__37144\,
            I => \N__37141\
        );

    \I__7603\ : LocalMux
    port map (
            O => \N__37141\,
            I => \SIG_DDS.tmp_buf_5\
        );

    \I__7602\ : InMux
    port map (
            O => \N__37138\,
            I => \N__37135\
        );

    \I__7601\ : LocalMux
    port map (
            O => \N__37135\,
            I => \N__37132\
        );

    \I__7600\ : Span4Mux_h
    port map (
            O => \N__37132\,
            I => \N__37129\
        );

    \I__7599\ : Odrv4
    port map (
            O => \N__37129\,
            I => \SIG_DDS.tmp_buf_6\
        );

    \I__7598\ : InMux
    port map (
            O => \N__37126\,
            I => \N__37122\
        );

    \I__7597\ : InMux
    port map (
            O => \N__37125\,
            I => \N__37119\
        );

    \I__7596\ : LocalMux
    port map (
            O => \N__37122\,
            I => \ADC_VDC.genclk.t0on_0\
        );

    \I__7595\ : LocalMux
    port map (
            O => \N__37119\,
            I => \ADC_VDC.genclk.t0on_0\
        );

    \I__7594\ : InMux
    port map (
            O => \N__37114\,
            I => \bfn_15_3_0_\
        );

    \I__7593\ : InMux
    port map (
            O => \N__37111\,
            I => \N__37107\
        );

    \I__7592\ : InMux
    port map (
            O => \N__37110\,
            I => \N__37104\
        );

    \I__7591\ : LocalMux
    port map (
            O => \N__37107\,
            I => \ADC_VDC.genclk.t0on_1\
        );

    \I__7590\ : LocalMux
    port map (
            O => \N__37104\,
            I => \ADC_VDC.genclk.t0on_1\
        );

    \I__7589\ : InMux
    port map (
            O => \N__37099\,
            I => \ADC_VDC.genclk.n19425\
        );

    \I__7588\ : CascadeMux
    port map (
            O => \N__37096\,
            I => \N__37093\
        );

    \I__7587\ : InMux
    port map (
            O => \N__37093\,
            I => \N__37089\
        );

    \I__7586\ : InMux
    port map (
            O => \N__37092\,
            I => \N__37086\
        );

    \I__7585\ : LocalMux
    port map (
            O => \N__37089\,
            I => \ADC_VDC.genclk.t0on_2\
        );

    \I__7584\ : LocalMux
    port map (
            O => \N__37086\,
            I => \ADC_VDC.genclk.t0on_2\
        );

    \I__7583\ : InMux
    port map (
            O => \N__37081\,
            I => \ADC_VDC.genclk.n19426\
        );

    \I__7582\ : InMux
    port map (
            O => \N__37078\,
            I => \N__37074\
        );

    \I__7581\ : InMux
    port map (
            O => \N__37077\,
            I => \N__37071\
        );

    \I__7580\ : LocalMux
    port map (
            O => \N__37074\,
            I => \ADC_VDC.genclk.t0on_3\
        );

    \I__7579\ : LocalMux
    port map (
            O => \N__37071\,
            I => \ADC_VDC.genclk.t0on_3\
        );

    \I__7578\ : InMux
    port map (
            O => \N__37066\,
            I => \ADC_VDC.genclk.n19427\
        );

    \I__7577\ : CascadeMux
    port map (
            O => \N__37063\,
            I => \N__37059\
        );

    \I__7576\ : CascadeMux
    port map (
            O => \N__37062\,
            I => \N__37056\
        );

    \I__7575\ : InMux
    port map (
            O => \N__37059\,
            I => \N__37053\
        );

    \I__7574\ : InMux
    port map (
            O => \N__37056\,
            I => \N__37050\
        );

    \I__7573\ : LocalMux
    port map (
            O => \N__37053\,
            I => \N__37047\
        );

    \I__7572\ : LocalMux
    port map (
            O => \N__37050\,
            I => \ADC_VDC.genclk.t0on_4\
        );

    \I__7571\ : Odrv4
    port map (
            O => \N__37047\,
            I => \ADC_VDC.genclk.t0on_4\
        );

    \I__7570\ : InMux
    port map (
            O => \N__37042\,
            I => \ADC_VDC.genclk.n19428\
        );

    \I__7569\ : CascadeMux
    port map (
            O => \N__37039\,
            I => \N__37035\
        );

    \I__7568\ : InMux
    port map (
            O => \N__37038\,
            I => \N__37032\
        );

    \I__7567\ : InMux
    port map (
            O => \N__37035\,
            I => \N__37029\
        );

    \I__7566\ : LocalMux
    port map (
            O => \N__37032\,
            I => \ADC_VDC.genclk.t0on_5\
        );

    \I__7565\ : LocalMux
    port map (
            O => \N__37029\,
            I => \ADC_VDC.genclk.t0on_5\
        );

    \I__7564\ : InMux
    port map (
            O => \N__37024\,
            I => \ADC_VDC.genclk.n19429\
        );

    \I__7563\ : CascadeMux
    port map (
            O => \N__37021\,
            I => \N__37018\
        );

    \I__7562\ : InMux
    port map (
            O => \N__37018\,
            I => \N__37014\
        );

    \I__7561\ : InMux
    port map (
            O => \N__37017\,
            I => \N__37011\
        );

    \I__7560\ : LocalMux
    port map (
            O => \N__37014\,
            I => \ADC_VDC.genclk.t0on_6\
        );

    \I__7559\ : LocalMux
    port map (
            O => \N__37011\,
            I => \ADC_VDC.genclk.t0on_6\
        );

    \I__7558\ : InMux
    port map (
            O => \N__37006\,
            I => \ADC_VDC.genclk.n19430\
        );

    \I__7557\ : CascadeMux
    port map (
            O => \N__37003\,
            I => \N__37000\
        );

    \I__7556\ : InMux
    port map (
            O => \N__37000\,
            I => \N__36997\
        );

    \I__7555\ : LocalMux
    port map (
            O => \N__36997\,
            I => \N__36994\
        );

    \I__7554\ : Odrv4
    port map (
            O => \N__36994\,
            I => n20949
        );

    \I__7553\ : InMux
    port map (
            O => \N__36991\,
            I => \N__36988\
        );

    \I__7552\ : LocalMux
    port map (
            O => \N__36988\,
            I => n26_adj_1623
        );

    \I__7551\ : CascadeMux
    port map (
            O => \N__36985\,
            I => \n21949_cascade_\
        );

    \I__7550\ : InMux
    port map (
            O => \N__36982\,
            I => \N__36979\
        );

    \I__7549\ : LocalMux
    port map (
            O => \N__36979\,
            I => \N__36974\
        );

    \I__7548\ : InMux
    port map (
            O => \N__36978\,
            I => \N__36969\
        );

    \I__7547\ : InMux
    port map (
            O => \N__36977\,
            I => \N__36969\
        );

    \I__7546\ : Odrv4
    port map (
            O => \N__36974\,
            I => \acadc_skipCount_7\
        );

    \I__7545\ : LocalMux
    port map (
            O => \N__36969\,
            I => \acadc_skipCount_7\
        );

    \I__7544\ : InMux
    port map (
            O => \N__36964\,
            I => \N__36961\
        );

    \I__7543\ : LocalMux
    port map (
            O => \N__36961\,
            I => \N__36958\
        );

    \I__7542\ : Span4Mux_h
    port map (
            O => \N__36958\,
            I => \N__36955\
        );

    \I__7541\ : Odrv4
    port map (
            O => \N__36955\,
            I => n21964
        );

    \I__7540\ : CascadeMux
    port map (
            O => \N__36952\,
            I => \n21952_cascade_\
        );

    \I__7539\ : InMux
    port map (
            O => \N__36949\,
            I => \N__36944\
        );

    \I__7538\ : InMux
    port map (
            O => \N__36948\,
            I => \N__36941\
        );

    \I__7537\ : InMux
    port map (
            O => \N__36947\,
            I => \N__36938\
        );

    \I__7536\ : LocalMux
    port map (
            O => \N__36944\,
            I => \N__36935\
        );

    \I__7535\ : LocalMux
    port map (
            O => \N__36941\,
            I => \N__36932\
        );

    \I__7534\ : LocalMux
    port map (
            O => \N__36938\,
            I => \acadc_skipCount_4\
        );

    \I__7533\ : Odrv4
    port map (
            O => \N__36935\,
            I => \acadc_skipCount_4\
        );

    \I__7532\ : Odrv4
    port map (
            O => \N__36932\,
            I => \acadc_skipCount_4\
        );

    \I__7531\ : InMux
    port map (
            O => \N__36925\,
            I => \N__36922\
        );

    \I__7530\ : LocalMux
    port map (
            O => \N__36922\,
            I => \N__36917\
        );

    \I__7529\ : CascadeMux
    port map (
            O => \N__36921\,
            I => \N__36914\
        );

    \I__7528\ : InMux
    port map (
            O => \N__36920\,
            I => \N__36911\
        );

    \I__7527\ : Span12Mux_h
    port map (
            O => \N__36917\,
            I => \N__36908\
        );

    \I__7526\ : InMux
    port map (
            O => \N__36914\,
            I => \N__36905\
        );

    \I__7525\ : LocalMux
    port map (
            O => \N__36911\,
            I => \acadc_skipCount_9\
        );

    \I__7524\ : Odrv12
    port map (
            O => \N__36908\,
            I => \acadc_skipCount_9\
        );

    \I__7523\ : LocalMux
    port map (
            O => \N__36905\,
            I => \acadc_skipCount_9\
        );

    \I__7522\ : InMux
    port map (
            O => \N__36898\,
            I => \N__36891\
        );

    \I__7521\ : CascadeMux
    port map (
            O => \N__36897\,
            I => \N__36888\
        );

    \I__7520\ : InMux
    port map (
            O => \N__36896\,
            I => \N__36885\
        );

    \I__7519\ : InMux
    port map (
            O => \N__36895\,
            I => \N__36882\
        );

    \I__7518\ : InMux
    port map (
            O => \N__36894\,
            I => \N__36877\
        );

    \I__7517\ : LocalMux
    port map (
            O => \N__36891\,
            I => \N__36874\
        );

    \I__7516\ : InMux
    port map (
            O => \N__36888\,
            I => \N__36871\
        );

    \I__7515\ : LocalMux
    port map (
            O => \N__36885\,
            I => \N__36868\
        );

    \I__7514\ : LocalMux
    port map (
            O => \N__36882\,
            I => \N__36865\
        );

    \I__7513\ : InMux
    port map (
            O => \N__36881\,
            I => \N__36862\
        );

    \I__7512\ : CascadeMux
    port map (
            O => \N__36880\,
            I => \N__36859\
        );

    \I__7511\ : LocalMux
    port map (
            O => \N__36877\,
            I => \N__36855\
        );

    \I__7510\ : Span4Mux_v
    port map (
            O => \N__36874\,
            I => \N__36850\
        );

    \I__7509\ : LocalMux
    port map (
            O => \N__36871\,
            I => \N__36850\
        );

    \I__7508\ : Span4Mux_h
    port map (
            O => \N__36868\,
            I => \N__36843\
        );

    \I__7507\ : Span4Mux_v
    port map (
            O => \N__36865\,
            I => \N__36843\
        );

    \I__7506\ : LocalMux
    port map (
            O => \N__36862\,
            I => \N__36843\
        );

    \I__7505\ : InMux
    port map (
            O => \N__36859\,
            I => \N__36840\
        );

    \I__7504\ : CascadeMux
    port map (
            O => \N__36858\,
            I => \N__36837\
        );

    \I__7503\ : Span12Mux_v
    port map (
            O => \N__36855\,
            I => \N__36834\
        );

    \I__7502\ : Span4Mux_h
    port map (
            O => \N__36850\,
            I => \N__36831\
        );

    \I__7501\ : Span4Mux_h
    port map (
            O => \N__36843\,
            I => \N__36826\
        );

    \I__7500\ : LocalMux
    port map (
            O => \N__36840\,
            I => \N__36826\
        );

    \I__7499\ : InMux
    port map (
            O => \N__36837\,
            I => \N__36823\
        );

    \I__7498\ : Odrv12
    port map (
            O => \N__36834\,
            I => comm_rx_buf_7
        );

    \I__7497\ : Odrv4
    port map (
            O => \N__36831\,
            I => comm_rx_buf_7
        );

    \I__7496\ : Odrv4
    port map (
            O => \N__36826\,
            I => comm_rx_buf_7
        );

    \I__7495\ : LocalMux
    port map (
            O => \N__36823\,
            I => comm_rx_buf_7
        );

    \I__7494\ : InMux
    port map (
            O => \N__36814\,
            I => \N__36811\
        );

    \I__7493\ : LocalMux
    port map (
            O => \N__36811\,
            I => n30_adj_1624
        );

    \I__7492\ : SRMux
    port map (
            O => \N__36808\,
            I => \N__36804\
        );

    \I__7491\ : SRMux
    port map (
            O => \N__36807\,
            I => \N__36800\
        );

    \I__7490\ : LocalMux
    port map (
            O => \N__36804\,
            I => \N__36797\
        );

    \I__7489\ : SRMux
    port map (
            O => \N__36803\,
            I => \N__36792\
        );

    \I__7488\ : LocalMux
    port map (
            O => \N__36800\,
            I => \N__36787\
        );

    \I__7487\ : Span4Mux_h
    port map (
            O => \N__36797\,
            I => \N__36784\
        );

    \I__7486\ : SRMux
    port map (
            O => \N__36796\,
            I => \N__36781\
        );

    \I__7485\ : SRMux
    port map (
            O => \N__36795\,
            I => \N__36777\
        );

    \I__7484\ : LocalMux
    port map (
            O => \N__36792\,
            I => \N__36774\
        );

    \I__7483\ : SRMux
    port map (
            O => \N__36791\,
            I => \N__36771\
        );

    \I__7482\ : SRMux
    port map (
            O => \N__36790\,
            I => \N__36768\
        );

    \I__7481\ : Span4Mux_v
    port map (
            O => \N__36787\,
            I => \N__36761\
        );

    \I__7480\ : Span4Mux_h
    port map (
            O => \N__36784\,
            I => \N__36761\
        );

    \I__7479\ : LocalMux
    port map (
            O => \N__36781\,
            I => \N__36761\
        );

    \I__7478\ : SRMux
    port map (
            O => \N__36780\,
            I => \N__36758\
        );

    \I__7477\ : LocalMux
    port map (
            O => \N__36777\,
            I => \N__36755\
        );

    \I__7476\ : Span4Mux_v
    port map (
            O => \N__36774\,
            I => \N__36752\
        );

    \I__7475\ : LocalMux
    port map (
            O => \N__36771\,
            I => \N__36749\
        );

    \I__7474\ : LocalMux
    port map (
            O => \N__36768\,
            I => \N__36742\
        );

    \I__7473\ : Span4Mux_v
    port map (
            O => \N__36761\,
            I => \N__36742\
        );

    \I__7472\ : LocalMux
    port map (
            O => \N__36758\,
            I => \N__36742\
        );

    \I__7471\ : Span4Mux_h
    port map (
            O => \N__36755\,
            I => \N__36737\
        );

    \I__7470\ : Span4Mux_h
    port map (
            O => \N__36752\,
            I => \N__36737\
        );

    \I__7469\ : Span4Mux_h
    port map (
            O => \N__36749\,
            I => \N__36734\
        );

    \I__7468\ : Sp12to4
    port map (
            O => \N__36742\,
            I => \N__36731\
        );

    \I__7467\ : Odrv4
    port map (
            O => \N__36737\,
            I => n14742
        );

    \I__7466\ : Odrv4
    port map (
            O => \N__36734\,
            I => n14742
        );

    \I__7465\ : Odrv12
    port map (
            O => \N__36731\,
            I => n14742
        );

    \I__7464\ : CascadeMux
    port map (
            O => \N__36724\,
            I => \N__36721\
        );

    \I__7463\ : InMux
    port map (
            O => \N__36721\,
            I => \N__36718\
        );

    \I__7462\ : LocalMux
    port map (
            O => \N__36718\,
            I => \N__36714\
        );

    \I__7461\ : InMux
    port map (
            O => \N__36717\,
            I => \N__36710\
        );

    \I__7460\ : Span4Mux_v
    port map (
            O => \N__36714\,
            I => \N__36707\
        );

    \I__7459\ : InMux
    port map (
            O => \N__36713\,
            I => \N__36704\
        );

    \I__7458\ : LocalMux
    port map (
            O => \N__36710\,
            I => buf_dds0_3
        );

    \I__7457\ : Odrv4
    port map (
            O => \N__36707\,
            I => buf_dds0_3
        );

    \I__7456\ : LocalMux
    port map (
            O => \N__36704\,
            I => buf_dds0_3
        );

    \I__7455\ : InMux
    port map (
            O => \N__36697\,
            I => \N__36694\
        );

    \I__7454\ : LocalMux
    port map (
            O => \N__36694\,
            I => \SIG_DDS.tmp_buf_2\
        );

    \I__7453\ : CascadeMux
    port map (
            O => \N__36691\,
            I => \N__36688\
        );

    \I__7452\ : InMux
    port map (
            O => \N__36688\,
            I => \N__36685\
        );

    \I__7451\ : LocalMux
    port map (
            O => \N__36685\,
            I => \SIG_DDS.tmp_buf_3\
        );

    \I__7450\ : InMux
    port map (
            O => \N__36682\,
            I => \N__36679\
        );

    \I__7449\ : LocalMux
    port map (
            O => \N__36679\,
            I => \N__36675\
        );

    \I__7448\ : InMux
    port map (
            O => \N__36678\,
            I => \N__36672\
        );

    \I__7447\ : Span4Mux_v
    port map (
            O => \N__36675\,
            I => \N__36669\
        );

    \I__7446\ : LocalMux
    port map (
            O => \N__36672\,
            I => data_idxvec_7
        );

    \I__7445\ : Odrv4
    port map (
            O => \N__36669\,
            I => data_idxvec_7
        );

    \I__7444\ : InMux
    port map (
            O => \N__36664\,
            I => \N__36661\
        );

    \I__7443\ : LocalMux
    port map (
            O => \N__36661\,
            I => \N__36658\
        );

    \I__7442\ : Span4Mux_v
    port map (
            O => \N__36658\,
            I => \N__36654\
        );

    \I__7441\ : InMux
    port map (
            O => \N__36657\,
            I => \N__36650\
        );

    \I__7440\ : Span4Mux_h
    port map (
            O => \N__36654\,
            I => \N__36647\
        );

    \I__7439\ : InMux
    port map (
            O => \N__36653\,
            I => \N__36644\
        );

    \I__7438\ : LocalMux
    port map (
            O => \N__36650\,
            I => \acadc_skipCount_14\
        );

    \I__7437\ : Odrv4
    port map (
            O => \N__36647\,
            I => \acadc_skipCount_14\
        );

    \I__7436\ : LocalMux
    port map (
            O => \N__36644\,
            I => \acadc_skipCount_14\
        );

    \I__7435\ : InMux
    port map (
            O => \N__36637\,
            I => \N__36631\
        );

    \I__7434\ : InMux
    port map (
            O => \N__36636\,
            I => \N__36631\
        );

    \I__7433\ : LocalMux
    port map (
            O => \N__36631\,
            I => n8_adj_1545
        );

    \I__7432\ : InMux
    port map (
            O => \N__36628\,
            I => \N__36624\
        );

    \I__7431\ : InMux
    port map (
            O => \N__36627\,
            I => \N__36621\
        );

    \I__7430\ : LocalMux
    port map (
            O => \N__36624\,
            I => \N__36618\
        );

    \I__7429\ : LocalMux
    port map (
            O => \N__36621\,
            I => acadc_skipcnt_9
        );

    \I__7428\ : Odrv4
    port map (
            O => \N__36618\,
            I => acadc_skipcnt_9
        );

    \I__7427\ : InMux
    port map (
            O => \N__36613\,
            I => \N__36609\
        );

    \I__7426\ : InMux
    port map (
            O => \N__36612\,
            I => \N__36606\
        );

    \I__7425\ : LocalMux
    port map (
            O => \N__36609\,
            I => \N__36603\
        );

    \I__7424\ : LocalMux
    port map (
            O => \N__36606\,
            I => acadc_skipcnt_15
        );

    \I__7423\ : Odrv4
    port map (
            O => \N__36603\,
            I => acadc_skipcnt_15
        );

    \I__7422\ : InMux
    port map (
            O => \N__36598\,
            I => \N__36595\
        );

    \I__7421\ : LocalMux
    port map (
            O => \N__36595\,
            I => \N__36592\
        );

    \I__7420\ : Span4Mux_h
    port map (
            O => \N__36592\,
            I => \N__36589\
        );

    \I__7419\ : Span4Mux_v
    port map (
            O => \N__36589\,
            I => \N__36584\
        );

    \I__7418\ : InMux
    port map (
            O => \N__36588\,
            I => \N__36579\
        );

    \I__7417\ : InMux
    port map (
            O => \N__36587\,
            I => \N__36579\
        );

    \I__7416\ : Odrv4
    port map (
            O => \N__36584\,
            I => \acadc_skipCount_15\
        );

    \I__7415\ : LocalMux
    port map (
            O => \N__36579\,
            I => \acadc_skipCount_15\
        );

    \I__7414\ : InMux
    port map (
            O => \N__36574\,
            I => \N__36571\
        );

    \I__7413\ : LocalMux
    port map (
            O => \N__36571\,
            I => n24
        );

    \I__7412\ : CascadeMux
    port map (
            O => \N__36568\,
            I => \N__36565\
        );

    \I__7411\ : InMux
    port map (
            O => \N__36565\,
            I => \N__36560\
        );

    \I__7410\ : InMux
    port map (
            O => \N__36564\,
            I => \N__36557\
        );

    \I__7409\ : InMux
    port map (
            O => \N__36563\,
            I => \N__36554\
        );

    \I__7408\ : LocalMux
    port map (
            O => \N__36560\,
            I => \N__36551\
        );

    \I__7407\ : LocalMux
    port map (
            O => \N__36557\,
            I => \N__36548\
        );

    \I__7406\ : LocalMux
    port map (
            O => \N__36554\,
            I => \N__36545\
        );

    \I__7405\ : Odrv4
    port map (
            O => \N__36551\,
            I => \acadc_skipCount_1\
        );

    \I__7404\ : Odrv4
    port map (
            O => \N__36548\,
            I => \acadc_skipCount_1\
        );

    \I__7403\ : Odrv12
    port map (
            O => \N__36545\,
            I => \acadc_skipCount_1\
        );

    \I__7402\ : InMux
    port map (
            O => \N__36538\,
            I => \N__36535\
        );

    \I__7401\ : LocalMux
    port map (
            O => \N__36535\,
            I => \N__36532\
        );

    \I__7400\ : Span4Mux_h
    port map (
            O => \N__36532\,
            I => \N__36529\
        );

    \I__7399\ : Odrv4
    port map (
            O => \N__36529\,
            I => n9_adj_1407
        );

    \I__7398\ : CascadeMux
    port map (
            O => \N__36526\,
            I => \N__36523\
        );

    \I__7397\ : CascadeBuf
    port map (
            O => \N__36523\,
            I => \N__36520\
        );

    \I__7396\ : CascadeMux
    port map (
            O => \N__36520\,
            I => \N__36517\
        );

    \I__7395\ : CascadeBuf
    port map (
            O => \N__36517\,
            I => \N__36514\
        );

    \I__7394\ : CascadeMux
    port map (
            O => \N__36514\,
            I => \N__36511\
        );

    \I__7393\ : CascadeBuf
    port map (
            O => \N__36511\,
            I => \N__36508\
        );

    \I__7392\ : CascadeMux
    port map (
            O => \N__36508\,
            I => \N__36505\
        );

    \I__7391\ : CascadeBuf
    port map (
            O => \N__36505\,
            I => \N__36502\
        );

    \I__7390\ : CascadeMux
    port map (
            O => \N__36502\,
            I => \N__36499\
        );

    \I__7389\ : CascadeBuf
    port map (
            O => \N__36499\,
            I => \N__36496\
        );

    \I__7388\ : CascadeMux
    port map (
            O => \N__36496\,
            I => \N__36493\
        );

    \I__7387\ : CascadeBuf
    port map (
            O => \N__36493\,
            I => \N__36490\
        );

    \I__7386\ : CascadeMux
    port map (
            O => \N__36490\,
            I => \N__36487\
        );

    \I__7385\ : CascadeBuf
    port map (
            O => \N__36487\,
            I => \N__36484\
        );

    \I__7384\ : CascadeMux
    port map (
            O => \N__36484\,
            I => \N__36481\
        );

    \I__7383\ : CascadeBuf
    port map (
            O => \N__36481\,
            I => \N__36478\
        );

    \I__7382\ : CascadeMux
    port map (
            O => \N__36478\,
            I => \N__36474\
        );

    \I__7381\ : CascadeMux
    port map (
            O => \N__36477\,
            I => \N__36471\
        );

    \I__7380\ : CascadeBuf
    port map (
            O => \N__36474\,
            I => \N__36468\
        );

    \I__7379\ : CascadeBuf
    port map (
            O => \N__36471\,
            I => \N__36465\
        );

    \I__7378\ : CascadeMux
    port map (
            O => \N__36468\,
            I => \N__36462\
        );

    \I__7377\ : CascadeMux
    port map (
            O => \N__36465\,
            I => \N__36459\
        );

    \I__7376\ : InMux
    port map (
            O => \N__36462\,
            I => \N__36456\
        );

    \I__7375\ : InMux
    port map (
            O => \N__36459\,
            I => \N__36453\
        );

    \I__7374\ : LocalMux
    port map (
            O => \N__36456\,
            I => \N__36450\
        );

    \I__7373\ : LocalMux
    port map (
            O => \N__36453\,
            I => \N__36447\
        );

    \I__7372\ : Span4Mux_v
    port map (
            O => \N__36450\,
            I => \N__36444\
        );

    \I__7371\ : Span4Mux_v
    port map (
            O => \N__36447\,
            I => \N__36441\
        );

    \I__7370\ : Span4Mux_h
    port map (
            O => \N__36444\,
            I => \N__36438\
        );

    \I__7369\ : Span4Mux_h
    port map (
            O => \N__36441\,
            I => \N__36433\
        );

    \I__7368\ : Span4Mux_h
    port map (
            O => \N__36438\,
            I => \N__36433\
        );

    \I__7367\ : Odrv4
    port map (
            O => \N__36433\,
            I => \data_index_9_N_212_2\
        );

    \I__7366\ : InMux
    port map (
            O => \N__36430\,
            I => \N__36427\
        );

    \I__7365\ : LocalMux
    port map (
            O => \N__36427\,
            I => \N__36423\
        );

    \I__7364\ : InMux
    port map (
            O => \N__36426\,
            I => \N__36420\
        );

    \I__7363\ : Span4Mux_v
    port map (
            O => \N__36423\,
            I => \N__36417\
        );

    \I__7362\ : LocalMux
    port map (
            O => \N__36420\,
            I => acadc_skipcnt_14
        );

    \I__7361\ : Odrv4
    port map (
            O => \N__36417\,
            I => acadc_skipcnt_14
        );

    \I__7360\ : InMux
    port map (
            O => \N__36412\,
            I => \N__36408\
        );

    \I__7359\ : InMux
    port map (
            O => \N__36411\,
            I => \N__36405\
        );

    \I__7358\ : LocalMux
    port map (
            O => \N__36408\,
            I => \N__36402\
        );

    \I__7357\ : LocalMux
    port map (
            O => \N__36405\,
            I => acadc_skipcnt_11
        );

    \I__7356\ : Odrv4
    port map (
            O => \N__36402\,
            I => acadc_skipcnt_11
        );

    \I__7355\ : InMux
    port map (
            O => \N__36397\,
            I => \N__36391\
        );

    \I__7354\ : CascadeMux
    port map (
            O => \N__36396\,
            I => \N__36388\
        );

    \I__7353\ : InMux
    port map (
            O => \N__36395\,
            I => \N__36385\
        );

    \I__7352\ : InMux
    port map (
            O => \N__36394\,
            I => \N__36382\
        );

    \I__7351\ : LocalMux
    port map (
            O => \N__36391\,
            I => \N__36379\
        );

    \I__7350\ : InMux
    port map (
            O => \N__36388\,
            I => \N__36375\
        );

    \I__7349\ : LocalMux
    port map (
            O => \N__36385\,
            I => \N__36370\
        );

    \I__7348\ : LocalMux
    port map (
            O => \N__36382\,
            I => \N__36370\
        );

    \I__7347\ : Span4Mux_v
    port map (
            O => \N__36379\,
            I => \N__36367\
        );

    \I__7346\ : InMux
    port map (
            O => \N__36378\,
            I => \N__36364\
        );

    \I__7345\ : LocalMux
    port map (
            O => \N__36375\,
            I => \N__36361\
        );

    \I__7344\ : Span12Mux_v
    port map (
            O => \N__36370\,
            I => \N__36358\
        );

    \I__7343\ : Span4Mux_h
    port map (
            O => \N__36367\,
            I => \N__36353\
        );

    \I__7342\ : LocalMux
    port map (
            O => \N__36364\,
            I => \N__36353\
        );

    \I__7341\ : Odrv12
    port map (
            O => \N__36361\,
            I => comm_buf_1_3
        );

    \I__7340\ : Odrv12
    port map (
            O => \N__36358\,
            I => comm_buf_1_3
        );

    \I__7339\ : Odrv4
    port map (
            O => \N__36353\,
            I => comm_buf_1_3
        );

    \I__7338\ : InMux
    port map (
            O => \N__36346\,
            I => \N__36340\
        );

    \I__7337\ : InMux
    port map (
            O => \N__36345\,
            I => \N__36340\
        );

    \I__7336\ : LocalMux
    port map (
            O => \N__36340\,
            I => \N__36337\
        );

    \I__7335\ : Odrv12
    port map (
            O => \N__36337\,
            I => n8_adj_1543
        );

    \I__7334\ : InMux
    port map (
            O => \N__36334\,
            I => \N__36330\
        );

    \I__7333\ : InMux
    port map (
            O => \N__36333\,
            I => \N__36327\
        );

    \I__7332\ : LocalMux
    port map (
            O => \N__36330\,
            I => \N__36324\
        );

    \I__7331\ : LocalMux
    port map (
            O => \N__36327\,
            I => acadc_skipcnt_2
        );

    \I__7330\ : Odrv4
    port map (
            O => \N__36324\,
            I => acadc_skipcnt_2
        );

    \I__7329\ : InMux
    port map (
            O => \N__36319\,
            I => \N__36315\
        );

    \I__7328\ : InMux
    port map (
            O => \N__36318\,
            I => \N__36312\
        );

    \I__7327\ : LocalMux
    port map (
            O => \N__36315\,
            I => \N__36309\
        );

    \I__7326\ : LocalMux
    port map (
            O => \N__36312\,
            I => acadc_skipcnt_7
        );

    \I__7325\ : Odrv4
    port map (
            O => \N__36309\,
            I => acadc_skipcnt_7
        );

    \I__7324\ : InMux
    port map (
            O => \N__36304\,
            I => \N__36299\
        );

    \I__7323\ : CascadeMux
    port map (
            O => \N__36303\,
            I => \N__36296\
        );

    \I__7322\ : InMux
    port map (
            O => \N__36302\,
            I => \N__36293\
        );

    \I__7321\ : LocalMux
    port map (
            O => \N__36299\,
            I => \N__36290\
        );

    \I__7320\ : InMux
    port map (
            O => \N__36296\,
            I => \N__36287\
        );

    \I__7319\ : LocalMux
    port map (
            O => \N__36293\,
            I => \acadc_skipCount_2\
        );

    \I__7318\ : Odrv4
    port map (
            O => \N__36290\,
            I => \acadc_skipCount_2\
        );

    \I__7317\ : LocalMux
    port map (
            O => \N__36287\,
            I => \acadc_skipCount_2\
        );

    \I__7316\ : InMux
    port map (
            O => \N__36280\,
            I => \N__36277\
        );

    \I__7315\ : LocalMux
    port map (
            O => \N__36277\,
            I => n23_adj_1586
        );

    \I__7314\ : CascadeMux
    port map (
            O => \N__36274\,
            I => \n22_cascade_\
        );

    \I__7313\ : InMux
    port map (
            O => \N__36271\,
            I => \N__36268\
        );

    \I__7312\ : LocalMux
    port map (
            O => \N__36268\,
            I => \N__36265\
        );

    \I__7311\ : Odrv4
    port map (
            O => \N__36265\,
            I => n30_adj_1571
        );

    \I__7310\ : CascadeMux
    port map (
            O => \N__36262\,
            I => \n30_adj_1478_cascade_\
        );

    \I__7309\ : InMux
    port map (
            O => \N__36259\,
            I => \N__36256\
        );

    \I__7308\ : LocalMux
    port map (
            O => \N__36256\,
            I => \N__36249\
        );

    \I__7307\ : InMux
    port map (
            O => \N__36255\,
            I => \N__36246\
        );

    \I__7306\ : InMux
    port map (
            O => \N__36254\,
            I => \N__36243\
        );

    \I__7305\ : InMux
    port map (
            O => \N__36253\,
            I => \N__36238\
        );

    \I__7304\ : InMux
    port map (
            O => \N__36252\,
            I => \N__36234\
        );

    \I__7303\ : Span4Mux_v
    port map (
            O => \N__36249\,
            I => \N__36228\
        );

    \I__7302\ : LocalMux
    port map (
            O => \N__36246\,
            I => \N__36228\
        );

    \I__7301\ : LocalMux
    port map (
            O => \N__36243\,
            I => \N__36225\
        );

    \I__7300\ : InMux
    port map (
            O => \N__36242\,
            I => \N__36222\
        );

    \I__7299\ : InMux
    port map (
            O => \N__36241\,
            I => \N__36219\
        );

    \I__7298\ : LocalMux
    port map (
            O => \N__36238\,
            I => \N__36216\
        );

    \I__7297\ : InMux
    port map (
            O => \N__36237\,
            I => \N__36213\
        );

    \I__7296\ : LocalMux
    port map (
            O => \N__36234\,
            I => \N__36210\
        );

    \I__7295\ : InMux
    port map (
            O => \N__36233\,
            I => \N__36207\
        );

    \I__7294\ : Span4Mux_v
    port map (
            O => \N__36228\,
            I => \N__36204\
        );

    \I__7293\ : Span4Mux_v
    port map (
            O => \N__36225\,
            I => \N__36199\
        );

    \I__7292\ : LocalMux
    port map (
            O => \N__36222\,
            I => \N__36199\
        );

    \I__7291\ : LocalMux
    port map (
            O => \N__36219\,
            I => \N__36188\
        );

    \I__7290\ : Span4Mux_v
    port map (
            O => \N__36216\,
            I => \N__36188\
        );

    \I__7289\ : LocalMux
    port map (
            O => \N__36213\,
            I => \N__36188\
        );

    \I__7288\ : Span4Mux_h
    port map (
            O => \N__36210\,
            I => \N__36188\
        );

    \I__7287\ : LocalMux
    port map (
            O => \N__36207\,
            I => \N__36188\
        );

    \I__7286\ : Span4Mux_h
    port map (
            O => \N__36204\,
            I => \N__36185\
        );

    \I__7285\ : Span4Mux_v
    port map (
            O => \N__36199\,
            I => \N__36182\
        );

    \I__7284\ : Span4Mux_v
    port map (
            O => \N__36188\,
            I => \N__36179\
        );

    \I__7283\ : Span4Mux_v
    port map (
            O => \N__36185\,
            I => \N__36176\
        );

    \I__7282\ : Span4Mux_v
    port map (
            O => \N__36182\,
            I => \N__36171\
        );

    \I__7281\ : Span4Mux_v
    port map (
            O => \N__36179\,
            I => \N__36171\
        );

    \I__7280\ : Odrv4
    port map (
            O => \N__36176\,
            I => comm_rx_buf_0
        );

    \I__7279\ : Odrv4
    port map (
            O => \N__36171\,
            I => comm_rx_buf_0
        );

    \I__7278\ : CascadeMux
    port map (
            O => \N__36166\,
            I => \N__36161\
        );

    \I__7277\ : InMux
    port map (
            O => \N__36165\,
            I => \N__36154\
        );

    \I__7276\ : InMux
    port map (
            O => \N__36164\,
            I => \N__36154\
        );

    \I__7275\ : InMux
    port map (
            O => \N__36161\,
            I => \N__36154\
        );

    \I__7274\ : LocalMux
    port map (
            O => \N__36154\,
            I => cmd_rdadctmp_13_adj_1430
        );

    \I__7273\ : InMux
    port map (
            O => \N__36151\,
            I => \N__36148\
        );

    \I__7272\ : LocalMux
    port map (
            O => \N__36148\,
            I => \N__36145\
        );

    \I__7271\ : Span4Mux_v
    port map (
            O => \N__36145\,
            I => \N__36140\
        );

    \I__7270\ : InMux
    port map (
            O => \N__36144\,
            I => \N__36137\
        );

    \I__7269\ : InMux
    port map (
            O => \N__36143\,
            I => \N__36134\
        );

    \I__7268\ : Span4Mux_h
    port map (
            O => \N__36140\,
            I => \N__36131\
        );

    \I__7267\ : LocalMux
    port map (
            O => \N__36137\,
            I => buf_dds1_4
        );

    \I__7266\ : LocalMux
    port map (
            O => \N__36134\,
            I => buf_dds1_4
        );

    \I__7265\ : Odrv4
    port map (
            O => \N__36131\,
            I => buf_dds1_4
        );

    \I__7264\ : InMux
    port map (
            O => \N__36124\,
            I => \N__36121\
        );

    \I__7263\ : LocalMux
    port map (
            O => \N__36121\,
            I => \N__36118\
        );

    \I__7262\ : Odrv4
    port map (
            O => \N__36118\,
            I => n16
        );

    \I__7261\ : InMux
    port map (
            O => \N__36115\,
            I => \N__36112\
        );

    \I__7260\ : LocalMux
    port map (
            O => \N__36112\,
            I => \N__36109\
        );

    \I__7259\ : Span4Mux_v
    port map (
            O => \N__36109\,
            I => \N__36105\
        );

    \I__7258\ : InMux
    port map (
            O => \N__36108\,
            I => \N__36101\
        );

    \I__7257\ : Span4Mux_h
    port map (
            O => \N__36105\,
            I => \N__36098\
        );

    \I__7256\ : InMux
    port map (
            O => \N__36104\,
            I => \N__36095\
        );

    \I__7255\ : LocalMux
    port map (
            O => \N__36101\,
            I => buf_dds1_6
        );

    \I__7254\ : Odrv4
    port map (
            O => \N__36098\,
            I => buf_dds1_6
        );

    \I__7253\ : LocalMux
    port map (
            O => \N__36095\,
            I => buf_dds1_6
        );

    \I__7252\ : InMux
    port map (
            O => \N__36088\,
            I => \N__36085\
        );

    \I__7251\ : LocalMux
    port map (
            O => \N__36085\,
            I => \N__36082\
        );

    \I__7250\ : Odrv4
    port map (
            O => \N__36082\,
            I => n16_adj_1488
        );

    \I__7249\ : CascadeMux
    port map (
            O => \N__36079\,
            I => \N__36076\
        );

    \I__7248\ : InMux
    port map (
            O => \N__36076\,
            I => \N__36073\
        );

    \I__7247\ : LocalMux
    port map (
            O => \N__36073\,
            I => \N__36070\
        );

    \I__7246\ : Odrv4
    port map (
            O => \N__36070\,
            I => n20824
        );

    \I__7245\ : InMux
    port map (
            O => \N__36067\,
            I => \N__36064\
        );

    \I__7244\ : LocalMux
    port map (
            O => \N__36064\,
            I => \N__36061\
        );

    \I__7243\ : Span4Mux_v
    port map (
            O => \N__36061\,
            I => \N__36058\
        );

    \I__7242\ : Span4Mux_h
    port map (
            O => \N__36058\,
            I => \N__36055\
        );

    \I__7241\ : Span4Mux_h
    port map (
            O => \N__36055\,
            I => \N__36052\
        );

    \I__7240\ : Odrv4
    port map (
            O => \N__36052\,
            I => n20836
        );

    \I__7239\ : CascadeMux
    port map (
            O => \N__36049\,
            I => \n22069_cascade_\
        );

    \I__7238\ : InMux
    port map (
            O => \N__36046\,
            I => \N__36043\
        );

    \I__7237\ : LocalMux
    port map (
            O => \N__36043\,
            I => n20837
        );

    \I__7236\ : InMux
    port map (
            O => \N__36040\,
            I => \N__36036\
        );

    \I__7235\ : InMux
    port map (
            O => \N__36039\,
            I => \N__36033\
        );

    \I__7234\ : LocalMux
    port map (
            O => \N__36036\,
            I => \N__36030\
        );

    \I__7233\ : LocalMux
    port map (
            O => \N__36033\,
            I => data_idxvec_1
        );

    \I__7232\ : Odrv4
    port map (
            O => \N__36030\,
            I => data_idxvec_1
        );

    \I__7231\ : CascadeMux
    port map (
            O => \N__36025\,
            I => \n26_adj_1509_cascade_\
        );

    \I__7230\ : InMux
    port map (
            O => \N__36022\,
            I => \N__36019\
        );

    \I__7229\ : LocalMux
    port map (
            O => \N__36019\,
            I => \N__36016\
        );

    \I__7228\ : Span4Mux_h
    port map (
            O => \N__36016\,
            I => \N__36013\
        );

    \I__7227\ : Span4Mux_v
    port map (
            O => \N__36013\,
            I => \N__36010\
        );

    \I__7226\ : Span4Mux_h
    port map (
            O => \N__36010\,
            I => \N__36007\
        );

    \I__7225\ : Span4Mux_h
    port map (
            O => \N__36007\,
            I => \N__36004\
        );

    \I__7224\ : Odrv4
    port map (
            O => \N__36004\,
            I => buf_data_iac_9
        );

    \I__7223\ : InMux
    port map (
            O => \N__36001\,
            I => \N__35998\
        );

    \I__7222\ : LocalMux
    port map (
            O => \N__35998\,
            I => n20825
        );

    \I__7221\ : InMux
    port map (
            O => \N__35995\,
            I => \N__35992\
        );

    \I__7220\ : LocalMux
    port map (
            O => \N__35992\,
            I => \N__35988\
        );

    \I__7219\ : InMux
    port map (
            O => \N__35991\,
            I => \N__35985\
        );

    \I__7218\ : Span4Mux_v
    port map (
            O => \N__35988\,
            I => \N__35982\
        );

    \I__7217\ : LocalMux
    port map (
            O => \N__35985\,
            I => \N__35979\
        );

    \I__7216\ : Span4Mux_h
    port map (
            O => \N__35982\,
            I => \N__35972\
        );

    \I__7215\ : Span4Mux_h
    port map (
            O => \N__35979\,
            I => \N__35972\
        );

    \I__7214\ : CascadeMux
    port map (
            O => \N__35978\,
            I => \N__35968\
        );

    \I__7213\ : InMux
    port map (
            O => \N__35977\,
            I => \N__35964\
        );

    \I__7212\ : Span4Mux_h
    port map (
            O => \N__35972\,
            I => \N__35961\
        );

    \I__7211\ : InMux
    port map (
            O => \N__35971\,
            I => \N__35958\
        );

    \I__7210\ : InMux
    port map (
            O => \N__35968\,
            I => \N__35955\
        );

    \I__7209\ : InMux
    port map (
            O => \N__35967\,
            I => \N__35952\
        );

    \I__7208\ : LocalMux
    port map (
            O => \N__35964\,
            I => \N__35948\
        );

    \I__7207\ : Span4Mux_h
    port map (
            O => \N__35961\,
            I => \N__35943\
        );

    \I__7206\ : LocalMux
    port map (
            O => \N__35958\,
            I => \N__35943\
        );

    \I__7205\ : LocalMux
    port map (
            O => \N__35955\,
            I => \N__35938\
        );

    \I__7204\ : LocalMux
    port map (
            O => \N__35952\,
            I => \N__35938\
        );

    \I__7203\ : InMux
    port map (
            O => \N__35951\,
            I => \N__35935\
        );

    \I__7202\ : Span4Mux_h
    port map (
            O => \N__35948\,
            I => \N__35930\
        );

    \I__7201\ : Span4Mux_v
    port map (
            O => \N__35943\,
            I => \N__35927\
        );

    \I__7200\ : Span4Mux_h
    port map (
            O => \N__35938\,
            I => \N__35922\
        );

    \I__7199\ : LocalMux
    port map (
            O => \N__35935\,
            I => \N__35922\
        );

    \I__7198\ : InMux
    port map (
            O => \N__35934\,
            I => \N__35919\
        );

    \I__7197\ : InMux
    port map (
            O => \N__35933\,
            I => \N__35916\
        );

    \I__7196\ : Odrv4
    port map (
            O => \N__35930\,
            I => comm_rx_buf_1
        );

    \I__7195\ : Odrv4
    port map (
            O => \N__35927\,
            I => comm_rx_buf_1
        );

    \I__7194\ : Odrv4
    port map (
            O => \N__35922\,
            I => comm_rx_buf_1
        );

    \I__7193\ : LocalMux
    port map (
            O => \N__35919\,
            I => comm_rx_buf_1
        );

    \I__7192\ : LocalMux
    port map (
            O => \N__35916\,
            I => comm_rx_buf_1
        );

    \I__7191\ : InMux
    port map (
            O => \N__35905\,
            I => \N__35902\
        );

    \I__7190\ : LocalMux
    port map (
            O => \N__35902\,
            I => n22072
        );

    \I__7189\ : InMux
    port map (
            O => \N__35899\,
            I => \N__35896\
        );

    \I__7188\ : LocalMux
    port map (
            O => \N__35896\,
            I => \N__35892\
        );

    \I__7187\ : InMux
    port map (
            O => \N__35895\,
            I => \N__35889\
        );

    \I__7186\ : Span4Mux_h
    port map (
            O => \N__35892\,
            I => \N__35886\
        );

    \I__7185\ : LocalMux
    port map (
            O => \N__35889\,
            I => data_idxvec_0
        );

    \I__7184\ : Odrv4
    port map (
            O => \N__35886\,
            I => data_idxvec_0
        );

    \I__7183\ : InMux
    port map (
            O => \N__35881\,
            I => \N__35878\
        );

    \I__7182\ : LocalMux
    port map (
            O => \N__35878\,
            I => \N__35875\
        );

    \I__7181\ : Span4Mux_h
    port map (
            O => \N__35875\,
            I => \N__35872\
        );

    \I__7180\ : Span4Mux_h
    port map (
            O => \N__35872\,
            I => \N__35869\
        );

    \I__7179\ : Span4Mux_h
    port map (
            O => \N__35869\,
            I => \N__35866\
        );

    \I__7178\ : Odrv4
    port map (
            O => \N__35866\,
            I => n21001
        );

    \I__7177\ : CascadeMux
    port map (
            O => \N__35863\,
            I => \n26_cascade_\
        );

    \I__7176\ : InMux
    port map (
            O => \N__35860\,
            I => \N__35857\
        );

    \I__7175\ : LocalMux
    port map (
            O => \N__35857\,
            I => \N__35852\
        );

    \I__7174\ : InMux
    port map (
            O => \N__35856\,
            I => \N__35849\
        );

    \I__7173\ : InMux
    port map (
            O => \N__35855\,
            I => \N__35846\
        );

    \I__7172\ : Span4Mux_v
    port map (
            O => \N__35852\,
            I => \N__35843\
        );

    \I__7171\ : LocalMux
    port map (
            O => \N__35849\,
            I => \N__35838\
        );

    \I__7170\ : LocalMux
    port map (
            O => \N__35846\,
            I => \N__35838\
        );

    \I__7169\ : Odrv4
    port map (
            O => \N__35843\,
            I => \acadc_skipCount_0\
        );

    \I__7168\ : Odrv4
    port map (
            O => \N__35838\,
            I => \acadc_skipCount_0\
        );

    \I__7167\ : CascadeMux
    port map (
            O => \N__35833\,
            I => \n22021_cascade_\
        );

    \I__7166\ : InMux
    port map (
            O => \N__35830\,
            I => \N__35827\
        );

    \I__7165\ : LocalMux
    port map (
            O => \N__35827\,
            I => n22024
        );

    \I__7164\ : InMux
    port map (
            O => \N__35824\,
            I => \N__35821\
        );

    \I__7163\ : LocalMux
    port map (
            O => \N__35821\,
            I => \N__35818\
        );

    \I__7162\ : Span12Mux_v
    port map (
            O => \N__35818\,
            I => \N__35815\
        );

    \I__7161\ : Odrv12
    port map (
            O => \N__35815\,
            I => n21976
        );

    \I__7160\ : InMux
    port map (
            O => \N__35812\,
            I => \N__35807\
        );

    \I__7159\ : CascadeMux
    port map (
            O => \N__35811\,
            I => \N__35803\
        );

    \I__7158\ : InMux
    port map (
            O => \N__35810\,
            I => \N__35799\
        );

    \I__7157\ : LocalMux
    port map (
            O => \N__35807\,
            I => \N__35795\
        );

    \I__7156\ : InMux
    port map (
            O => \N__35806\,
            I => \N__35792\
        );

    \I__7155\ : InMux
    port map (
            O => \N__35803\,
            I => \N__35789\
        );

    \I__7154\ : InMux
    port map (
            O => \N__35802\,
            I => \N__35786\
        );

    \I__7153\ : LocalMux
    port map (
            O => \N__35799\,
            I => \N__35783\
        );

    \I__7152\ : InMux
    port map (
            O => \N__35798\,
            I => \N__35780\
        );

    \I__7151\ : Span4Mux_h
    port map (
            O => \N__35795\,
            I => \N__35776\
        );

    \I__7150\ : LocalMux
    port map (
            O => \N__35792\,
            I => \N__35773\
        );

    \I__7149\ : LocalMux
    port map (
            O => \N__35789\,
            I => \N__35770\
        );

    \I__7148\ : LocalMux
    port map (
            O => \N__35786\,
            I => \N__35767\
        );

    \I__7147\ : Span4Mux_v
    port map (
            O => \N__35783\,
            I => \N__35762\
        );

    \I__7146\ : LocalMux
    port map (
            O => \N__35780\,
            I => \N__35762\
        );

    \I__7145\ : InMux
    port map (
            O => \N__35779\,
            I => \N__35759\
        );

    \I__7144\ : Span4Mux_v
    port map (
            O => \N__35776\,
            I => \N__35754\
        );

    \I__7143\ : Span4Mux_v
    port map (
            O => \N__35773\,
            I => \N__35751\
        );

    \I__7142\ : Span4Mux_h
    port map (
            O => \N__35770\,
            I => \N__35748\
        );

    \I__7141\ : Span4Mux_h
    port map (
            O => \N__35767\,
            I => \N__35745\
        );

    \I__7140\ : Span4Mux_h
    port map (
            O => \N__35762\,
            I => \N__35742\
        );

    \I__7139\ : LocalMux
    port map (
            O => \N__35759\,
            I => \N__35739\
        );

    \I__7138\ : InMux
    port map (
            O => \N__35758\,
            I => \N__35736\
        );

    \I__7137\ : InMux
    port map (
            O => \N__35757\,
            I => \N__35733\
        );

    \I__7136\ : Odrv4
    port map (
            O => \N__35754\,
            I => comm_rx_buf_6
        );

    \I__7135\ : Odrv4
    port map (
            O => \N__35751\,
            I => comm_rx_buf_6
        );

    \I__7134\ : Odrv4
    port map (
            O => \N__35748\,
            I => comm_rx_buf_6
        );

    \I__7133\ : Odrv4
    port map (
            O => \N__35745\,
            I => comm_rx_buf_6
        );

    \I__7132\ : Odrv4
    port map (
            O => \N__35742\,
            I => comm_rx_buf_6
        );

    \I__7131\ : Odrv12
    port map (
            O => \N__35739\,
            I => comm_rx_buf_6
        );

    \I__7130\ : LocalMux
    port map (
            O => \N__35736\,
            I => comm_rx_buf_6
        );

    \I__7129\ : LocalMux
    port map (
            O => \N__35733\,
            I => comm_rx_buf_6
        );

    \I__7128\ : InMux
    port map (
            O => \N__35716\,
            I => \N__35713\
        );

    \I__7127\ : LocalMux
    port map (
            O => \N__35713\,
            I => \N__35710\
        );

    \I__7126\ : Span4Mux_h
    port map (
            O => \N__35710\,
            I => \N__35707\
        );

    \I__7125\ : Span4Mux_h
    port map (
            O => \N__35707\,
            I => \N__35704\
        );

    \I__7124\ : Odrv4
    port map (
            O => \N__35704\,
            I => buf_data_vac_6
        );

    \I__7123\ : InMux
    port map (
            O => \N__35701\,
            I => \N__35698\
        );

    \I__7122\ : LocalMux
    port map (
            O => \N__35698\,
            I => \N__35695\
        );

    \I__7121\ : Span4Mux_v
    port map (
            O => \N__35695\,
            I => \N__35692\
        );

    \I__7120\ : Odrv4
    port map (
            O => \N__35692\,
            I => comm_buf_5_6
        );

    \I__7119\ : InMux
    port map (
            O => \N__35689\,
            I => \N__35686\
        );

    \I__7118\ : LocalMux
    port map (
            O => \N__35686\,
            I => \N__35683\
        );

    \I__7117\ : Span4Mux_h
    port map (
            O => \N__35683\,
            I => \N__35680\
        );

    \I__7116\ : Span4Mux_h
    port map (
            O => \N__35680\,
            I => \N__35677\
        );

    \I__7115\ : Odrv4
    port map (
            O => \N__35677\,
            I => buf_data_vac_5
        );

    \I__7114\ : InMux
    port map (
            O => \N__35674\,
            I => \N__35671\
        );

    \I__7113\ : LocalMux
    port map (
            O => \N__35671\,
            I => comm_buf_5_5
        );

    \I__7112\ : InMux
    port map (
            O => \N__35668\,
            I => \N__35665\
        );

    \I__7111\ : LocalMux
    port map (
            O => \N__35665\,
            I => \N__35658\
        );

    \I__7110\ : InMux
    port map (
            O => \N__35664\,
            I => \N__35655\
        );

    \I__7109\ : CascadeMux
    port map (
            O => \N__35663\,
            I => \N__35652\
        );

    \I__7108\ : InMux
    port map (
            O => \N__35662\,
            I => \N__35649\
        );

    \I__7107\ : InMux
    port map (
            O => \N__35661\,
            I => \N__35646\
        );

    \I__7106\ : Span4Mux_h
    port map (
            O => \N__35658\,
            I => \N__35641\
        );

    \I__7105\ : LocalMux
    port map (
            O => \N__35655\,
            I => \N__35641\
        );

    \I__7104\ : InMux
    port map (
            O => \N__35652\,
            I => \N__35637\
        );

    \I__7103\ : LocalMux
    port map (
            O => \N__35649\,
            I => \N__35633\
        );

    \I__7102\ : LocalMux
    port map (
            O => \N__35646\,
            I => \N__35628\
        );

    \I__7101\ : Span4Mux_h
    port map (
            O => \N__35641\,
            I => \N__35628\
        );

    \I__7100\ : InMux
    port map (
            O => \N__35640\,
            I => \N__35625\
        );

    \I__7099\ : LocalMux
    port map (
            O => \N__35637\,
            I => \N__35622\
        );

    \I__7098\ : InMux
    port map (
            O => \N__35636\,
            I => \N__35619\
        );

    \I__7097\ : Span4Mux_h
    port map (
            O => \N__35633\,
            I => \N__35614\
        );

    \I__7096\ : Sp12to4
    port map (
            O => \N__35628\,
            I => \N__35611\
        );

    \I__7095\ : LocalMux
    port map (
            O => \N__35625\,
            I => \N__35608\
        );

    \I__7094\ : Span4Mux_h
    port map (
            O => \N__35622\,
            I => \N__35603\
        );

    \I__7093\ : LocalMux
    port map (
            O => \N__35619\,
            I => \N__35603\
        );

    \I__7092\ : InMux
    port map (
            O => \N__35618\,
            I => \N__35600\
        );

    \I__7091\ : InMux
    port map (
            O => \N__35617\,
            I => \N__35597\
        );

    \I__7090\ : Odrv4
    port map (
            O => \N__35614\,
            I => comm_rx_buf_4
        );

    \I__7089\ : Odrv12
    port map (
            O => \N__35611\,
            I => comm_rx_buf_4
        );

    \I__7088\ : Odrv12
    port map (
            O => \N__35608\,
            I => comm_rx_buf_4
        );

    \I__7087\ : Odrv4
    port map (
            O => \N__35603\,
            I => comm_rx_buf_4
        );

    \I__7086\ : LocalMux
    port map (
            O => \N__35600\,
            I => comm_rx_buf_4
        );

    \I__7085\ : LocalMux
    port map (
            O => \N__35597\,
            I => comm_rx_buf_4
        );

    \I__7084\ : InMux
    port map (
            O => \N__35584\,
            I => \N__35581\
        );

    \I__7083\ : LocalMux
    port map (
            O => \N__35581\,
            I => \N__35578\
        );

    \I__7082\ : Span4Mux_h
    port map (
            O => \N__35578\,
            I => \N__35575\
        );

    \I__7081\ : Span4Mux_h
    port map (
            O => \N__35575\,
            I => \N__35572\
        );

    \I__7080\ : Odrv4
    port map (
            O => \N__35572\,
            I => buf_data_vac_4
        );

    \I__7079\ : InMux
    port map (
            O => \N__35569\,
            I => \N__35564\
        );

    \I__7078\ : CascadeMux
    port map (
            O => \N__35568\,
            I => \N__35560\
        );

    \I__7077\ : CascadeMux
    port map (
            O => \N__35567\,
            I => \N__35555\
        );

    \I__7076\ : LocalMux
    port map (
            O => \N__35564\,
            I => \N__35552\
        );

    \I__7075\ : InMux
    port map (
            O => \N__35563\,
            I => \N__35549\
        );

    \I__7074\ : InMux
    port map (
            O => \N__35560\,
            I => \N__35546\
        );

    \I__7073\ : InMux
    port map (
            O => \N__35559\,
            I => \N__35543\
        );

    \I__7072\ : InMux
    port map (
            O => \N__35558\,
            I => \N__35540\
        );

    \I__7071\ : InMux
    port map (
            O => \N__35555\,
            I => \N__35537\
        );

    \I__7070\ : Span4Mux_v
    port map (
            O => \N__35552\,
            I => \N__35534\
        );

    \I__7069\ : LocalMux
    port map (
            O => \N__35549\,
            I => \N__35531\
        );

    \I__7068\ : LocalMux
    port map (
            O => \N__35546\,
            I => \N__35525\
        );

    \I__7067\ : LocalMux
    port map (
            O => \N__35543\,
            I => \N__35525\
        );

    \I__7066\ : LocalMux
    port map (
            O => \N__35540\,
            I => \N__35522\
        );

    \I__7065\ : LocalMux
    port map (
            O => \N__35537\,
            I => \N__35519\
        );

    \I__7064\ : Span4Mux_v
    port map (
            O => \N__35534\,
            I => \N__35514\
        );

    \I__7063\ : Span4Mux_h
    port map (
            O => \N__35531\,
            I => \N__35514\
        );

    \I__7062\ : InMux
    port map (
            O => \N__35530\,
            I => \N__35511\
        );

    \I__7061\ : Span4Mux_v
    port map (
            O => \N__35525\,
            I => \N__35502\
        );

    \I__7060\ : Span4Mux_h
    port map (
            O => \N__35522\,
            I => \N__35502\
        );

    \I__7059\ : Span4Mux_v
    port map (
            O => \N__35519\,
            I => \N__35502\
        );

    \I__7058\ : Span4Mux_h
    port map (
            O => \N__35514\,
            I => \N__35497\
        );

    \I__7057\ : LocalMux
    port map (
            O => \N__35511\,
            I => \N__35497\
        );

    \I__7056\ : InMux
    port map (
            O => \N__35510\,
            I => \N__35494\
        );

    \I__7055\ : InMux
    port map (
            O => \N__35509\,
            I => \N__35491\
        );

    \I__7054\ : Odrv4
    port map (
            O => \N__35502\,
            I => comm_rx_buf_3
        );

    \I__7053\ : Odrv4
    port map (
            O => \N__35497\,
            I => comm_rx_buf_3
        );

    \I__7052\ : LocalMux
    port map (
            O => \N__35494\,
            I => comm_rx_buf_3
        );

    \I__7051\ : LocalMux
    port map (
            O => \N__35491\,
            I => comm_rx_buf_3
        );

    \I__7050\ : InMux
    port map (
            O => \N__35482\,
            I => \N__35479\
        );

    \I__7049\ : LocalMux
    port map (
            O => \N__35479\,
            I => \N__35476\
        );

    \I__7048\ : Span4Mux_h
    port map (
            O => \N__35476\,
            I => \N__35473\
        );

    \I__7047\ : Span4Mux_v
    port map (
            O => \N__35473\,
            I => \N__35470\
        );

    \I__7046\ : Span4Mux_h
    port map (
            O => \N__35470\,
            I => \N__35467\
        );

    \I__7045\ : Span4Mux_h
    port map (
            O => \N__35467\,
            I => \N__35464\
        );

    \I__7044\ : Odrv4
    port map (
            O => \N__35464\,
            I => buf_data_vac_3
        );

    \I__7043\ : InMux
    port map (
            O => \N__35461\,
            I => \N__35458\
        );

    \I__7042\ : LocalMux
    port map (
            O => \N__35458\,
            I => \N__35455\
        );

    \I__7041\ : Odrv4
    port map (
            O => \N__35455\,
            I => comm_buf_5_3
        );

    \I__7040\ : InMux
    port map (
            O => \N__35452\,
            I => \N__35445\
        );

    \I__7039\ : InMux
    port map (
            O => \N__35451\,
            I => \N__35442\
        );

    \I__7038\ : InMux
    port map (
            O => \N__35450\,
            I => \N__35438\
        );

    \I__7037\ : InMux
    port map (
            O => \N__35449\,
            I => \N__35433\
        );

    \I__7036\ : InMux
    port map (
            O => \N__35448\,
            I => \N__35433\
        );

    \I__7035\ : LocalMux
    port map (
            O => \N__35445\,
            I => \N__35428\
        );

    \I__7034\ : LocalMux
    port map (
            O => \N__35442\,
            I => \N__35428\
        );

    \I__7033\ : InMux
    port map (
            O => \N__35441\,
            I => \N__35425\
        );

    \I__7032\ : LocalMux
    port map (
            O => \N__35438\,
            I => \N__35422\
        );

    \I__7031\ : LocalMux
    port map (
            O => \N__35433\,
            I => \N__35417\
        );

    \I__7030\ : Span4Mux_v
    port map (
            O => \N__35428\,
            I => \N__35414\
        );

    \I__7029\ : LocalMux
    port map (
            O => \N__35425\,
            I => \N__35411\
        );

    \I__7028\ : Span4Mux_v
    port map (
            O => \N__35422\,
            I => \N__35408\
        );

    \I__7027\ : InMux
    port map (
            O => \N__35421\,
            I => \N__35405\
        );

    \I__7026\ : CascadeMux
    port map (
            O => \N__35420\,
            I => \N__35402\
        );

    \I__7025\ : Span4Mux_v
    port map (
            O => \N__35417\,
            I => \N__35398\
        );

    \I__7024\ : Sp12to4
    port map (
            O => \N__35414\,
            I => \N__35395\
        );

    \I__7023\ : Span4Mux_h
    port map (
            O => \N__35411\,
            I => \N__35392\
        );

    \I__7022\ : Span4Mux_h
    port map (
            O => \N__35408\,
            I => \N__35387\
        );

    \I__7021\ : LocalMux
    port map (
            O => \N__35405\,
            I => \N__35387\
        );

    \I__7020\ : InMux
    port map (
            O => \N__35402\,
            I => \N__35384\
        );

    \I__7019\ : InMux
    port map (
            O => \N__35401\,
            I => \N__35381\
        );

    \I__7018\ : Odrv4
    port map (
            O => \N__35398\,
            I => comm_rx_buf_2
        );

    \I__7017\ : Odrv12
    port map (
            O => \N__35395\,
            I => comm_rx_buf_2
        );

    \I__7016\ : Odrv4
    port map (
            O => \N__35392\,
            I => comm_rx_buf_2
        );

    \I__7015\ : Odrv4
    port map (
            O => \N__35387\,
            I => comm_rx_buf_2
        );

    \I__7014\ : LocalMux
    port map (
            O => \N__35384\,
            I => comm_rx_buf_2
        );

    \I__7013\ : LocalMux
    port map (
            O => \N__35381\,
            I => comm_rx_buf_2
        );

    \I__7012\ : InMux
    port map (
            O => \N__35368\,
            I => \N__35365\
        );

    \I__7011\ : LocalMux
    port map (
            O => \N__35365\,
            I => \N__35362\
        );

    \I__7010\ : Span12Mux_v
    port map (
            O => \N__35362\,
            I => \N__35359\
        );

    \I__7009\ : Odrv12
    port map (
            O => \N__35359\,
            I => buf_data_vac_2
        );

    \I__7008\ : InMux
    port map (
            O => \N__35356\,
            I => \N__35353\
        );

    \I__7007\ : LocalMux
    port map (
            O => \N__35353\,
            I => \N__35350\
        );

    \I__7006\ : Odrv12
    port map (
            O => \N__35350\,
            I => comm_buf_5_2
        );

    \I__7005\ : InMux
    port map (
            O => \N__35347\,
            I => \N__35344\
        );

    \I__7004\ : LocalMux
    port map (
            O => \N__35344\,
            I => \N__35341\
        );

    \I__7003\ : Span12Mux_v
    port map (
            O => \N__35341\,
            I => \N__35338\
        );

    \I__7002\ : Odrv12
    port map (
            O => \N__35338\,
            I => buf_data_vac_1
        );

    \I__7001\ : InMux
    port map (
            O => \N__35335\,
            I => \N__35332\
        );

    \I__7000\ : LocalMux
    port map (
            O => \N__35332\,
            I => \N__35329\
        );

    \I__6999\ : Span4Mux_v
    port map (
            O => \N__35329\,
            I => \N__35326\
        );

    \I__6998\ : Span4Mux_h
    port map (
            O => \N__35326\,
            I => \N__35322\
        );

    \I__6997\ : CascadeMux
    port map (
            O => \N__35325\,
            I => \N__35319\
        );

    \I__6996\ : Span4Mux_h
    port map (
            O => \N__35322\,
            I => \N__35316\
        );

    \I__6995\ : InMux
    port map (
            O => \N__35319\,
            I => \N__35313\
        );

    \I__6994\ : Odrv4
    port map (
            O => \N__35316\,
            I => \buf_readRTD_1\
        );

    \I__6993\ : LocalMux
    port map (
            O => \N__35313\,
            I => \buf_readRTD_1\
        );

    \I__6992\ : InMux
    port map (
            O => \N__35308\,
            I => \N__35305\
        );

    \I__6991\ : LocalMux
    port map (
            O => \N__35305\,
            I => \N__35302\
        );

    \I__6990\ : Span4Mux_v
    port map (
            O => \N__35302\,
            I => \N__35298\
        );

    \I__6989\ : CascadeMux
    port map (
            O => \N__35301\,
            I => \N__35295\
        );

    \I__6988\ : Span4Mux_h
    port map (
            O => \N__35298\,
            I => \N__35292\
        );

    \I__6987\ : InMux
    port map (
            O => \N__35295\,
            I => \N__35289\
        );

    \I__6986\ : Odrv4
    port map (
            O => \N__35292\,
            I => buf_adcdata_vdc_9
        );

    \I__6985\ : LocalMux
    port map (
            O => \N__35289\,
            I => buf_adcdata_vdc_9
        );

    \I__6984\ : InMux
    port map (
            O => \N__35284\,
            I => \N__35280\
        );

    \I__6983\ : InMux
    port map (
            O => \N__35283\,
            I => \N__35277\
        );

    \I__6982\ : LocalMux
    port map (
            O => \N__35280\,
            I => \N__35273\
        );

    \I__6981\ : LocalMux
    port map (
            O => \N__35277\,
            I => \N__35270\
        );

    \I__6980\ : CascadeMux
    port map (
            O => \N__35276\,
            I => \N__35267\
        );

    \I__6979\ : Span4Mux_v
    port map (
            O => \N__35273\,
            I => \N__35264\
        );

    \I__6978\ : Span4Mux_v
    port map (
            O => \N__35270\,
            I => \N__35261\
        );

    \I__6977\ : InMux
    port map (
            O => \N__35267\,
            I => \N__35258\
        );

    \I__6976\ : Span4Mux_h
    port map (
            O => \N__35264\,
            I => \N__35255\
        );

    \I__6975\ : Span4Mux_h
    port map (
            O => \N__35261\,
            I => \N__35252\
        );

    \I__6974\ : LocalMux
    port map (
            O => \N__35258\,
            I => buf_adcdata_vac_9
        );

    \I__6973\ : Odrv4
    port map (
            O => \N__35255\,
            I => buf_adcdata_vac_9
        );

    \I__6972\ : Odrv4
    port map (
            O => \N__35252\,
            I => buf_adcdata_vac_9
        );

    \I__6971\ : InMux
    port map (
            O => \N__35245\,
            I => \N__35242\
        );

    \I__6970\ : LocalMux
    port map (
            O => \N__35242\,
            I => n19_adj_1508
        );

    \I__6969\ : InMux
    port map (
            O => \N__35239\,
            I => \N__35236\
        );

    \I__6968\ : LocalMux
    port map (
            O => \N__35236\,
            I => \N__35233\
        );

    \I__6967\ : Odrv12
    port map (
            O => \N__35233\,
            I => n30_adj_1475
        );

    \I__6966\ : InMux
    port map (
            O => \N__35230\,
            I => \N__35227\
        );

    \I__6965\ : LocalMux
    port map (
            O => \N__35227\,
            I => \N__35224\
        );

    \I__6964\ : Odrv12
    port map (
            O => \N__35224\,
            I => comm_buf_2_7
        );

    \I__6963\ : InMux
    port map (
            O => \N__35221\,
            I => \N__35218\
        );

    \I__6962\ : LocalMux
    port map (
            O => \N__35218\,
            I => \N__35215\
        );

    \I__6961\ : Odrv4
    port map (
            O => \N__35215\,
            I => n30_adj_1595
        );

    \I__6960\ : InMux
    port map (
            O => \N__35212\,
            I => \N__35209\
        );

    \I__6959\ : LocalMux
    port map (
            O => \N__35209\,
            I => \N__35206\
        );

    \I__6958\ : Odrv4
    port map (
            O => \N__35206\,
            I => comm_buf_2_6
        );

    \I__6957\ : InMux
    port map (
            O => \N__35203\,
            I => \N__35200\
        );

    \I__6956\ : LocalMux
    port map (
            O => \N__35200\,
            I => \N__35197\
        );

    \I__6955\ : Span12Mux_h
    port map (
            O => \N__35197\,
            I => \N__35194\
        );

    \I__6954\ : Odrv12
    port map (
            O => \N__35194\,
            I => n30_adj_1612
        );

    \I__6953\ : InMux
    port map (
            O => \N__35191\,
            I => \N__35188\
        );

    \I__6952\ : LocalMux
    port map (
            O => \N__35188\,
            I => comm_buf_2_3
        );

    \I__6951\ : InMux
    port map (
            O => \N__35185\,
            I => \N__35182\
        );

    \I__6950\ : LocalMux
    port map (
            O => \N__35182\,
            I => \N__35179\
        );

    \I__6949\ : Span12Mux_h
    port map (
            O => \N__35179\,
            I => \N__35176\
        );

    \I__6948\ : Odrv12
    port map (
            O => \N__35176\,
            I => n30_adj_1615
        );

    \I__6947\ : InMux
    port map (
            O => \N__35173\,
            I => \N__35170\
        );

    \I__6946\ : LocalMux
    port map (
            O => \N__35170\,
            I => \N__35167\
        );

    \I__6945\ : Odrv4
    port map (
            O => \N__35167\,
            I => comm_buf_2_2
        );

    \I__6944\ : InMux
    port map (
            O => \N__35164\,
            I => \N__35161\
        );

    \I__6943\ : LocalMux
    port map (
            O => \N__35161\,
            I => \N__35158\
        );

    \I__6942\ : Span4Mux_v
    port map (
            O => \N__35158\,
            I => \N__35155\
        );

    \I__6941\ : Span4Mux_h
    port map (
            O => \N__35155\,
            I => \N__35152\
        );

    \I__6940\ : Odrv4
    port map (
            O => \N__35152\,
            I => n30_adj_1619
        );

    \I__6939\ : InMux
    port map (
            O => \N__35149\,
            I => \N__35146\
        );

    \I__6938\ : LocalMux
    port map (
            O => \N__35146\,
            I => comm_buf_2_1
        );

    \I__6937\ : InMux
    port map (
            O => \N__35143\,
            I => \N__35140\
        );

    \I__6936\ : LocalMux
    port map (
            O => \N__35140\,
            I => \N__35137\
        );

    \I__6935\ : Span12Mux_v
    port map (
            O => \N__35137\,
            I => \N__35134\
        );

    \I__6934\ : Odrv12
    port map (
            O => \N__35134\,
            I => buf_data_vac_0
        );

    \I__6933\ : InMux
    port map (
            O => \N__35131\,
            I => \N__35128\
        );

    \I__6932\ : LocalMux
    port map (
            O => \N__35128\,
            I => \N__35125\
        );

    \I__6931\ : Span4Mux_h
    port map (
            O => \N__35125\,
            I => \N__35122\
        );

    \I__6930\ : Odrv4
    port map (
            O => \N__35122\,
            I => comm_buf_5_0
        );

    \I__6929\ : InMux
    port map (
            O => \N__35119\,
            I => \N__35116\
        );

    \I__6928\ : LocalMux
    port map (
            O => \N__35116\,
            I => \N__35113\
        );

    \I__6927\ : Odrv12
    port map (
            O => \N__35113\,
            I => buf_data_vac_7
        );

    \I__6926\ : InMux
    port map (
            O => \N__35110\,
            I => \N__35107\
        );

    \I__6925\ : LocalMux
    port map (
            O => \N__35107\,
            I => \N__35104\
        );

    \I__6924\ : Span4Mux_h
    port map (
            O => \N__35104\,
            I => \N__35101\
        );

    \I__6923\ : Odrv4
    port map (
            O => \N__35101\,
            I => comm_buf_5_7
        );

    \I__6922\ : InMux
    port map (
            O => \N__35098\,
            I => \N__35095\
        );

    \I__6921\ : LocalMux
    port map (
            O => \N__35095\,
            I => \N__35092\
        );

    \I__6920\ : Span4Mux_h
    port map (
            O => \N__35092\,
            I => \N__35089\
        );

    \I__6919\ : Odrv4
    port map (
            O => \N__35089\,
            I => comm_buf_4_2
        );

    \I__6918\ : InMux
    port map (
            O => \N__35086\,
            I => \N__35083\
        );

    \I__6917\ : LocalMux
    port map (
            O => \N__35083\,
            I => \N__35079\
        );

    \I__6916\ : InMux
    port map (
            O => \N__35082\,
            I => \N__35076\
        );

    \I__6915\ : Span4Mux_v
    port map (
            O => \N__35079\,
            I => \N__35073\
        );

    \I__6914\ : LocalMux
    port map (
            O => \N__35076\,
            I => \N__35070\
        );

    \I__6913\ : Span4Mux_h
    port map (
            O => \N__35073\,
            I => \N__35067\
        );

    \I__6912\ : Odrv4
    port map (
            O => \N__35070\,
            I => comm_buf_6_2
        );

    \I__6911\ : Odrv4
    port map (
            O => \N__35067\,
            I => comm_buf_6_2
        );

    \I__6910\ : CascadeMux
    port map (
            O => \N__35062\,
            I => \n4_adj_1568_cascade_\
        );

    \I__6909\ : InMux
    port map (
            O => \N__35059\,
            I => \N__35056\
        );

    \I__6908\ : LocalMux
    port map (
            O => \N__35056\,
            I => n20786
        );

    \I__6907\ : InMux
    port map (
            O => \N__35053\,
            I => \N__35050\
        );

    \I__6906\ : LocalMux
    port map (
            O => \N__35050\,
            I => n4_adj_1560
        );

    \I__6905\ : CascadeMux
    port map (
            O => \N__35047\,
            I => \n21276_cascade_\
        );

    \I__6904\ : InMux
    port map (
            O => \N__35044\,
            I => \N__35041\
        );

    \I__6903\ : LocalMux
    port map (
            O => \N__35041\,
            I => n22105
        );

    \I__6902\ : InMux
    port map (
            O => \N__35038\,
            I => \N__35035\
        );

    \I__6901\ : LocalMux
    port map (
            O => \N__35035\,
            I => \N__35032\
        );

    \I__6900\ : Span4Mux_h
    port map (
            O => \N__35032\,
            I => \N__35029\
        );

    \I__6899\ : Odrv4
    port map (
            O => \N__35029\,
            I => comm_buf_3_2
        );

    \I__6898\ : CascadeMux
    port map (
            O => \N__35026\,
            I => \n21985_cascade_\
        );

    \I__6897\ : CascadeMux
    port map (
            O => \N__35023\,
            I => \n21988_cascade_\
        );

    \I__6896\ : InMux
    port map (
            O => \N__35020\,
            I => \N__35017\
        );

    \I__6895\ : LocalMux
    port map (
            O => \N__35017\,
            I => \N__35014\
        );

    \I__6894\ : Span4Mux_v
    port map (
            O => \N__35014\,
            I => \N__35011\
        );

    \I__6893\ : Odrv4
    port map (
            O => \N__35011\,
            I => comm_buf_3_0
        );

    \I__6892\ : CascadeMux
    port map (
            O => \N__35008\,
            I => \n17304_cascade_\
        );

    \I__6891\ : CascadeMux
    port map (
            O => \N__35005\,
            I => \n20906_cascade_\
        );

    \I__6890\ : InMux
    port map (
            O => \N__35002\,
            I => \N__34999\
        );

    \I__6889\ : LocalMux
    port map (
            O => \N__34999\,
            I => \ADC_VDC.genclk.n27_adj_1402\
        );

    \I__6888\ : InMux
    port map (
            O => \N__34996\,
            I => \N__34991\
        );

    \I__6887\ : InMux
    port map (
            O => \N__34995\,
            I => \N__34988\
        );

    \I__6886\ : InMux
    port map (
            O => \N__34994\,
            I => \N__34985\
        );

    \I__6885\ : LocalMux
    port map (
            O => \N__34991\,
            I => \N__34980\
        );

    \I__6884\ : LocalMux
    port map (
            O => \N__34988\,
            I => \N__34980\
        );

    \I__6883\ : LocalMux
    port map (
            O => \N__34985\,
            I => \comm_spi.n14586\
        );

    \I__6882\ : Odrv4
    port map (
            O => \N__34980\,
            I => \comm_spi.n14586\
        );

    \I__6881\ : CascadeMux
    port map (
            O => \N__34975\,
            I => \N__34971\
        );

    \I__6880\ : InMux
    port map (
            O => \N__34974\,
            I => \N__34967\
        );

    \I__6879\ : InMux
    port map (
            O => \N__34971\,
            I => \N__34964\
        );

    \I__6878\ : InMux
    port map (
            O => \N__34970\,
            I => \N__34959\
        );

    \I__6877\ : LocalMux
    port map (
            O => \N__34967\,
            I => \N__34956\
        );

    \I__6876\ : LocalMux
    port map (
            O => \N__34964\,
            I => \N__34953\
        );

    \I__6875\ : InMux
    port map (
            O => \N__34963\,
            I => \N__34950\
        );

    \I__6874\ : InMux
    port map (
            O => \N__34962\,
            I => \N__34947\
        );

    \I__6873\ : LocalMux
    port map (
            O => \N__34959\,
            I => \ADC_VDC.genclk.div_state_0\
        );

    \I__6872\ : Odrv4
    port map (
            O => \N__34956\,
            I => \ADC_VDC.genclk.div_state_0\
        );

    \I__6871\ : Odrv12
    port map (
            O => \N__34953\,
            I => \ADC_VDC.genclk.div_state_0\
        );

    \I__6870\ : LocalMux
    port map (
            O => \N__34950\,
            I => \ADC_VDC.genclk.div_state_0\
        );

    \I__6869\ : LocalMux
    port map (
            O => \N__34947\,
            I => \ADC_VDC.genclk.div_state_0\
        );

    \I__6868\ : CascadeMux
    port map (
            O => \N__34936\,
            I => \N__34932\
        );

    \I__6867\ : InMux
    port map (
            O => \N__34935\,
            I => \N__34927\
        );

    \I__6866\ : InMux
    port map (
            O => \N__34932\,
            I => \N__34922\
        );

    \I__6865\ : InMux
    port map (
            O => \N__34931\,
            I => \N__34922\
        );

    \I__6864\ : InMux
    port map (
            O => \N__34930\,
            I => \N__34919\
        );

    \I__6863\ : LocalMux
    port map (
            O => \N__34927\,
            I => \N__34915\
        );

    \I__6862\ : LocalMux
    port map (
            O => \N__34922\,
            I => \N__34908\
        );

    \I__6861\ : LocalMux
    port map (
            O => \N__34919\,
            I => \N__34908\
        );

    \I__6860\ : InMux
    port map (
            O => \N__34918\,
            I => \N__34905\
        );

    \I__6859\ : Span4Mux_h
    port map (
            O => \N__34915\,
            I => \N__34902\
        );

    \I__6858\ : InMux
    port map (
            O => \N__34914\,
            I => \N__34897\
        );

    \I__6857\ : InMux
    port map (
            O => \N__34913\,
            I => \N__34897\
        );

    \I__6856\ : Span4Mux_h
    port map (
            O => \N__34908\,
            I => \N__34894\
        );

    \I__6855\ : LocalMux
    port map (
            O => \N__34905\,
            I => \ADC_VDC.genclk.div_state_1\
        );

    \I__6854\ : Odrv4
    port map (
            O => \N__34902\,
            I => \ADC_VDC.genclk.div_state_1\
        );

    \I__6853\ : LocalMux
    port map (
            O => \N__34897\,
            I => \ADC_VDC.genclk.div_state_1\
        );

    \I__6852\ : Odrv4
    port map (
            O => \N__34894\,
            I => \ADC_VDC.genclk.div_state_1\
        );

    \I__6851\ : CEMux
    port map (
            O => \N__34885\,
            I => \N__34882\
        );

    \I__6850\ : LocalMux
    port map (
            O => \N__34882\,
            I => \ADC_VDC.genclk.n6\
        );

    \I__6849\ : CascadeMux
    port map (
            O => \N__34879\,
            I => \N__34873\
        );

    \I__6848\ : CascadeMux
    port map (
            O => \N__34878\,
            I => \N__34869\
        );

    \I__6847\ : CascadeMux
    port map (
            O => \N__34877\,
            I => \N__34866\
        );

    \I__6846\ : InMux
    port map (
            O => \N__34876\,
            I => \N__34861\
        );

    \I__6845\ : InMux
    port map (
            O => \N__34873\,
            I => \N__34858\
        );

    \I__6844\ : InMux
    port map (
            O => \N__34872\,
            I => \N__34855\
        );

    \I__6843\ : InMux
    port map (
            O => \N__34869\,
            I => \N__34850\
        );

    \I__6842\ : InMux
    port map (
            O => \N__34866\,
            I => \N__34850\
        );

    \I__6841\ : InMux
    port map (
            O => \N__34865\,
            I => \N__34847\
        );

    \I__6840\ : CascadeMux
    port map (
            O => \N__34864\,
            I => \N__34841\
        );

    \I__6839\ : LocalMux
    port map (
            O => \N__34861\,
            I => \N__34838\
        );

    \I__6838\ : LocalMux
    port map (
            O => \N__34858\,
            I => \N__34835\
        );

    \I__6837\ : LocalMux
    port map (
            O => \N__34855\,
            I => \N__34832\
        );

    \I__6836\ : LocalMux
    port map (
            O => \N__34850\,
            I => \N__34827\
        );

    \I__6835\ : LocalMux
    port map (
            O => \N__34847\,
            I => \N__34827\
        );

    \I__6834\ : InMux
    port map (
            O => \N__34846\,
            I => \N__34820\
        );

    \I__6833\ : InMux
    port map (
            O => \N__34845\,
            I => \N__34820\
        );

    \I__6832\ : InMux
    port map (
            O => \N__34844\,
            I => \N__34820\
        );

    \I__6831\ : InMux
    port map (
            O => \N__34841\,
            I => \N__34817\
        );

    \I__6830\ : Span4Mux_v
    port map (
            O => \N__34838\,
            I => \N__34812\
        );

    \I__6829\ : Span4Mux_v
    port map (
            O => \N__34835\,
            I => \N__34812\
        );

    \I__6828\ : Span4Mux_h
    port map (
            O => \N__34832\,
            I => \N__34805\
        );

    \I__6827\ : Span4Mux_v
    port map (
            O => \N__34827\,
            I => \N__34805\
        );

    \I__6826\ : LocalMux
    port map (
            O => \N__34820\,
            I => \N__34805\
        );

    \I__6825\ : LocalMux
    port map (
            O => \N__34817\,
            I => \N__34802\
        );

    \I__6824\ : Span4Mux_v
    port map (
            O => \N__34812\,
            I => \N__34799\
        );

    \I__6823\ : Span4Mux_h
    port map (
            O => \N__34805\,
            I => \N__34796\
        );

    \I__6822\ : Span12Mux_v
    port map (
            O => \N__34802\,
            I => \N__34793\
        );

    \I__6821\ : Span4Mux_h
    port map (
            O => \N__34799\,
            I => \N__34790\
        );

    \I__6820\ : Span4Mux_v
    port map (
            O => \N__34796\,
            I => \N__34787\
        );

    \I__6819\ : Span12Mux_h
    port map (
            O => \N__34793\,
            I => \N__34784\
        );

    \I__6818\ : Sp12to4
    port map (
            O => \N__34790\,
            I => \N__34779\
        );

    \I__6817\ : Sp12to4
    port map (
            O => \N__34787\,
            I => \N__34779\
        );

    \I__6816\ : Odrv12
    port map (
            O => \N__34784\,
            I => \VDC_SDO\
        );

    \I__6815\ : Odrv12
    port map (
            O => \N__34779\,
            I => \VDC_SDO\
        );

    \I__6814\ : InMux
    port map (
            O => \N__34774\,
            I => \N__34765\
        );

    \I__6813\ : InMux
    port map (
            O => \N__34773\,
            I => \N__34762\
        );

    \I__6812\ : InMux
    port map (
            O => \N__34772\,
            I => \N__34755\
        );

    \I__6811\ : InMux
    port map (
            O => \N__34771\,
            I => \N__34755\
        );

    \I__6810\ : InMux
    port map (
            O => \N__34770\,
            I => \N__34755\
        );

    \I__6809\ : InMux
    port map (
            O => \N__34769\,
            I => \N__34752\
        );

    \I__6808\ : CascadeMux
    port map (
            O => \N__34768\,
            I => \N__34748\
        );

    \I__6807\ : LocalMux
    port map (
            O => \N__34765\,
            I => \N__34736\
        );

    \I__6806\ : LocalMux
    port map (
            O => \N__34762\,
            I => \N__34731\
        );

    \I__6805\ : LocalMux
    port map (
            O => \N__34755\,
            I => \N__34731\
        );

    \I__6804\ : LocalMux
    port map (
            O => \N__34752\,
            I => \N__34728\
        );

    \I__6803\ : CascadeMux
    port map (
            O => \N__34751\,
            I => \N__34725\
        );

    \I__6802\ : InMux
    port map (
            O => \N__34748\,
            I => \N__34720\
        );

    \I__6801\ : InMux
    port map (
            O => \N__34747\,
            I => \N__34717\
        );

    \I__6800\ : CascadeMux
    port map (
            O => \N__34746\,
            I => \N__34713\
        );

    \I__6799\ : InMux
    port map (
            O => \N__34745\,
            I => \N__34709\
        );

    \I__6798\ : InMux
    port map (
            O => \N__34744\,
            I => \N__34704\
        );

    \I__6797\ : InMux
    port map (
            O => \N__34743\,
            I => \N__34704\
        );

    \I__6796\ : InMux
    port map (
            O => \N__34742\,
            I => \N__34701\
        );

    \I__6795\ : InMux
    port map (
            O => \N__34741\,
            I => \N__34698\
        );

    \I__6794\ : InMux
    port map (
            O => \N__34740\,
            I => \N__34693\
        );

    \I__6793\ : InMux
    port map (
            O => \N__34739\,
            I => \N__34693\
        );

    \I__6792\ : Span4Mux_v
    port map (
            O => \N__34736\,
            I => \N__34686\
        );

    \I__6791\ : Span4Mux_v
    port map (
            O => \N__34731\,
            I => \N__34686\
        );

    \I__6790\ : Span4Mux_v
    port map (
            O => \N__34728\,
            I => \N__34686\
        );

    \I__6789\ : InMux
    port map (
            O => \N__34725\,
            I => \N__34679\
        );

    \I__6788\ : InMux
    port map (
            O => \N__34724\,
            I => \N__34679\
        );

    \I__6787\ : InMux
    port map (
            O => \N__34723\,
            I => \N__34679\
        );

    \I__6786\ : LocalMux
    port map (
            O => \N__34720\,
            I => \N__34674\
        );

    \I__6785\ : LocalMux
    port map (
            O => \N__34717\,
            I => \N__34674\
        );

    \I__6784\ : InMux
    port map (
            O => \N__34716\,
            I => \N__34667\
        );

    \I__6783\ : InMux
    port map (
            O => \N__34713\,
            I => \N__34667\
        );

    \I__6782\ : InMux
    port map (
            O => \N__34712\,
            I => \N__34667\
        );

    \I__6781\ : LocalMux
    port map (
            O => \N__34709\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__6780\ : LocalMux
    port map (
            O => \N__34704\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__6779\ : LocalMux
    port map (
            O => \N__34701\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__6778\ : LocalMux
    port map (
            O => \N__34698\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__6777\ : LocalMux
    port map (
            O => \N__34693\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__6776\ : Odrv4
    port map (
            O => \N__34686\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__6775\ : LocalMux
    port map (
            O => \N__34679\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__6774\ : Odrv4
    port map (
            O => \N__34674\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__6773\ : LocalMux
    port map (
            O => \N__34667\,
            I => \ADC_VDC.adc_state_0\
        );

    \I__6772\ : InMux
    port map (
            O => \N__34648\,
            I => \N__34645\
        );

    \I__6771\ : LocalMux
    port map (
            O => \N__34645\,
            I => \ADC_VDC.n62\
        );

    \I__6770\ : CascadeMux
    port map (
            O => \N__34642\,
            I => \N__34621\
        );

    \I__6769\ : InMux
    port map (
            O => \N__34641\,
            I => \N__34617\
        );

    \I__6768\ : InMux
    port map (
            O => \N__34640\,
            I => \N__34602\
        );

    \I__6767\ : InMux
    port map (
            O => \N__34639\,
            I => \N__34602\
        );

    \I__6766\ : InMux
    port map (
            O => \N__34638\,
            I => \N__34602\
        );

    \I__6765\ : InMux
    port map (
            O => \N__34637\,
            I => \N__34602\
        );

    \I__6764\ : InMux
    port map (
            O => \N__34636\,
            I => \N__34602\
        );

    \I__6763\ : InMux
    port map (
            O => \N__34635\,
            I => \N__34602\
        );

    \I__6762\ : InMux
    port map (
            O => \N__34634\,
            I => \N__34602\
        );

    \I__6761\ : InMux
    port map (
            O => \N__34633\,
            I => \N__34595\
        );

    \I__6760\ : InMux
    port map (
            O => \N__34632\,
            I => \N__34595\
        );

    \I__6759\ : InMux
    port map (
            O => \N__34631\,
            I => \N__34595\
        );

    \I__6758\ : CascadeMux
    port map (
            O => \N__34630\,
            I => \N__34590\
        );

    \I__6757\ : InMux
    port map (
            O => \N__34629\,
            I => \N__34585\
        );

    \I__6756\ : InMux
    port map (
            O => \N__34628\,
            I => \N__34575\
        );

    \I__6755\ : InMux
    port map (
            O => \N__34627\,
            I => \N__34575\
        );

    \I__6754\ : InMux
    port map (
            O => \N__34626\,
            I => \N__34575\
        );

    \I__6753\ : InMux
    port map (
            O => \N__34625\,
            I => \N__34575\
        );

    \I__6752\ : InMux
    port map (
            O => \N__34624\,
            I => \N__34556\
        );

    \I__6751\ : InMux
    port map (
            O => \N__34621\,
            I => \N__34556\
        );

    \I__6750\ : CascadeMux
    port map (
            O => \N__34620\,
            I => \N__34553\
        );

    \I__6749\ : LocalMux
    port map (
            O => \N__34617\,
            I => \N__34546\
        );

    \I__6748\ : LocalMux
    port map (
            O => \N__34602\,
            I => \N__34546\
        );

    \I__6747\ : LocalMux
    port map (
            O => \N__34595\,
            I => \N__34546\
        );

    \I__6746\ : InMux
    port map (
            O => \N__34594\,
            I => \N__34541\
        );

    \I__6745\ : InMux
    port map (
            O => \N__34593\,
            I => \N__34541\
        );

    \I__6744\ : InMux
    port map (
            O => \N__34590\,
            I => \N__34536\
        );

    \I__6743\ : InMux
    port map (
            O => \N__34589\,
            I => \N__34536\
        );

    \I__6742\ : InMux
    port map (
            O => \N__34588\,
            I => \N__34533\
        );

    \I__6741\ : LocalMux
    port map (
            O => \N__34585\,
            I => \N__34530\
        );

    \I__6740\ : InMux
    port map (
            O => \N__34584\,
            I => \N__34527\
        );

    \I__6739\ : LocalMux
    port map (
            O => \N__34575\,
            I => \N__34524\
        );

    \I__6738\ : InMux
    port map (
            O => \N__34574\,
            I => \N__34507\
        );

    \I__6737\ : InMux
    port map (
            O => \N__34573\,
            I => \N__34507\
        );

    \I__6736\ : InMux
    port map (
            O => \N__34572\,
            I => \N__34507\
        );

    \I__6735\ : InMux
    port map (
            O => \N__34571\,
            I => \N__34507\
        );

    \I__6734\ : InMux
    port map (
            O => \N__34570\,
            I => \N__34507\
        );

    \I__6733\ : InMux
    port map (
            O => \N__34569\,
            I => \N__34507\
        );

    \I__6732\ : InMux
    port map (
            O => \N__34568\,
            I => \N__34507\
        );

    \I__6731\ : InMux
    port map (
            O => \N__34567\,
            I => \N__34507\
        );

    \I__6730\ : InMux
    port map (
            O => \N__34566\,
            I => \N__34504\
        );

    \I__6729\ : CascadeMux
    port map (
            O => \N__34565\,
            I => \N__34500\
        );

    \I__6728\ : CascadeMux
    port map (
            O => \N__34564\,
            I => \N__34497\
        );

    \I__6727\ : CascadeMux
    port map (
            O => \N__34563\,
            I => \N__34494\
        );

    \I__6726\ : CascadeMux
    port map (
            O => \N__34562\,
            I => \N__34491\
        );

    \I__6725\ : CascadeMux
    port map (
            O => \N__34561\,
            I => \N__34482\
        );

    \I__6724\ : LocalMux
    port map (
            O => \N__34556\,
            I => \N__34479\
        );

    \I__6723\ : InMux
    port map (
            O => \N__34553\,
            I => \N__34476\
        );

    \I__6722\ : Span4Mux_v
    port map (
            O => \N__34546\,
            I => \N__34467\
        );

    \I__6721\ : LocalMux
    port map (
            O => \N__34541\,
            I => \N__34467\
        );

    \I__6720\ : LocalMux
    port map (
            O => \N__34536\,
            I => \N__34467\
        );

    \I__6719\ : LocalMux
    port map (
            O => \N__34533\,
            I => \N__34467\
        );

    \I__6718\ : Span4Mux_h
    port map (
            O => \N__34530\,
            I => \N__34456\
        );

    \I__6717\ : LocalMux
    port map (
            O => \N__34527\,
            I => \N__34456\
        );

    \I__6716\ : Span4Mux_h
    port map (
            O => \N__34524\,
            I => \N__34456\
        );

    \I__6715\ : LocalMux
    port map (
            O => \N__34507\,
            I => \N__34456\
        );

    \I__6714\ : LocalMux
    port map (
            O => \N__34504\,
            I => \N__34453\
        );

    \I__6713\ : InMux
    port map (
            O => \N__34503\,
            I => \N__34446\
        );

    \I__6712\ : InMux
    port map (
            O => \N__34500\,
            I => \N__34446\
        );

    \I__6711\ : InMux
    port map (
            O => \N__34497\,
            I => \N__34446\
        );

    \I__6710\ : InMux
    port map (
            O => \N__34494\,
            I => \N__34443\
        );

    \I__6709\ : InMux
    port map (
            O => \N__34491\,
            I => \N__34436\
        );

    \I__6708\ : InMux
    port map (
            O => \N__34490\,
            I => \N__34436\
        );

    \I__6707\ : InMux
    port map (
            O => \N__34489\,
            I => \N__34436\
        );

    \I__6706\ : InMux
    port map (
            O => \N__34488\,
            I => \N__34425\
        );

    \I__6705\ : InMux
    port map (
            O => \N__34487\,
            I => \N__34425\
        );

    \I__6704\ : InMux
    port map (
            O => \N__34486\,
            I => \N__34425\
        );

    \I__6703\ : InMux
    port map (
            O => \N__34485\,
            I => \N__34425\
        );

    \I__6702\ : InMux
    port map (
            O => \N__34482\,
            I => \N__34425\
        );

    \I__6701\ : Span4Mux_h
    port map (
            O => \N__34479\,
            I => \N__34418\
        );

    \I__6700\ : LocalMux
    port map (
            O => \N__34476\,
            I => \N__34418\
        );

    \I__6699\ : Span4Mux_h
    port map (
            O => \N__34467\,
            I => \N__34418\
        );

    \I__6698\ : InMux
    port map (
            O => \N__34466\,
            I => \N__34413\
        );

    \I__6697\ : InMux
    port map (
            O => \N__34465\,
            I => \N__34413\
        );

    \I__6696\ : Span4Mux_v
    port map (
            O => \N__34456\,
            I => \N__34406\
        );

    \I__6695\ : Span4Mux_v
    port map (
            O => \N__34453\,
            I => \N__34406\
        );

    \I__6694\ : LocalMux
    port map (
            O => \N__34446\,
            I => \N__34406\
        );

    \I__6693\ : LocalMux
    port map (
            O => \N__34443\,
            I => adc_state_2
        );

    \I__6692\ : LocalMux
    port map (
            O => \N__34436\,
            I => adc_state_2
        );

    \I__6691\ : LocalMux
    port map (
            O => \N__34425\,
            I => adc_state_2
        );

    \I__6690\ : Odrv4
    port map (
            O => \N__34418\,
            I => adc_state_2
        );

    \I__6689\ : LocalMux
    port map (
            O => \N__34413\,
            I => adc_state_2
        );

    \I__6688\ : Odrv4
    port map (
            O => \N__34406\,
            I => adc_state_2
        );

    \I__6687\ : CascadeMux
    port map (
            O => \N__34393\,
            I => \N__34390\
        );

    \I__6686\ : InMux
    port map (
            O => \N__34390\,
            I => \N__34387\
        );

    \I__6685\ : LocalMux
    port map (
            O => \N__34387\,
            I => \N__34381\
        );

    \I__6684\ : InMux
    port map (
            O => \N__34386\,
            I => \N__34376\
        );

    \I__6683\ : InMux
    port map (
            O => \N__34385\,
            I => \N__34376\
        );

    \I__6682\ : CascadeMux
    port map (
            O => \N__34384\,
            I => \N__34357\
        );

    \I__6681\ : Span4Mux_h
    port map (
            O => \N__34381\,
            I => \N__34350\
        );

    \I__6680\ : LocalMux
    port map (
            O => \N__34376\,
            I => \N__34350\
        );

    \I__6679\ : InMux
    port map (
            O => \N__34375\,
            I => \N__34347\
        );

    \I__6678\ : InMux
    port map (
            O => \N__34374\,
            I => \N__34336\
        );

    \I__6677\ : InMux
    port map (
            O => \N__34373\,
            I => \N__34336\
        );

    \I__6676\ : InMux
    port map (
            O => \N__34372\,
            I => \N__34336\
        );

    \I__6675\ : InMux
    port map (
            O => \N__34371\,
            I => \N__34336\
        );

    \I__6674\ : InMux
    port map (
            O => \N__34370\,
            I => \N__34336\
        );

    \I__6673\ : InMux
    port map (
            O => \N__34369\,
            I => \N__34333\
        );

    \I__6672\ : InMux
    port map (
            O => \N__34368\,
            I => \N__34330\
        );

    \I__6671\ : InMux
    port map (
            O => \N__34367\,
            I => \N__34317\
        );

    \I__6670\ : InMux
    port map (
            O => \N__34366\,
            I => \N__34317\
        );

    \I__6669\ : InMux
    port map (
            O => \N__34365\,
            I => \N__34317\
        );

    \I__6668\ : InMux
    port map (
            O => \N__34364\,
            I => \N__34317\
        );

    \I__6667\ : InMux
    port map (
            O => \N__34363\,
            I => \N__34317\
        );

    \I__6666\ : InMux
    port map (
            O => \N__34362\,
            I => \N__34317\
        );

    \I__6665\ : InMux
    port map (
            O => \N__34361\,
            I => \N__34314\
        );

    \I__6664\ : InMux
    port map (
            O => \N__34360\,
            I => \N__34311\
        );

    \I__6663\ : InMux
    port map (
            O => \N__34357\,
            I => \N__34308\
        );

    \I__6662\ : CascadeMux
    port map (
            O => \N__34356\,
            I => \N__34296\
        );

    \I__6661\ : InMux
    port map (
            O => \N__34355\,
            I => \N__34286\
        );

    \I__6660\ : Span4Mux_v
    port map (
            O => \N__34350\,
            I => \N__34281\
        );

    \I__6659\ : LocalMux
    port map (
            O => \N__34347\,
            I => \N__34281\
        );

    \I__6658\ : LocalMux
    port map (
            O => \N__34336\,
            I => \N__34276\
        );

    \I__6657\ : LocalMux
    port map (
            O => \N__34333\,
            I => \N__34276\
        );

    \I__6656\ : LocalMux
    port map (
            O => \N__34330\,
            I => \N__34273\
        );

    \I__6655\ : LocalMux
    port map (
            O => \N__34317\,
            I => \N__34268\
        );

    \I__6654\ : LocalMux
    port map (
            O => \N__34314\,
            I => \N__34268\
        );

    \I__6653\ : LocalMux
    port map (
            O => \N__34311\,
            I => \N__34263\
        );

    \I__6652\ : LocalMux
    port map (
            O => \N__34308\,
            I => \N__34263\
        );

    \I__6651\ : InMux
    port map (
            O => \N__34307\,
            I => \N__34252\
        );

    \I__6650\ : InMux
    port map (
            O => \N__34306\,
            I => \N__34239\
        );

    \I__6649\ : InMux
    port map (
            O => \N__34305\,
            I => \N__34239\
        );

    \I__6648\ : InMux
    port map (
            O => \N__34304\,
            I => \N__34239\
        );

    \I__6647\ : InMux
    port map (
            O => \N__34303\,
            I => \N__34239\
        );

    \I__6646\ : InMux
    port map (
            O => \N__34302\,
            I => \N__34239\
        );

    \I__6645\ : InMux
    port map (
            O => \N__34301\,
            I => \N__34239\
        );

    \I__6644\ : InMux
    port map (
            O => \N__34300\,
            I => \N__34236\
        );

    \I__6643\ : InMux
    port map (
            O => \N__34299\,
            I => \N__34233\
        );

    \I__6642\ : InMux
    port map (
            O => \N__34296\,
            I => \N__34224\
        );

    \I__6641\ : InMux
    port map (
            O => \N__34295\,
            I => \N__34224\
        );

    \I__6640\ : InMux
    port map (
            O => \N__34294\,
            I => \N__34224\
        );

    \I__6639\ : InMux
    port map (
            O => \N__34293\,
            I => \N__34224\
        );

    \I__6638\ : InMux
    port map (
            O => \N__34292\,
            I => \N__34215\
        );

    \I__6637\ : InMux
    port map (
            O => \N__34291\,
            I => \N__34215\
        );

    \I__6636\ : InMux
    port map (
            O => \N__34290\,
            I => \N__34215\
        );

    \I__6635\ : InMux
    port map (
            O => \N__34289\,
            I => \N__34215\
        );

    \I__6634\ : LocalMux
    port map (
            O => \N__34286\,
            I => \N__34210\
        );

    \I__6633\ : Span4Mux_h
    port map (
            O => \N__34281\,
            I => \N__34210\
        );

    \I__6632\ : Span4Mux_v
    port map (
            O => \N__34276\,
            I => \N__34201\
        );

    \I__6631\ : Span4Mux_v
    port map (
            O => \N__34273\,
            I => \N__34201\
        );

    \I__6630\ : Span4Mux_v
    port map (
            O => \N__34268\,
            I => \N__34201\
        );

    \I__6629\ : Span4Mux_h
    port map (
            O => \N__34263\,
            I => \N__34201\
        );

    \I__6628\ : InMux
    port map (
            O => \N__34262\,
            I => \N__34184\
        );

    \I__6627\ : InMux
    port map (
            O => \N__34261\,
            I => \N__34184\
        );

    \I__6626\ : InMux
    port map (
            O => \N__34260\,
            I => \N__34184\
        );

    \I__6625\ : InMux
    port map (
            O => \N__34259\,
            I => \N__34184\
        );

    \I__6624\ : InMux
    port map (
            O => \N__34258\,
            I => \N__34184\
        );

    \I__6623\ : InMux
    port map (
            O => \N__34257\,
            I => \N__34184\
        );

    \I__6622\ : InMux
    port map (
            O => \N__34256\,
            I => \N__34184\
        );

    \I__6621\ : InMux
    port map (
            O => \N__34255\,
            I => \N__34184\
        );

    \I__6620\ : LocalMux
    port map (
            O => \N__34252\,
            I => \N__34181\
        );

    \I__6619\ : LocalMux
    port map (
            O => \N__34239\,
            I => adc_state_3
        );

    \I__6618\ : LocalMux
    port map (
            O => \N__34236\,
            I => adc_state_3
        );

    \I__6617\ : LocalMux
    port map (
            O => \N__34233\,
            I => adc_state_3
        );

    \I__6616\ : LocalMux
    port map (
            O => \N__34224\,
            I => adc_state_3
        );

    \I__6615\ : LocalMux
    port map (
            O => \N__34215\,
            I => adc_state_3
        );

    \I__6614\ : Odrv4
    port map (
            O => \N__34210\,
            I => adc_state_3
        );

    \I__6613\ : Odrv4
    port map (
            O => \N__34201\,
            I => adc_state_3
        );

    \I__6612\ : LocalMux
    port map (
            O => \N__34184\,
            I => adc_state_3
        );

    \I__6611\ : Odrv4
    port map (
            O => \N__34181\,
            I => adc_state_3
        );

    \I__6610\ : CascadeMux
    port map (
            O => \N__34162\,
            I => \ADC_VDC.n62_cascade_\
        );

    \I__6609\ : InMux
    port map (
            O => \N__34159\,
            I => \N__34142\
        );

    \I__6608\ : InMux
    port map (
            O => \N__34158\,
            I => \N__34142\
        );

    \I__6607\ : InMux
    port map (
            O => \N__34157\,
            I => \N__34136\
        );

    \I__6606\ : InMux
    port map (
            O => \N__34156\,
            I => \N__34136\
        );

    \I__6605\ : InMux
    port map (
            O => \N__34155\,
            I => \N__34133\
        );

    \I__6604\ : InMux
    port map (
            O => \N__34154\,
            I => \N__34128\
        );

    \I__6603\ : InMux
    port map (
            O => \N__34153\,
            I => \N__34128\
        );

    \I__6602\ : InMux
    port map (
            O => \N__34152\,
            I => \N__34123\
        );

    \I__6601\ : InMux
    port map (
            O => \N__34151\,
            I => \N__34123\
        );

    \I__6600\ : InMux
    port map (
            O => \N__34150\,
            I => \N__34115\
        );

    \I__6599\ : InMux
    port map (
            O => \N__34149\,
            I => \N__34115\
        );

    \I__6598\ : CascadeMux
    port map (
            O => \N__34148\,
            I => \N__34109\
        );

    \I__6597\ : CascadeMux
    port map (
            O => \N__34147\,
            I => \N__34106\
        );

    \I__6596\ : LocalMux
    port map (
            O => \N__34142\,
            I => \N__34103\
        );

    \I__6595\ : InMux
    port map (
            O => \N__34141\,
            I => \N__34100\
        );

    \I__6594\ : LocalMux
    port map (
            O => \N__34136\,
            I => \N__34097\
        );

    \I__6593\ : LocalMux
    port map (
            O => \N__34133\,
            I => \N__34089\
        );

    \I__6592\ : LocalMux
    port map (
            O => \N__34128\,
            I => \N__34089\
        );

    \I__6591\ : LocalMux
    port map (
            O => \N__34123\,
            I => \N__34086\
        );

    \I__6590\ : InMux
    port map (
            O => \N__34122\,
            I => \N__34083\
        );

    \I__6589\ : InMux
    port map (
            O => \N__34121\,
            I => \N__34080\
        );

    \I__6588\ : InMux
    port map (
            O => \N__34120\,
            I => \N__34077\
        );

    \I__6587\ : LocalMux
    port map (
            O => \N__34115\,
            I => \N__34074\
        );

    \I__6586\ : InMux
    port map (
            O => \N__34114\,
            I => \N__34071\
        );

    \I__6585\ : InMux
    port map (
            O => \N__34113\,
            I => \N__34066\
        );

    \I__6584\ : InMux
    port map (
            O => \N__34112\,
            I => \N__34066\
        );

    \I__6583\ : InMux
    port map (
            O => \N__34109\,
            I => \N__34063\
        );

    \I__6582\ : InMux
    port map (
            O => \N__34106\,
            I => \N__34060\
        );

    \I__6581\ : Span4Mux_v
    port map (
            O => \N__34103\,
            I => \N__34057\
        );

    \I__6580\ : LocalMux
    port map (
            O => \N__34100\,
            I => \N__34052\
        );

    \I__6579\ : Span4Mux_h
    port map (
            O => \N__34097\,
            I => \N__34052\
        );

    \I__6578\ : InMux
    port map (
            O => \N__34096\,
            I => \N__34045\
        );

    \I__6577\ : InMux
    port map (
            O => \N__34095\,
            I => \N__34045\
        );

    \I__6576\ : InMux
    port map (
            O => \N__34094\,
            I => \N__34045\
        );

    \I__6575\ : Span4Mux_v
    port map (
            O => \N__34089\,
            I => \N__34042\
        );

    \I__6574\ : Span4Mux_h
    port map (
            O => \N__34086\,
            I => \N__34037\
        );

    \I__6573\ : LocalMux
    port map (
            O => \N__34083\,
            I => \N__34037\
        );

    \I__6572\ : LocalMux
    port map (
            O => \N__34080\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__6571\ : LocalMux
    port map (
            O => \N__34077\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__6570\ : Odrv12
    port map (
            O => \N__34074\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__6569\ : LocalMux
    port map (
            O => \N__34071\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__6568\ : LocalMux
    port map (
            O => \N__34066\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__6567\ : LocalMux
    port map (
            O => \N__34063\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__6566\ : LocalMux
    port map (
            O => \N__34060\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__6565\ : Odrv4
    port map (
            O => \N__34057\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__6564\ : Odrv4
    port map (
            O => \N__34052\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__6563\ : LocalMux
    port map (
            O => \N__34045\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__6562\ : Odrv4
    port map (
            O => \N__34042\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__6561\ : Odrv4
    port map (
            O => \N__34037\,
            I => \ADC_VDC.adc_state_1\
        );

    \I__6560\ : CEMux
    port map (
            O => \N__34012\,
            I => \N__34009\
        );

    \I__6559\ : LocalMux
    port map (
            O => \N__34009\,
            I => \N__34006\
        );

    \I__6558\ : Odrv4
    port map (
            O => \N__34006\,
            I => \ADC_VDC.n11736\
        );

    \I__6557\ : InMux
    port map (
            O => \N__34003\,
            I => \N__34000\
        );

    \I__6556\ : LocalMux
    port map (
            O => \N__34000\,
            I => \N__33997\
        );

    \I__6555\ : Span4Mux_h
    port map (
            O => \N__33997\,
            I => \N__33994\
        );

    \I__6554\ : Span4Mux_h
    port map (
            O => \N__33994\,
            I => \N__33991\
        );

    \I__6553\ : Odrv4
    port map (
            O => \N__33991\,
            I => comm_buf_3_7
        );

    \I__6552\ : InMux
    port map (
            O => \N__33988\,
            I => \N__33985\
        );

    \I__6551\ : LocalMux
    port map (
            O => \N__33985\,
            I => \N__33982\
        );

    \I__6550\ : Odrv4
    port map (
            O => \N__33982\,
            I => n1
        );

    \I__6549\ : CascadeMux
    port map (
            O => \N__33979\,
            I => \n2_adj_1559_cascade_\
        );

    \I__6548\ : InMux
    port map (
            O => \N__33976\,
            I => \N__33973\
        );

    \I__6547\ : LocalMux
    port map (
            O => \N__33973\,
            I => \N__33970\
        );

    \I__6546\ : Span4Mux_h
    port map (
            O => \N__33970\,
            I => \N__33967\
        );

    \I__6545\ : Odrv4
    port map (
            O => \N__33967\,
            I => comm_buf_4_7
        );

    \I__6544\ : InMux
    port map (
            O => \N__33964\,
            I => \N__33961\
        );

    \I__6543\ : LocalMux
    port map (
            O => \N__33961\,
            I => \N__33957\
        );

    \I__6542\ : CascadeMux
    port map (
            O => \N__33960\,
            I => \N__33954\
        );

    \I__6541\ : Span4Mux_h
    port map (
            O => \N__33957\,
            I => \N__33951\
        );

    \I__6540\ : InMux
    port map (
            O => \N__33954\,
            I => \N__33948\
        );

    \I__6539\ : Span4Mux_v
    port map (
            O => \N__33951\,
            I => \N__33945\
        );

    \I__6538\ : LocalMux
    port map (
            O => \N__33948\,
            I => comm_buf_6_7
        );

    \I__6537\ : Odrv4
    port map (
            O => \N__33945\,
            I => comm_buf_6_7
        );

    \I__6536\ : InMux
    port map (
            O => \N__33940\,
            I => n19325
        );

    \I__6535\ : CEMux
    port map (
            O => \N__33937\,
            I => \N__33933\
        );

    \I__6534\ : CEMux
    port map (
            O => \N__33936\,
            I => \N__33930\
        );

    \I__6533\ : LocalMux
    port map (
            O => \N__33933\,
            I => \N__33927\
        );

    \I__6532\ : LocalMux
    port map (
            O => \N__33930\,
            I => \N__33924\
        );

    \I__6531\ : Span4Mux_v
    port map (
            O => \N__33927\,
            I => \N__33918\
        );

    \I__6530\ : Span4Mux_h
    port map (
            O => \N__33924\,
            I => \N__33918\
        );

    \I__6529\ : CEMux
    port map (
            O => \N__33923\,
            I => \N__33915\
        );

    \I__6528\ : Span4Mux_h
    port map (
            O => \N__33918\,
            I => \N__33911\
        );

    \I__6527\ : LocalMux
    port map (
            O => \N__33915\,
            I => \N__33908\
        );

    \I__6526\ : InMux
    port map (
            O => \N__33914\,
            I => \N__33905\
        );

    \I__6525\ : Odrv4
    port map (
            O => \N__33911\,
            I => n11538
        );

    \I__6524\ : Odrv12
    port map (
            O => \N__33908\,
            I => n11538
        );

    \I__6523\ : LocalMux
    port map (
            O => \N__33905\,
            I => n11538
        );

    \I__6522\ : SRMux
    port map (
            O => \N__33898\,
            I => \N__33895\
        );

    \I__6521\ : LocalMux
    port map (
            O => \N__33895\,
            I => \N__33891\
        );

    \I__6520\ : SRMux
    port map (
            O => \N__33894\,
            I => \N__33888\
        );

    \I__6519\ : Span4Mux_h
    port map (
            O => \N__33891\,
            I => \N__33885\
        );

    \I__6518\ : LocalMux
    port map (
            O => \N__33888\,
            I => \N__33882\
        );

    \I__6517\ : Odrv4
    port map (
            O => \N__33885\,
            I => n14639
        );

    \I__6516\ : Odrv4
    port map (
            O => \N__33882\,
            I => n14639
        );

    \I__6515\ : CascadeMux
    port map (
            O => \N__33877\,
            I => \N__33874\
        );

    \I__6514\ : InMux
    port map (
            O => \N__33874\,
            I => \N__33871\
        );

    \I__6513\ : LocalMux
    port map (
            O => \N__33871\,
            I => \SIG_DDS.tmp_buf_11\
        );

    \I__6512\ : InMux
    port map (
            O => \N__33868\,
            I => \N__33865\
        );

    \I__6511\ : LocalMux
    port map (
            O => \N__33865\,
            I => \N__33861\
        );

    \I__6510\ : InMux
    port map (
            O => \N__33864\,
            I => \N__33858\
        );

    \I__6509\ : Span4Mux_h
    port map (
            O => \N__33861\,
            I => \N__33854\
        );

    \I__6508\ : LocalMux
    port map (
            O => \N__33858\,
            I => \N__33851\
        );

    \I__6507\ : InMux
    port map (
            O => \N__33857\,
            I => \N__33848\
        );

    \I__6506\ : Sp12to4
    port map (
            O => \N__33854\,
            I => \N__33843\
        );

    \I__6505\ : Span12Mux_h
    port map (
            O => \N__33851\,
            I => \N__33843\
        );

    \I__6504\ : LocalMux
    port map (
            O => \N__33848\,
            I => buf_dds0_12
        );

    \I__6503\ : Odrv12
    port map (
            O => \N__33843\,
            I => buf_dds0_12
        );

    \I__6502\ : CascadeMux
    port map (
            O => \N__33838\,
            I => \N__33835\
        );

    \I__6501\ : InMux
    port map (
            O => \N__33835\,
            I => \N__33832\
        );

    \I__6500\ : LocalMux
    port map (
            O => \N__33832\,
            I => \SIG_DDS.tmp_buf_12\
        );

    \I__6499\ : CascadeMux
    port map (
            O => \N__33829\,
            I => \N__33826\
        );

    \I__6498\ : InMux
    port map (
            O => \N__33826\,
            I => \N__33823\
        );

    \I__6497\ : LocalMux
    port map (
            O => \N__33823\,
            I => \SIG_DDS.tmp_buf_1\
        );

    \I__6496\ : InMux
    port map (
            O => \N__33820\,
            I => \N__33815\
        );

    \I__6495\ : InMux
    port map (
            O => \N__33819\,
            I => \N__33812\
        );

    \I__6494\ : InMux
    port map (
            O => \N__33818\,
            I => \N__33809\
        );

    \I__6493\ : LocalMux
    port map (
            O => \N__33815\,
            I => \comm_spi.n22632\
        );

    \I__6492\ : LocalMux
    port map (
            O => \N__33812\,
            I => \comm_spi.n22632\
        );

    \I__6491\ : LocalMux
    port map (
            O => \N__33809\,
            I => \comm_spi.n22632\
        );

    \I__6490\ : InMux
    port map (
            O => \N__33802\,
            I => \N__33799\
        );

    \I__6489\ : LocalMux
    port map (
            O => \N__33799\,
            I => \comm_spi.n14600\
        );

    \I__6488\ : SRMux
    port map (
            O => \N__33796\,
            I => \N__33793\
        );

    \I__6487\ : LocalMux
    port map (
            O => \N__33793\,
            I => \N__33790\
        );

    \I__6486\ : Sp12to4
    port map (
            O => \N__33790\,
            I => \N__33787\
        );

    \I__6485\ : Odrv12
    port map (
            O => \N__33787\,
            I => \comm_spi.DOUT_7__N_739\
        );

    \I__6484\ : CascadeMux
    port map (
            O => \N__33784\,
            I => \ADC_VDC.genclk.n21172_cascade_\
        );

    \I__6483\ : InMux
    port map (
            O => \N__33781\,
            I => \N__33777\
        );

    \I__6482\ : InMux
    port map (
            O => \N__33780\,
            I => \N__33774\
        );

    \I__6481\ : LocalMux
    port map (
            O => \N__33777\,
            I => \ADC_VDC.genclk.n21166\
        );

    \I__6480\ : LocalMux
    port map (
            O => \N__33774\,
            I => \ADC_VDC.genclk.n21166\
        );

    \I__6479\ : InMux
    port map (
            O => \N__33769\,
            I => \N__33766\
        );

    \I__6478\ : LocalMux
    port map (
            O => \N__33766\,
            I => \N__33763\
        );

    \I__6477\ : Odrv4
    port map (
            O => \N__33763\,
            I => \ADC_VDC.genclk.n28_adj_1400\
        );

    \I__6476\ : InMux
    port map (
            O => \N__33760\,
            I => \N__33757\
        );

    \I__6475\ : LocalMux
    port map (
            O => \N__33757\,
            I => \ADC_VDC.genclk.n26_adj_1401\
        );

    \I__6474\ : CascadeMux
    port map (
            O => \N__33754\,
            I => \N__33750\
        );

    \I__6473\ : InMux
    port map (
            O => \N__33753\,
            I => \N__33747\
        );

    \I__6472\ : InMux
    port map (
            O => \N__33750\,
            I => \N__33744\
        );

    \I__6471\ : LocalMux
    port map (
            O => \N__33747\,
            I => acadc_skipcnt_6
        );

    \I__6470\ : LocalMux
    port map (
            O => \N__33744\,
            I => acadc_skipcnt_6
        );

    \I__6469\ : InMux
    port map (
            O => \N__33739\,
            I => n19316
        );

    \I__6468\ : InMux
    port map (
            O => \N__33736\,
            I => n19317
        );

    \I__6467\ : InMux
    port map (
            O => \N__33733\,
            I => \N__33730\
        );

    \I__6466\ : LocalMux
    port map (
            O => \N__33730\,
            I => \N__33726\
        );

    \I__6465\ : InMux
    port map (
            O => \N__33729\,
            I => \N__33723\
        );

    \I__6464\ : Span4Mux_h
    port map (
            O => \N__33726\,
            I => \N__33720\
        );

    \I__6463\ : LocalMux
    port map (
            O => \N__33723\,
            I => acadc_skipcnt_8
        );

    \I__6462\ : Odrv4
    port map (
            O => \N__33720\,
            I => acadc_skipcnt_8
        );

    \I__6461\ : InMux
    port map (
            O => \N__33715\,
            I => n19318
        );

    \I__6460\ : InMux
    port map (
            O => \N__33712\,
            I => \bfn_13_18_0_\
        );

    \I__6459\ : InMux
    port map (
            O => \N__33709\,
            I => n19320
        );

    \I__6458\ : InMux
    port map (
            O => \N__33706\,
            I => n19321
        );

    \I__6457\ : InMux
    port map (
            O => \N__33703\,
            I => n19322
        );

    \I__6456\ : InMux
    port map (
            O => \N__33700\,
            I => \N__33697\
        );

    \I__6455\ : LocalMux
    port map (
            O => \N__33697\,
            I => \N__33693\
        );

    \I__6454\ : InMux
    port map (
            O => \N__33696\,
            I => \N__33690\
        );

    \I__6453\ : Span4Mux_h
    port map (
            O => \N__33693\,
            I => \N__33687\
        );

    \I__6452\ : LocalMux
    port map (
            O => \N__33690\,
            I => acadc_skipcnt_13
        );

    \I__6451\ : Odrv4
    port map (
            O => \N__33687\,
            I => acadc_skipcnt_13
        );

    \I__6450\ : InMux
    port map (
            O => \N__33682\,
            I => n19323
        );

    \I__6449\ : InMux
    port map (
            O => \N__33679\,
            I => n19324
        );

    \I__6448\ : InMux
    port map (
            O => \N__33676\,
            I => \N__33672\
        );

    \I__6447\ : InMux
    port map (
            O => \N__33675\,
            I => \N__33669\
        );

    \I__6446\ : LocalMux
    port map (
            O => \N__33672\,
            I => \N__33666\
        );

    \I__6445\ : LocalMux
    port map (
            O => \N__33669\,
            I => acadc_skipcnt_1
        );

    \I__6444\ : Odrv4
    port map (
            O => \N__33666\,
            I => acadc_skipcnt_1
        );

    \I__6443\ : InMux
    port map (
            O => \N__33661\,
            I => \bfn_13_17_0_\
        );

    \I__6442\ : InMux
    port map (
            O => \N__33658\,
            I => n19312
        );

    \I__6441\ : InMux
    port map (
            O => \N__33655\,
            I => \N__33651\
        );

    \I__6440\ : InMux
    port map (
            O => \N__33654\,
            I => \N__33648\
        );

    \I__6439\ : LocalMux
    port map (
            O => \N__33651\,
            I => \N__33645\
        );

    \I__6438\ : LocalMux
    port map (
            O => \N__33648\,
            I => \N__33640\
        );

    \I__6437\ : Span4Mux_v
    port map (
            O => \N__33645\,
            I => \N__33640\
        );

    \I__6436\ : Odrv4
    port map (
            O => \N__33640\,
            I => acadc_skipcnt_3
        );

    \I__6435\ : InMux
    port map (
            O => \N__33637\,
            I => n19313
        );

    \I__6434\ : CascadeMux
    port map (
            O => \N__33634\,
            I => \N__33631\
        );

    \I__6433\ : InMux
    port map (
            O => \N__33631\,
            I => \N__33627\
        );

    \I__6432\ : InMux
    port map (
            O => \N__33630\,
            I => \N__33624\
        );

    \I__6431\ : LocalMux
    port map (
            O => \N__33627\,
            I => \N__33621\
        );

    \I__6430\ : LocalMux
    port map (
            O => \N__33624\,
            I => \N__33616\
        );

    \I__6429\ : Span4Mux_h
    port map (
            O => \N__33621\,
            I => \N__33616\
        );

    \I__6428\ : Odrv4
    port map (
            O => \N__33616\,
            I => acadc_skipcnt_4
        );

    \I__6427\ : InMux
    port map (
            O => \N__33613\,
            I => n19314
        );

    \I__6426\ : InMux
    port map (
            O => \N__33610\,
            I => \N__33607\
        );

    \I__6425\ : LocalMux
    port map (
            O => \N__33607\,
            I => \N__33603\
        );

    \I__6424\ : InMux
    port map (
            O => \N__33606\,
            I => \N__33600\
        );

    \I__6423\ : Span4Mux_h
    port map (
            O => \N__33603\,
            I => \N__33597\
        );

    \I__6422\ : LocalMux
    port map (
            O => \N__33600\,
            I => acadc_skipcnt_5
        );

    \I__6421\ : Odrv4
    port map (
            O => \N__33597\,
            I => acadc_skipcnt_5
        );

    \I__6420\ : InMux
    port map (
            O => \N__33592\,
            I => n19315
        );

    \I__6419\ : CascadeMux
    port map (
            O => \N__33589\,
            I => \n22198_cascade_\
        );

    \I__6418\ : CascadeMux
    port map (
            O => \N__33586\,
            I => \n30_adj_1503_cascade_\
        );

    \I__6417\ : InMux
    port map (
            O => \N__33583\,
            I => \N__33580\
        );

    \I__6416\ : LocalMux
    port map (
            O => \N__33580\,
            I => \N__33577\
        );

    \I__6415\ : Span4Mux_h
    port map (
            O => \N__33577\,
            I => \N__33574\
        );

    \I__6414\ : Odrv4
    port map (
            O => \N__33574\,
            I => n19_adj_1501
        );

    \I__6413\ : CascadeMux
    port map (
            O => \N__33571\,
            I => \N__33568\
        );

    \I__6412\ : InMux
    port map (
            O => \N__33568\,
            I => \N__33565\
        );

    \I__6411\ : LocalMux
    port map (
            O => \N__33565\,
            I => \N__33562\
        );

    \I__6410\ : Span4Mux_h
    port map (
            O => \N__33562\,
            I => \N__33559\
        );

    \I__6409\ : Sp12to4
    port map (
            O => \N__33559\,
            I => \N__33555\
        );

    \I__6408\ : CascadeMux
    port map (
            O => \N__33558\,
            I => \N__33552\
        );

    \I__6407\ : Span12Mux_v
    port map (
            O => \N__33555\,
            I => \N__33549\
        );

    \I__6406\ : InMux
    port map (
            O => \N__33552\,
            I => \N__33546\
        );

    \I__6405\ : Odrv12
    port map (
            O => \N__33549\,
            I => \buf_readRTD_3\
        );

    \I__6404\ : LocalMux
    port map (
            O => \N__33546\,
            I => \buf_readRTD_3\
        );

    \I__6403\ : InMux
    port map (
            O => \N__33541\,
            I => \N__33538\
        );

    \I__6402\ : LocalMux
    port map (
            O => \N__33538\,
            I => \N__33535\
        );

    \I__6401\ : Span4Mux_h
    port map (
            O => \N__33535\,
            I => \N__33530\
        );

    \I__6400\ : InMux
    port map (
            O => \N__33534\,
            I => \N__33527\
        );

    \I__6399\ : InMux
    port map (
            O => \N__33533\,
            I => \N__33524\
        );

    \I__6398\ : Span4Mux_h
    port map (
            O => \N__33530\,
            I => \N__33521\
        );

    \I__6397\ : LocalMux
    port map (
            O => \N__33527\,
            I => buf_adcdata_iac_11
        );

    \I__6396\ : LocalMux
    port map (
            O => \N__33524\,
            I => buf_adcdata_iac_11
        );

    \I__6395\ : Odrv4
    port map (
            O => \N__33521\,
            I => buf_adcdata_iac_11
        );

    \I__6394\ : CascadeMux
    port map (
            O => \N__33514\,
            I => \n22009_cascade_\
        );

    \I__6393\ : InMux
    port map (
            O => \N__33511\,
            I => \N__33508\
        );

    \I__6392\ : LocalMux
    port map (
            O => \N__33508\,
            I => \N__33505\
        );

    \I__6391\ : Odrv12
    port map (
            O => \N__33505\,
            I => n16_adj_1500
        );

    \I__6390\ : InMux
    port map (
            O => \N__33502\,
            I => \N__33499\
        );

    \I__6389\ : LocalMux
    port map (
            O => \N__33499\,
            I => n22012
        );

    \I__6388\ : CascadeMux
    port map (
            O => \N__33496\,
            I => \N__33493\
        );

    \I__6387\ : InMux
    port map (
            O => \N__33493\,
            I => \N__33489\
        );

    \I__6386\ : InMux
    port map (
            O => \N__33492\,
            I => \N__33486\
        );

    \I__6385\ : LocalMux
    port map (
            O => \N__33489\,
            I => acadc_skipcnt_0
        );

    \I__6384\ : LocalMux
    port map (
            O => \N__33486\,
            I => acadc_skipcnt_0
        );

    \I__6383\ : SRMux
    port map (
            O => \N__33481\,
            I => \N__33478\
        );

    \I__6382\ : LocalMux
    port map (
            O => \N__33478\,
            I => \N__33475\
        );

    \I__6381\ : Span4Mux_h
    port map (
            O => \N__33475\,
            I => \N__33472\
        );

    \I__6380\ : Odrv4
    port map (
            O => \N__33472\,
            I => n20757
        );

    \I__6379\ : InMux
    port map (
            O => \N__33469\,
            I => \N__33466\
        );

    \I__6378\ : LocalMux
    port map (
            O => \N__33466\,
            I => \N__33463\
        );

    \I__6377\ : Span4Mux_v
    port map (
            O => \N__33463\,
            I => \N__33458\
        );

    \I__6376\ : InMux
    port map (
            O => \N__33462\,
            I => \N__33455\
        );

    \I__6375\ : InMux
    port map (
            O => \N__33461\,
            I => \N__33452\
        );

    \I__6374\ : Span4Mux_h
    port map (
            O => \N__33458\,
            I => \N__33449\
        );

    \I__6373\ : LocalMux
    port map (
            O => \N__33455\,
            I => buf_adcdata_iac_12
        );

    \I__6372\ : LocalMux
    port map (
            O => \N__33452\,
            I => buf_adcdata_iac_12
        );

    \I__6371\ : Odrv4
    port map (
            O => \N__33449\,
            I => buf_adcdata_iac_12
        );

    \I__6370\ : CascadeMux
    port map (
            O => \N__33442\,
            I => \n22081_cascade_\
        );

    \I__6369\ : CascadeMux
    port map (
            O => \N__33439\,
            I => \N__33435\
        );

    \I__6368\ : InMux
    port map (
            O => \N__33438\,
            I => \N__33432\
        );

    \I__6367\ : InMux
    port map (
            O => \N__33435\,
            I => \N__33429\
        );

    \I__6366\ : LocalMux
    port map (
            O => \N__33432\,
            I => \N__33426\
        );

    \I__6365\ : LocalMux
    port map (
            O => \N__33429\,
            I => data_idxvec_4
        );

    \I__6364\ : Odrv4
    port map (
            O => \N__33426\,
            I => data_idxvec_4
        );

    \I__6363\ : InMux
    port map (
            O => \N__33421\,
            I => \N__33418\
        );

    \I__6362\ : LocalMux
    port map (
            O => \N__33418\,
            I => \N__33415\
        );

    \I__6361\ : Span4Mux_h
    port map (
            O => \N__33415\,
            I => \N__33412\
        );

    \I__6360\ : Odrv4
    port map (
            O => \N__33412\,
            I => n21261
        );

    \I__6359\ : CascadeMux
    port map (
            O => \N__33409\,
            I => \n26_adj_1484_cascade_\
        );

    \I__6358\ : CascadeMux
    port map (
            O => \N__33406\,
            I => \n22159_cascade_\
        );

    \I__6357\ : InMux
    port map (
            O => \N__33403\,
            I => \N__33400\
        );

    \I__6356\ : LocalMux
    port map (
            O => \N__33400\,
            I => n22084
        );

    \I__6355\ : CascadeMux
    port map (
            O => \N__33397\,
            I => \n22162_cascade_\
        );

    \I__6354\ : CascadeMux
    port map (
            O => \N__33394\,
            I => \n30_adj_1493_cascade_\
        );

    \I__6353\ : InMux
    port map (
            O => \N__33391\,
            I => \N__33387\
        );

    \I__6352\ : InMux
    port map (
            O => \N__33390\,
            I => \N__33384\
        );

    \I__6351\ : LocalMux
    port map (
            O => \N__33387\,
            I => \N__33381\
        );

    \I__6350\ : LocalMux
    port map (
            O => \N__33384\,
            I => data_idxvec_3
        );

    \I__6349\ : Odrv4
    port map (
            O => \N__33381\,
            I => data_idxvec_3
        );

    \I__6348\ : InMux
    port map (
            O => \N__33376\,
            I => \N__33373\
        );

    \I__6347\ : LocalMux
    port map (
            O => \N__33373\,
            I => \N__33370\
        );

    \I__6346\ : Span4Mux_h
    port map (
            O => \N__33370\,
            I => \N__33367\
        );

    \I__6345\ : Span4Mux_h
    port map (
            O => \N__33367\,
            I => \N__33364\
        );

    \I__6344\ : Odrv4
    port map (
            O => \N__33364\,
            I => n21285
        );

    \I__6343\ : CascadeMux
    port map (
            O => \N__33361\,
            I => \n26_adj_1502_cascade_\
        );

    \I__6342\ : CascadeMux
    port map (
            O => \N__33358\,
            I => \n22195_cascade_\
        );

    \I__6341\ : InMux
    port map (
            O => \N__33355\,
            I => \N__33350\
        );

    \I__6340\ : InMux
    port map (
            O => \N__33354\,
            I => \N__33345\
        );

    \I__6339\ : InMux
    port map (
            O => \N__33353\,
            I => \N__33345\
        );

    \I__6338\ : LocalMux
    port map (
            O => \N__33350\,
            I => \acadc_skipCount_3\
        );

    \I__6337\ : LocalMux
    port map (
            O => \N__33345\,
            I => \acadc_skipCount_3\
        );

    \I__6336\ : CascadeMux
    port map (
            O => \N__33340\,
            I => \N__33337\
        );

    \I__6335\ : InMux
    port map (
            O => \N__33337\,
            I => \N__33333\
        );

    \I__6334\ : InMux
    port map (
            O => \N__33336\,
            I => \N__33330\
        );

    \I__6333\ : LocalMux
    port map (
            O => \N__33333\,
            I => data_idxvec_2
        );

    \I__6332\ : LocalMux
    port map (
            O => \N__33330\,
            I => data_idxvec_2
        );

    \I__6331\ : CascadeMux
    port map (
            O => \N__33325\,
            I => \n26_adj_1506_cascade_\
        );

    \I__6330\ : InMux
    port map (
            O => \N__33322\,
            I => \N__33319\
        );

    \I__6329\ : LocalMux
    port map (
            O => \N__33319\,
            I => \N__33316\
        );

    \I__6328\ : Span4Mux_v
    port map (
            O => \N__33316\,
            I => \N__33313\
        );

    \I__6327\ : Span4Mux_h
    port map (
            O => \N__33313\,
            I => \N__33310\
        );

    \I__6326\ : Span4Mux_h
    port map (
            O => \N__33310\,
            I => \N__33307\
        );

    \I__6325\ : Odrv4
    port map (
            O => \N__33307\,
            I => buf_data_iac_10
        );

    \I__6324\ : CascadeMux
    port map (
            O => \N__33304\,
            I => \n20816_cascade_\
        );

    \I__6323\ : InMux
    port map (
            O => \N__33301\,
            I => \N__33298\
        );

    \I__6322\ : LocalMux
    port map (
            O => \N__33298\,
            I => \N__33295\
        );

    \I__6321\ : Span4Mux_v
    port map (
            O => \N__33295\,
            I => \N__33292\
        );

    \I__6320\ : Span4Mux_h
    port map (
            O => \N__33292\,
            I => \N__33289\
        );

    \I__6319\ : Odrv4
    port map (
            O => \N__33289\,
            I => n20845
        );

    \I__6318\ : CascadeMux
    port map (
            O => \N__33286\,
            I => \n22087_cascade_\
        );

    \I__6317\ : CascadeMux
    port map (
            O => \N__33283\,
            I => \n22090_cascade_\
        );

    \I__6316\ : InMux
    port map (
            O => \N__33280\,
            I => \N__33277\
        );

    \I__6315\ : LocalMux
    port map (
            O => \N__33277\,
            I => \N__33274\
        );

    \I__6314\ : Odrv12
    port map (
            O => \N__33274\,
            I => n19_adj_1505
        );

    \I__6313\ : InMux
    port map (
            O => \N__33271\,
            I => \N__33268\
        );

    \I__6312\ : LocalMux
    port map (
            O => \N__33268\,
            I => \N__33265\
        );

    \I__6311\ : Span4Mux_v
    port map (
            O => \N__33265\,
            I => \N__33262\
        );

    \I__6310\ : Span4Mux_h
    port map (
            O => \N__33262\,
            I => \N__33258\
        );

    \I__6309\ : CascadeMux
    port map (
            O => \N__33261\,
            I => \N__33255\
        );

    \I__6308\ : Span4Mux_h
    port map (
            O => \N__33258\,
            I => \N__33252\
        );

    \I__6307\ : InMux
    port map (
            O => \N__33255\,
            I => \N__33249\
        );

    \I__6306\ : Odrv4
    port map (
            O => \N__33252\,
            I => \buf_readRTD_2\
        );

    \I__6305\ : LocalMux
    port map (
            O => \N__33249\,
            I => \buf_readRTD_2\
        );

    \I__6304\ : InMux
    port map (
            O => \N__33244\,
            I => \N__33241\
        );

    \I__6303\ : LocalMux
    port map (
            O => \N__33241\,
            I => n20846
        );

    \I__6302\ : InMux
    port map (
            O => \N__33238\,
            I => \N__33235\
        );

    \I__6301\ : LocalMux
    port map (
            O => \N__33235\,
            I => n20815
        );

    \I__6300\ : InMux
    port map (
            O => \N__33232\,
            I => \N__33229\
        );

    \I__6299\ : LocalMux
    port map (
            O => \N__33229\,
            I => \N__33226\
        );

    \I__6298\ : Span4Mux_v
    port map (
            O => \N__33226\,
            I => \N__33223\
        );

    \I__6297\ : Span4Mux_h
    port map (
            O => \N__33223\,
            I => \N__33220\
        );

    \I__6296\ : Odrv4
    port map (
            O => \N__33220\,
            I => n19
        );

    \I__6295\ : CascadeMux
    port map (
            O => \N__33217\,
            I => \N__33214\
        );

    \I__6294\ : InMux
    port map (
            O => \N__33214\,
            I => \N__33211\
        );

    \I__6293\ : LocalMux
    port map (
            O => \N__33211\,
            I => \N__33208\
        );

    \I__6292\ : Span4Mux_v
    port map (
            O => \N__33208\,
            I => \N__33204\
        );

    \I__6291\ : CascadeMux
    port map (
            O => \N__33207\,
            I => \N__33201\
        );

    \I__6290\ : Sp12to4
    port map (
            O => \N__33204\,
            I => \N__33198\
        );

    \I__6289\ : InMux
    port map (
            O => \N__33201\,
            I => \N__33195\
        );

    \I__6288\ : Odrv12
    port map (
            O => \N__33198\,
            I => \buf_readRTD_4\
        );

    \I__6287\ : LocalMux
    port map (
            O => \N__33195\,
            I => \buf_readRTD_4\
        );

    \I__6286\ : InMux
    port map (
            O => \N__33190\,
            I => \N__33187\
        );

    \I__6285\ : LocalMux
    port map (
            O => \N__33187\,
            I => \N__33184\
        );

    \I__6284\ : Span4Mux_v
    port map (
            O => \N__33184\,
            I => \N__33181\
        );

    \I__6283\ : Span4Mux_h
    port map (
            O => \N__33181\,
            I => \N__33178\
        );

    \I__6282\ : Odrv4
    port map (
            O => \N__33178\,
            I => comm_buf_3_5
        );

    \I__6281\ : CascadeMux
    port map (
            O => \N__33175\,
            I => \n17331_cascade_\
        );

    \I__6280\ : CascadeMux
    port map (
            O => \N__33172\,
            I => \n20903_cascade_\
        );

    \I__6279\ : CascadeMux
    port map (
            O => \N__33169\,
            I => \n1_adj_1561_cascade_\
        );

    \I__6278\ : CascadeMux
    port map (
            O => \N__33166\,
            I => \N__33163\
        );

    \I__6277\ : InMux
    port map (
            O => \N__33163\,
            I => \N__33159\
        );

    \I__6276\ : InMux
    port map (
            O => \N__33162\,
            I => \N__33156\
        );

    \I__6275\ : LocalMux
    port map (
            O => \N__33159\,
            I => \N__33151\
        );

    \I__6274\ : LocalMux
    port map (
            O => \N__33156\,
            I => \N__33151\
        );

    \I__6273\ : Odrv12
    port map (
            O => \N__33151\,
            I => comm_buf_6_6
        );

    \I__6272\ : CascadeMux
    port map (
            O => \N__33148\,
            I => \N__33145\
        );

    \I__6271\ : InMux
    port map (
            O => \N__33145\,
            I => \N__33142\
        );

    \I__6270\ : LocalMux
    port map (
            O => \N__33142\,
            I => \N__33139\
        );

    \I__6269\ : Span4Mux_v
    port map (
            O => \N__33139\,
            I => \N__33136\
        );

    \I__6268\ : Odrv4
    port map (
            O => \N__33136\,
            I => comm_buf_3_6
        );

    \I__6267\ : InMux
    port map (
            O => \N__33133\,
            I => \N__33130\
        );

    \I__6266\ : LocalMux
    port map (
            O => \N__33130\,
            I => n2_adj_1562
        );

    \I__6265\ : InMux
    port map (
            O => \N__33127\,
            I => \N__33124\
        );

    \I__6264\ : LocalMux
    port map (
            O => \N__33124\,
            I => comm_buf_4_6
        );

    \I__6263\ : InMux
    port map (
            O => \N__33121\,
            I => \N__33118\
        );

    \I__6262\ : LocalMux
    port map (
            O => \N__33118\,
            I => n21051
        );

    \I__6261\ : CascadeMux
    port map (
            O => \N__33115\,
            I => \n4_adj_1563_cascade_\
        );

    \I__6260\ : InMux
    port map (
            O => \N__33112\,
            I => \N__33109\
        );

    \I__6259\ : LocalMux
    port map (
            O => \N__33109\,
            I => n22093
        );

    \I__6258\ : SRMux
    port map (
            O => \N__33106\,
            I => \N__33103\
        );

    \I__6257\ : LocalMux
    port map (
            O => \N__33103\,
            I => n14763
        );

    \I__6256\ : CascadeMux
    port map (
            O => \N__33100\,
            I => \N__33097\
        );

    \I__6255\ : InMux
    port map (
            O => \N__33097\,
            I => \N__33094\
        );

    \I__6254\ : LocalMux
    port map (
            O => \N__33094\,
            I => \N__33091\
        );

    \I__6253\ : Span4Mux_h
    port map (
            O => \N__33091\,
            I => \N__33088\
        );

    \I__6252\ : Odrv4
    port map (
            O => \N__33088\,
            I => comm_buf_3_3
        );

    \I__6251\ : CascadeMux
    port map (
            O => \N__33085\,
            I => \n21979_cascade_\
        );

    \I__6250\ : InMux
    port map (
            O => \N__33082\,
            I => \N__33079\
        );

    \I__6249\ : LocalMux
    port map (
            O => \N__33079\,
            I => comm_buf_4_3
        );

    \I__6248\ : InMux
    port map (
            O => \N__33076\,
            I => \N__33072\
        );

    \I__6247\ : InMux
    port map (
            O => \N__33075\,
            I => \N__33069\
        );

    \I__6246\ : LocalMux
    port map (
            O => \N__33072\,
            I => \N__33066\
        );

    \I__6245\ : LocalMux
    port map (
            O => \N__33069\,
            I => comm_buf_6_3
        );

    \I__6244\ : Odrv4
    port map (
            O => \N__33066\,
            I => comm_buf_6_3
        );

    \I__6243\ : CascadeMux
    port map (
            O => \N__33061\,
            I => \n4_adj_1567_cascade_\
        );

    \I__6242\ : CascadeMux
    port map (
            O => \N__33058\,
            I => \n20783_cascade_\
        );

    \I__6241\ : InMux
    port map (
            O => \N__33055\,
            I => \N__33052\
        );

    \I__6240\ : LocalMux
    port map (
            O => \N__33052\,
            I => n21982
        );

    \I__6239\ : SRMux
    port map (
            O => \N__33049\,
            I => \N__33046\
        );

    \I__6238\ : LocalMux
    port map (
            O => \N__33046\,
            I => \N__33043\
        );

    \I__6237\ : Odrv12
    port map (
            O => \N__33043\,
            I => \comm_spi.data_tx_7__N_762\
        );

    \I__6236\ : CEMux
    port map (
            O => \N__33040\,
            I => \N__33037\
        );

    \I__6235\ : LocalMux
    port map (
            O => \N__33037\,
            I => n11727
        );

    \I__6234\ : InMux
    port map (
            O => \N__33034\,
            I => \N__33024\
        );

    \I__6233\ : InMux
    port map (
            O => \N__33033\,
            I => \N__33024\
        );

    \I__6232\ : InMux
    port map (
            O => \N__33032\,
            I => \N__33024\
        );

    \I__6231\ : InMux
    port map (
            O => \N__33031\,
            I => \N__33021\
        );

    \I__6230\ : LocalMux
    port map (
            O => \N__33024\,
            I => \comm_spi.bit_cnt_1\
        );

    \I__6229\ : LocalMux
    port map (
            O => \N__33021\,
            I => \comm_spi.bit_cnt_1\
        );

    \I__6228\ : CascadeMux
    port map (
            O => \N__33016\,
            I => \N__33012\
        );

    \I__6227\ : InMux
    port map (
            O => \N__33015\,
            I => \N__33006\
        );

    \I__6226\ : InMux
    port map (
            O => \N__33012\,
            I => \N__32997\
        );

    \I__6225\ : InMux
    port map (
            O => \N__33011\,
            I => \N__32997\
        );

    \I__6224\ : InMux
    port map (
            O => \N__33010\,
            I => \N__32997\
        );

    \I__6223\ : InMux
    port map (
            O => \N__33009\,
            I => \N__32997\
        );

    \I__6222\ : LocalMux
    port map (
            O => \N__33006\,
            I => \N__32994\
        );

    \I__6221\ : LocalMux
    port map (
            O => \N__32997\,
            I => \comm_spi.bit_cnt_0\
        );

    \I__6220\ : Odrv4
    port map (
            O => \N__32994\,
            I => \comm_spi.bit_cnt_0\
        );

    \I__6219\ : InMux
    port map (
            O => \N__32989\,
            I => \N__32984\
        );

    \I__6218\ : InMux
    port map (
            O => \N__32988\,
            I => \N__32979\
        );

    \I__6217\ : InMux
    port map (
            O => \N__32987\,
            I => \N__32979\
        );

    \I__6216\ : LocalMux
    port map (
            O => \N__32984\,
            I => \N__32976\
        );

    \I__6215\ : LocalMux
    port map (
            O => \N__32979\,
            I => \comm_spi.bit_cnt_2\
        );

    \I__6214\ : Odrv4
    port map (
            O => \N__32976\,
            I => \comm_spi.bit_cnt_2\
        );

    \I__6213\ : CascadeMux
    port map (
            O => \N__32971\,
            I => \N__32968\
        );

    \I__6212\ : InMux
    port map (
            O => \N__32968\,
            I => \N__32965\
        );

    \I__6211\ : LocalMux
    port map (
            O => \N__32965\,
            I => \N__32962\
        );

    \I__6210\ : Span4Mux_h
    port map (
            O => \N__32962\,
            I => \N__32959\
        );

    \I__6209\ : Odrv4
    port map (
            O => \N__32959\,
            I => comm_buf_3_1
        );

    \I__6208\ : CascadeMux
    port map (
            O => \N__32956\,
            I => \n21991_cascade_\
        );

    \I__6207\ : InMux
    port map (
            O => \N__32953\,
            I => \N__32948\
        );

    \I__6206\ : InMux
    port map (
            O => \N__32952\,
            I => \N__32943\
        );

    \I__6205\ : InMux
    port map (
            O => \N__32951\,
            I => \N__32943\
        );

    \I__6204\ : LocalMux
    port map (
            O => \N__32948\,
            I => \ADC_VDC.bit_cnt_6\
        );

    \I__6203\ : LocalMux
    port map (
            O => \N__32943\,
            I => \ADC_VDC.bit_cnt_6\
        );

    \I__6202\ : InMux
    port map (
            O => \N__32938\,
            I => \ADC_VDC.n19474\
        );

    \I__6201\ : InMux
    port map (
            O => \N__32935\,
            I => \ADC_VDC.n19475\
        );

    \I__6200\ : InMux
    port map (
            O => \N__32932\,
            I => \N__32927\
        );

    \I__6199\ : InMux
    port map (
            O => \N__32931\,
            I => \N__32924\
        );

    \I__6198\ : InMux
    port map (
            O => \N__32930\,
            I => \N__32921\
        );

    \I__6197\ : LocalMux
    port map (
            O => \N__32927\,
            I => \ADC_VDC.bit_cnt_7\
        );

    \I__6196\ : LocalMux
    port map (
            O => \N__32924\,
            I => \ADC_VDC.bit_cnt_7\
        );

    \I__6195\ : LocalMux
    port map (
            O => \N__32921\,
            I => \ADC_VDC.bit_cnt_7\
        );

    \I__6194\ : IoInMux
    port map (
            O => \N__32914\,
            I => \N__32909\
        );

    \I__6193\ : ClkMux
    port map (
            O => \N__32913\,
            I => \N__32905\
        );

    \I__6192\ : ClkMux
    port map (
            O => \N__32912\,
            I => \N__32900\
        );

    \I__6191\ : LocalMux
    port map (
            O => \N__32909\,
            I => \N__32897\
        );

    \I__6190\ : ClkMux
    port map (
            O => \N__32908\,
            I => \N__32890\
        );

    \I__6189\ : LocalMux
    port map (
            O => \N__32905\,
            I => \N__32887\
        );

    \I__6188\ : ClkMux
    port map (
            O => \N__32904\,
            I => \N__32881\
        );

    \I__6187\ : ClkMux
    port map (
            O => \N__32903\,
            I => \N__32877\
        );

    \I__6186\ : LocalMux
    port map (
            O => \N__32900\,
            I => \N__32874\
        );

    \I__6185\ : IoSpan4Mux
    port map (
            O => \N__32897\,
            I => \N__32868\
        );

    \I__6184\ : ClkMux
    port map (
            O => \N__32896\,
            I => \N__32865\
        );

    \I__6183\ : ClkMux
    port map (
            O => \N__32895\,
            I => \N__32862\
        );

    \I__6182\ : ClkMux
    port map (
            O => \N__32894\,
            I => \N__32858\
        );

    \I__6181\ : ClkMux
    port map (
            O => \N__32893\,
            I => \N__32855\
        );

    \I__6180\ : LocalMux
    port map (
            O => \N__32890\,
            I => \N__32850\
        );

    \I__6179\ : Span4Mux_h
    port map (
            O => \N__32887\,
            I => \N__32850\
        );

    \I__6178\ : ClkMux
    port map (
            O => \N__32886\,
            I => \N__32847\
        );

    \I__6177\ : ClkMux
    port map (
            O => \N__32885\,
            I => \N__32843\
        );

    \I__6176\ : ClkMux
    port map (
            O => \N__32884\,
            I => \N__32839\
        );

    \I__6175\ : LocalMux
    port map (
            O => \N__32881\,
            I => \N__32836\
        );

    \I__6174\ : ClkMux
    port map (
            O => \N__32880\,
            I => \N__32833\
        );

    \I__6173\ : LocalMux
    port map (
            O => \N__32877\,
            I => \N__32830\
        );

    \I__6172\ : Span4Mux_h
    port map (
            O => \N__32874\,
            I => \N__32827\
        );

    \I__6171\ : ClkMux
    port map (
            O => \N__32873\,
            I => \N__32824\
        );

    \I__6170\ : ClkMux
    port map (
            O => \N__32872\,
            I => \N__32821\
        );

    \I__6169\ : ClkMux
    port map (
            O => \N__32871\,
            I => \N__32818\
        );

    \I__6168\ : Span4Mux_s3_h
    port map (
            O => \N__32868\,
            I => \N__32815\
        );

    \I__6167\ : LocalMux
    port map (
            O => \N__32865\,
            I => \N__32810\
        );

    \I__6166\ : LocalMux
    port map (
            O => \N__32862\,
            I => \N__32810\
        );

    \I__6165\ : ClkMux
    port map (
            O => \N__32861\,
            I => \N__32807\
        );

    \I__6164\ : LocalMux
    port map (
            O => \N__32858\,
            I => \N__32801\
        );

    \I__6163\ : LocalMux
    port map (
            O => \N__32855\,
            I => \N__32801\
        );

    \I__6162\ : Span4Mux_h
    port map (
            O => \N__32850\,
            I => \N__32796\
        );

    \I__6161\ : LocalMux
    port map (
            O => \N__32847\,
            I => \N__32796\
        );

    \I__6160\ : ClkMux
    port map (
            O => \N__32846\,
            I => \N__32793\
        );

    \I__6159\ : LocalMux
    port map (
            O => \N__32843\,
            I => \N__32790\
        );

    \I__6158\ : ClkMux
    port map (
            O => \N__32842\,
            I => \N__32787\
        );

    \I__6157\ : LocalMux
    port map (
            O => \N__32839\,
            I => \N__32784\
        );

    \I__6156\ : Span4Mux_h
    port map (
            O => \N__32836\,
            I => \N__32779\
        );

    \I__6155\ : LocalMux
    port map (
            O => \N__32833\,
            I => \N__32779\
        );

    \I__6154\ : Span4Mux_h
    port map (
            O => \N__32830\,
            I => \N__32775\
        );

    \I__6153\ : Span4Mux_v
    port map (
            O => \N__32827\,
            I => \N__32770\
        );

    \I__6152\ : LocalMux
    port map (
            O => \N__32824\,
            I => \N__32770\
        );

    \I__6151\ : LocalMux
    port map (
            O => \N__32821\,
            I => \N__32765\
        );

    \I__6150\ : LocalMux
    port map (
            O => \N__32818\,
            I => \N__32765\
        );

    \I__6149\ : Span4Mux_h
    port map (
            O => \N__32815\,
            I => \N__32762\
        );

    \I__6148\ : Span4Mux_h
    port map (
            O => \N__32810\,
            I => \N__32757\
        );

    \I__6147\ : LocalMux
    port map (
            O => \N__32807\,
            I => \N__32757\
        );

    \I__6146\ : ClkMux
    port map (
            O => \N__32806\,
            I => \N__32754\
        );

    \I__6145\ : Span4Mux_h
    port map (
            O => \N__32801\,
            I => \N__32751\
        );

    \I__6144\ : Span4Mux_v
    port map (
            O => \N__32796\,
            I => \N__32746\
        );

    \I__6143\ : LocalMux
    port map (
            O => \N__32793\,
            I => \N__32746\
        );

    \I__6142\ : Span4Mux_v
    port map (
            O => \N__32790\,
            I => \N__32741\
        );

    \I__6141\ : LocalMux
    port map (
            O => \N__32787\,
            I => \N__32741\
        );

    \I__6140\ : Span4Mux_h
    port map (
            O => \N__32784\,
            I => \N__32736\
        );

    \I__6139\ : Span4Mux_h
    port map (
            O => \N__32779\,
            I => \N__32736\
        );

    \I__6138\ : ClkMux
    port map (
            O => \N__32778\,
            I => \N__32733\
        );

    \I__6137\ : Span4Mux_v
    port map (
            O => \N__32775\,
            I => \N__32728\
        );

    \I__6136\ : Span4Mux_h
    port map (
            O => \N__32770\,
            I => \N__32728\
        );

    \I__6135\ : Span4Mux_h
    port map (
            O => \N__32765\,
            I => \N__32724\
        );

    \I__6134\ : Span4Mux_h
    port map (
            O => \N__32762\,
            I => \N__32719\
        );

    \I__6133\ : Span4Mux_v
    port map (
            O => \N__32757\,
            I => \N__32719\
        );

    \I__6132\ : LocalMux
    port map (
            O => \N__32754\,
            I => \N__32716\
        );

    \I__6131\ : Span4Mux_v
    port map (
            O => \N__32751\,
            I => \N__32711\
        );

    \I__6130\ : Span4Mux_h
    port map (
            O => \N__32746\,
            I => \N__32711\
        );

    \I__6129\ : Span4Mux_h
    port map (
            O => \N__32741\,
            I => \N__32704\
        );

    \I__6128\ : Span4Mux_v
    port map (
            O => \N__32736\,
            I => \N__32704\
        );

    \I__6127\ : LocalMux
    port map (
            O => \N__32733\,
            I => \N__32704\
        );

    \I__6126\ : Span4Mux_v
    port map (
            O => \N__32728\,
            I => \N__32701\
        );

    \I__6125\ : ClkMux
    port map (
            O => \N__32727\,
            I => \N__32698\
        );

    \I__6124\ : Span4Mux_v
    port map (
            O => \N__32724\,
            I => \N__32693\
        );

    \I__6123\ : Span4Mux_h
    port map (
            O => \N__32719\,
            I => \N__32693\
        );

    \I__6122\ : Span4Mux_h
    port map (
            O => \N__32716\,
            I => \N__32688\
        );

    \I__6121\ : Span4Mux_v
    port map (
            O => \N__32711\,
            I => \N__32688\
        );

    \I__6120\ : Sp12to4
    port map (
            O => \N__32704\,
            I => \N__32685\
        );

    \I__6119\ : Span4Mux_h
    port map (
            O => \N__32701\,
            I => \N__32680\
        );

    \I__6118\ : LocalMux
    port map (
            O => \N__32698\,
            I => \N__32680\
        );

    \I__6117\ : Odrv4
    port map (
            O => \N__32693\,
            I => \VDC_CLK\
        );

    \I__6116\ : Odrv4
    port map (
            O => \N__32688\,
            I => \VDC_CLK\
        );

    \I__6115\ : Odrv12
    port map (
            O => \N__32685\,
            I => \VDC_CLK\
        );

    \I__6114\ : Odrv4
    port map (
            O => \N__32680\,
            I => \VDC_CLK\
        );

    \I__6113\ : SRMux
    port map (
            O => \N__32671\,
            I => \N__32668\
        );

    \I__6112\ : LocalMux
    port map (
            O => \N__32668\,
            I => \N__32665\
        );

    \I__6111\ : Span4Mux_h
    port map (
            O => \N__32665\,
            I => \N__32662\
        );

    \I__6110\ : Odrv4
    port map (
            O => \N__32662\,
            I => \ADC_VDC.n18381\
        );

    \I__6109\ : InMux
    port map (
            O => \N__32659\,
            I => \N__32656\
        );

    \I__6108\ : LocalMux
    port map (
            O => \N__32656\,
            I => \N__32653\
        );

    \I__6107\ : Span4Mux_v
    port map (
            O => \N__32653\,
            I => \N__32650\
        );

    \I__6106\ : Span4Mux_h
    port map (
            O => \N__32650\,
            I => \N__32647\
        );

    \I__6105\ : Span4Mux_h
    port map (
            O => \N__32647\,
            I => \N__32644\
        );

    \I__6104\ : Odrv4
    port map (
            O => \N__32644\,
            I => buf_data_iac_6
        );

    \I__6103\ : InMux
    port map (
            O => \N__32641\,
            I => \N__32637\
        );

    \I__6102\ : CascadeMux
    port map (
            O => \N__32640\,
            I => \N__32634\
        );

    \I__6101\ : LocalMux
    port map (
            O => \N__32637\,
            I => \N__32629\
        );

    \I__6100\ : InMux
    port map (
            O => \N__32634\,
            I => \N__32626\
        );

    \I__6099\ : InMux
    port map (
            O => \N__32633\,
            I => \N__32622\
        );

    \I__6098\ : InMux
    port map (
            O => \N__32632\,
            I => \N__32619\
        );

    \I__6097\ : Span4Mux_v
    port map (
            O => \N__32629\,
            I => \N__32616\
        );

    \I__6096\ : LocalMux
    port map (
            O => \N__32626\,
            I => \N__32613\
        );

    \I__6095\ : InMux
    port map (
            O => \N__32625\,
            I => \N__32610\
        );

    \I__6094\ : LocalMux
    port map (
            O => \N__32622\,
            I => \ADC_VDC.bit_cnt_3\
        );

    \I__6093\ : LocalMux
    port map (
            O => \N__32619\,
            I => \ADC_VDC.bit_cnt_3\
        );

    \I__6092\ : Odrv4
    port map (
            O => \N__32616\,
            I => \ADC_VDC.bit_cnt_3\
        );

    \I__6091\ : Odrv4
    port map (
            O => \N__32613\,
            I => \ADC_VDC.bit_cnt_3\
        );

    \I__6090\ : LocalMux
    port map (
            O => \N__32610\,
            I => \ADC_VDC.bit_cnt_3\
        );

    \I__6089\ : InMux
    port map (
            O => \N__32599\,
            I => \N__32596\
        );

    \I__6088\ : LocalMux
    port map (
            O => \N__32596\,
            I => \N__32592\
        );

    \I__6087\ : InMux
    port map (
            O => \N__32595\,
            I => \N__32586\
        );

    \I__6086\ : Span4Mux_v
    port map (
            O => \N__32592\,
            I => \N__32583\
        );

    \I__6085\ : InMux
    port map (
            O => \N__32591\,
            I => \N__32580\
        );

    \I__6084\ : InMux
    port map (
            O => \N__32590\,
            I => \N__32575\
        );

    \I__6083\ : InMux
    port map (
            O => \N__32589\,
            I => \N__32575\
        );

    \I__6082\ : LocalMux
    port map (
            O => \N__32586\,
            I => \ADC_VDC.bit_cnt_2\
        );

    \I__6081\ : Odrv4
    port map (
            O => \N__32583\,
            I => \ADC_VDC.bit_cnt_2\
        );

    \I__6080\ : LocalMux
    port map (
            O => \N__32580\,
            I => \ADC_VDC.bit_cnt_2\
        );

    \I__6079\ : LocalMux
    port map (
            O => \N__32575\,
            I => \ADC_VDC.bit_cnt_2\
        );

    \I__6078\ : InMux
    port map (
            O => \N__32566\,
            I => \N__32563\
        );

    \I__6077\ : LocalMux
    port map (
            O => \N__32563\,
            I => \ADC_VDC.n6_adj_1404\
        );

    \I__6076\ : CascadeMux
    port map (
            O => \N__32560\,
            I => \ADC_VDC.n11_cascade_\
        );

    \I__6075\ : InMux
    port map (
            O => \N__32557\,
            I => \N__32554\
        );

    \I__6074\ : LocalMux
    port map (
            O => \N__32554\,
            I => \ADC_VDC.n17359\
        );

    \I__6073\ : InMux
    port map (
            O => \N__32551\,
            I => \N__32548\
        );

    \I__6072\ : LocalMux
    port map (
            O => \N__32548\,
            I => \N__32543\
        );

    \I__6071\ : InMux
    port map (
            O => \N__32547\,
            I => \N__32538\
        );

    \I__6070\ : InMux
    port map (
            O => \N__32546\,
            I => \N__32535\
        );

    \I__6069\ : Span4Mux_h
    port map (
            O => \N__32543\,
            I => \N__32532\
        );

    \I__6068\ : InMux
    port map (
            O => \N__32542\,
            I => \N__32527\
        );

    \I__6067\ : InMux
    port map (
            O => \N__32541\,
            I => \N__32527\
        );

    \I__6066\ : LocalMux
    port map (
            O => \N__32538\,
            I => \ADC_VDC.bit_cnt_0\
        );

    \I__6065\ : LocalMux
    port map (
            O => \N__32535\,
            I => \ADC_VDC.bit_cnt_0\
        );

    \I__6064\ : Odrv4
    port map (
            O => \N__32532\,
            I => \ADC_VDC.bit_cnt_0\
        );

    \I__6063\ : LocalMux
    port map (
            O => \N__32527\,
            I => \ADC_VDC.bit_cnt_0\
        );

    \I__6062\ : InMux
    port map (
            O => \N__32518\,
            I => \bfn_13_6_0_\
        );

    \I__6061\ : InMux
    port map (
            O => \N__32515\,
            I => \N__32512\
        );

    \I__6060\ : LocalMux
    port map (
            O => \N__32512\,
            I => \N__32506\
        );

    \I__6059\ : CascadeMux
    port map (
            O => \N__32511\,
            I => \N__32502\
        );

    \I__6058\ : InMux
    port map (
            O => \N__32510\,
            I => \N__32499\
        );

    \I__6057\ : InMux
    port map (
            O => \N__32509\,
            I => \N__32496\
        );

    \I__6056\ : Span4Mux_h
    port map (
            O => \N__32506\,
            I => \N__32493\
        );

    \I__6055\ : InMux
    port map (
            O => \N__32505\,
            I => \N__32488\
        );

    \I__6054\ : InMux
    port map (
            O => \N__32502\,
            I => \N__32488\
        );

    \I__6053\ : LocalMux
    port map (
            O => \N__32499\,
            I => \ADC_VDC.bit_cnt_1\
        );

    \I__6052\ : LocalMux
    port map (
            O => \N__32496\,
            I => \ADC_VDC.bit_cnt_1\
        );

    \I__6051\ : Odrv4
    port map (
            O => \N__32493\,
            I => \ADC_VDC.bit_cnt_1\
        );

    \I__6050\ : LocalMux
    port map (
            O => \N__32488\,
            I => \ADC_VDC.bit_cnt_1\
        );

    \I__6049\ : InMux
    port map (
            O => \N__32479\,
            I => \ADC_VDC.n19469\
        );

    \I__6048\ : InMux
    port map (
            O => \N__32476\,
            I => \ADC_VDC.n19470\
        );

    \I__6047\ : InMux
    port map (
            O => \N__32473\,
            I => \ADC_VDC.n19471\
        );

    \I__6046\ : InMux
    port map (
            O => \N__32470\,
            I => \N__32467\
        );

    \I__6045\ : LocalMux
    port map (
            O => \N__32467\,
            I => \N__32460\
        );

    \I__6044\ : InMux
    port map (
            O => \N__32466\,
            I => \N__32457\
        );

    \I__6043\ : InMux
    port map (
            O => \N__32465\,
            I => \N__32450\
        );

    \I__6042\ : InMux
    port map (
            O => \N__32464\,
            I => \N__32450\
        );

    \I__6041\ : InMux
    port map (
            O => \N__32463\,
            I => \N__32450\
        );

    \I__6040\ : Span4Mux_h
    port map (
            O => \N__32460\,
            I => \N__32447\
        );

    \I__6039\ : LocalMux
    port map (
            O => \N__32457\,
            I => \ADC_VDC.bit_cnt_4\
        );

    \I__6038\ : LocalMux
    port map (
            O => \N__32450\,
            I => \ADC_VDC.bit_cnt_4\
        );

    \I__6037\ : Odrv4
    port map (
            O => \N__32447\,
            I => \ADC_VDC.bit_cnt_4\
        );

    \I__6036\ : InMux
    port map (
            O => \N__32440\,
            I => \ADC_VDC.n19472\
        );

    \I__6035\ : InMux
    port map (
            O => \N__32437\,
            I => \N__32432\
        );

    \I__6034\ : InMux
    port map (
            O => \N__32436\,
            I => \N__32429\
        );

    \I__6033\ : InMux
    port map (
            O => \N__32435\,
            I => \N__32426\
        );

    \I__6032\ : LocalMux
    port map (
            O => \N__32432\,
            I => \ADC_VDC.bit_cnt_5\
        );

    \I__6031\ : LocalMux
    port map (
            O => \N__32429\,
            I => \ADC_VDC.bit_cnt_5\
        );

    \I__6030\ : LocalMux
    port map (
            O => \N__32426\,
            I => \ADC_VDC.bit_cnt_5\
        );

    \I__6029\ : InMux
    port map (
            O => \N__32419\,
            I => \ADC_VDC.n19473\
        );

    \I__6028\ : CascadeMux
    port map (
            O => \N__32416\,
            I => \comm_spi.n22632_cascade_\
        );

    \I__6027\ : CascadeMux
    port map (
            O => \N__32413\,
            I => \comm_spi.imosi_cascade_\
        );

    \I__6026\ : InMux
    port map (
            O => \N__32410\,
            I => \N__32404\
        );

    \I__6025\ : InMux
    port map (
            O => \N__32409\,
            I => \N__32404\
        );

    \I__6024\ : LocalMux
    port map (
            O => \N__32404\,
            I => \comm_spi.imosi\
        );

    \I__6023\ : InMux
    port map (
            O => \N__32401\,
            I => \N__32398\
        );

    \I__6022\ : LocalMux
    port map (
            O => \N__32398\,
            I => \comm_spi.n14599\
        );

    \I__6021\ : SRMux
    port map (
            O => \N__32395\,
            I => \N__32392\
        );

    \I__6020\ : LocalMux
    port map (
            O => \N__32392\,
            I => \N__32389\
        );

    \I__6019\ : Span4Mux_h
    port map (
            O => \N__32389\,
            I => \N__32386\
        );

    \I__6018\ : Odrv4
    port map (
            O => \N__32386\,
            I => \comm_spi.DOUT_7__N_738\
        );

    \I__6017\ : InMux
    port map (
            O => \N__32383\,
            I => \N__32379\
        );

    \I__6016\ : InMux
    port map (
            O => \N__32382\,
            I => \N__32376\
        );

    \I__6015\ : LocalMux
    port map (
            O => \N__32379\,
            I => \ADC_VDC.genclk.n21167\
        );

    \I__6014\ : LocalMux
    port map (
            O => \N__32376\,
            I => \ADC_VDC.genclk.n21167\
        );

    \I__6013\ : InMux
    port map (
            O => \N__32371\,
            I => \N__32367\
        );

    \I__6012\ : CascadeMux
    port map (
            O => \N__32370\,
            I => \N__32363\
        );

    \I__6011\ : LocalMux
    port map (
            O => \N__32367\,
            I => \N__32360\
        );

    \I__6010\ : InMux
    port map (
            O => \N__32366\,
            I => \N__32355\
        );

    \I__6009\ : InMux
    port map (
            O => \N__32363\,
            I => \N__32355\
        );

    \I__6008\ : Odrv4
    port map (
            O => \N__32360\,
            I => buf_dds0_10
        );

    \I__6007\ : LocalMux
    port map (
            O => \N__32355\,
            I => buf_dds0_10
        );

    \I__6006\ : InMux
    port map (
            O => \N__32350\,
            I => \N__32347\
        );

    \I__6005\ : LocalMux
    port map (
            O => \N__32347\,
            I => \SIG_DDS.tmp_buf_10\
        );

    \I__6004\ : InMux
    port map (
            O => \N__32344\,
            I => \N__32341\
        );

    \I__6003\ : LocalMux
    port map (
            O => \N__32341\,
            I => \N__32338\
        );

    \I__6002\ : Span4Mux_h
    port map (
            O => \N__32338\,
            I => \N__32333\
        );

    \I__6001\ : InMux
    port map (
            O => \N__32337\,
            I => \N__32330\
        );

    \I__6000\ : InMux
    port map (
            O => \N__32336\,
            I => \N__32327\
        );

    \I__5999\ : Odrv4
    port map (
            O => \N__32333\,
            I => buf_dds0_9
        );

    \I__5998\ : LocalMux
    port map (
            O => \N__32330\,
            I => buf_dds0_9
        );

    \I__5997\ : LocalMux
    port map (
            O => \N__32327\,
            I => buf_dds0_9
        );

    \I__5996\ : CascadeMux
    port map (
            O => \N__32320\,
            I => \N__32317\
        );

    \I__5995\ : InMux
    port map (
            O => \N__32317\,
            I => \N__32314\
        );

    \I__5994\ : LocalMux
    port map (
            O => \N__32314\,
            I => \SIG_DDS.tmp_buf_9\
        );

    \I__5993\ : InMux
    port map (
            O => \N__32311\,
            I => \N__32307\
        );

    \I__5992\ : InMux
    port map (
            O => \N__32310\,
            I => \N__32304\
        );

    \I__5991\ : LocalMux
    port map (
            O => \N__32307\,
            I => \N__32301\
        );

    \I__5990\ : LocalMux
    port map (
            O => \N__32304\,
            I => \N__32297\
        );

    \I__5989\ : Span4Mux_h
    port map (
            O => \N__32301\,
            I => \N__32294\
        );

    \I__5988\ : InMux
    port map (
            O => \N__32300\,
            I => \N__32291\
        );

    \I__5987\ : Span4Mux_v
    port map (
            O => \N__32297\,
            I => \N__32288\
        );

    \I__5986\ : Odrv4
    port map (
            O => \N__32294\,
            I => buf_dds0_13
        );

    \I__5985\ : LocalMux
    port map (
            O => \N__32291\,
            I => buf_dds0_13
        );

    \I__5984\ : Odrv4
    port map (
            O => \N__32288\,
            I => buf_dds0_13
        );

    \I__5983\ : CascadeMux
    port map (
            O => \N__32281\,
            I => \N__32278\
        );

    \I__5982\ : InMux
    port map (
            O => \N__32278\,
            I => \N__32275\
        );

    \I__5981\ : LocalMux
    port map (
            O => \N__32275\,
            I => \SIG_DDS.tmp_buf_13\
        );

    \I__5980\ : CascadeMux
    port map (
            O => \N__32272\,
            I => \N__32268\
        );

    \I__5979\ : InMux
    port map (
            O => \N__32271\,
            I => \N__32265\
        );

    \I__5978\ : InMux
    port map (
            O => \N__32268\,
            I => \N__32262\
        );

    \I__5977\ : LocalMux
    port map (
            O => \N__32265\,
            I => \N__32259\
        );

    \I__5976\ : LocalMux
    port map (
            O => \N__32262\,
            I => \N__32255\
        );

    \I__5975\ : Span4Mux_v
    port map (
            O => \N__32259\,
            I => \N__32252\
        );

    \I__5974\ : InMux
    port map (
            O => \N__32258\,
            I => \N__32249\
        );

    \I__5973\ : Span4Mux_h
    port map (
            O => \N__32255\,
            I => \N__32246\
        );

    \I__5972\ : Odrv4
    port map (
            O => \N__32252\,
            I => buf_dds0_14
        );

    \I__5971\ : LocalMux
    port map (
            O => \N__32249\,
            I => buf_dds0_14
        );

    \I__5970\ : Odrv4
    port map (
            O => \N__32246\,
            I => buf_dds0_14
        );

    \I__5969\ : InMux
    port map (
            O => \N__32239\,
            I => \N__32235\
        );

    \I__5968\ : InMux
    port map (
            O => \N__32238\,
            I => \N__32232\
        );

    \I__5967\ : LocalMux
    port map (
            O => \N__32235\,
            I => \N__32228\
        );

    \I__5966\ : LocalMux
    port map (
            O => \N__32232\,
            I => \N__32225\
        );

    \I__5965\ : InMux
    port map (
            O => \N__32231\,
            I => \N__32222\
        );

    \I__5964\ : Span4Mux_v
    port map (
            O => \N__32228\,
            I => \N__32219\
        );

    \I__5963\ : Odrv4
    port map (
            O => \N__32225\,
            I => buf_dds0_1
        );

    \I__5962\ : LocalMux
    port map (
            O => \N__32222\,
            I => buf_dds0_1
        );

    \I__5961\ : Odrv4
    port map (
            O => \N__32219\,
            I => buf_dds0_1
        );

    \I__5960\ : CascadeMux
    port map (
            O => \N__32212\,
            I => \N__32209\
        );

    \I__5959\ : InMux
    port map (
            O => \N__32209\,
            I => \N__32206\
        );

    \I__5958\ : LocalMux
    port map (
            O => \N__32206\,
            I => \SIG_DDS.tmp_buf_7\
        );

    \I__5957\ : CascadeMux
    port map (
            O => \N__32203\,
            I => \N__32200\
        );

    \I__5956\ : InMux
    port map (
            O => \N__32200\,
            I => \N__32197\
        );

    \I__5955\ : LocalMux
    port map (
            O => \N__32197\,
            I => \SIG_DDS.tmp_buf_8\
        );

    \I__5954\ : InMux
    port map (
            O => \N__32194\,
            I => \N__32191\
        );

    \I__5953\ : LocalMux
    port map (
            O => \N__32191\,
            I => \comm_spi.n22629\
        );

    \I__5952\ : CascadeMux
    port map (
            O => \N__32188\,
            I => \comm_spi.n22629_cascade_\
        );

    \I__5951\ : CascadeMux
    port map (
            O => \N__32185\,
            I => \N__32182\
        );

    \I__5950\ : InMux
    port map (
            O => \N__32182\,
            I => \N__32173\
        );

    \I__5949\ : InMux
    port map (
            O => \N__32181\,
            I => \N__32173\
        );

    \I__5948\ : InMux
    port map (
            O => \N__32180\,
            I => \N__32170\
        );

    \I__5947\ : InMux
    port map (
            O => \N__32179\,
            I => \N__32165\
        );

    \I__5946\ : InMux
    port map (
            O => \N__32178\,
            I => \N__32165\
        );

    \I__5945\ : LocalMux
    port map (
            O => \N__32173\,
            I => \N__32152\
        );

    \I__5944\ : LocalMux
    port map (
            O => \N__32170\,
            I => \N__32147\
        );

    \I__5943\ : LocalMux
    port map (
            O => \N__32165\,
            I => \N__32147\
        );

    \I__5942\ : InMux
    port map (
            O => \N__32164\,
            I => \N__32138\
        );

    \I__5941\ : InMux
    port map (
            O => \N__32163\,
            I => \N__32138\
        );

    \I__5940\ : InMux
    port map (
            O => \N__32162\,
            I => \N__32138\
        );

    \I__5939\ : InMux
    port map (
            O => \N__32161\,
            I => \N__32138\
        );

    \I__5938\ : InMux
    port map (
            O => \N__32160\,
            I => \N__32131\
        );

    \I__5937\ : InMux
    port map (
            O => \N__32159\,
            I => \N__32131\
        );

    \I__5936\ : InMux
    port map (
            O => \N__32158\,
            I => \N__32131\
        );

    \I__5935\ : InMux
    port map (
            O => \N__32157\,
            I => \N__32128\
        );

    \I__5934\ : InMux
    port map (
            O => \N__32156\,
            I => \N__32125\
        );

    \I__5933\ : InMux
    port map (
            O => \N__32155\,
            I => \N__32122\
        );

    \I__5932\ : Span4Mux_v
    port map (
            O => \N__32152\,
            I => \N__32117\
        );

    \I__5931\ : Span4Mux_v
    port map (
            O => \N__32147\,
            I => \N__32117\
        );

    \I__5930\ : LocalMux
    port map (
            O => \N__32138\,
            I => \N__32108\
        );

    \I__5929\ : LocalMux
    port map (
            O => \N__32131\,
            I => \N__32108\
        );

    \I__5928\ : LocalMux
    port map (
            O => \N__32128\,
            I => \N__32108\
        );

    \I__5927\ : LocalMux
    port map (
            O => \N__32125\,
            I => \N__32108\
        );

    \I__5926\ : LocalMux
    port map (
            O => \N__32122\,
            I => \eis_end_N_716\
        );

    \I__5925\ : Odrv4
    port map (
            O => \N__32117\,
            I => \eis_end_N_716\
        );

    \I__5924\ : Odrv12
    port map (
            O => \N__32108\,
            I => \eis_end_N_716\
        );

    \I__5923\ : InMux
    port map (
            O => \N__32101\,
            I => \N__32096\
        );

    \I__5922\ : InMux
    port map (
            O => \N__32100\,
            I => \N__32091\
        );

    \I__5921\ : SRMux
    port map (
            O => \N__32099\,
            I => \N__32088\
        );

    \I__5920\ : LocalMux
    port map (
            O => \N__32096\,
            I => \N__32084\
        );

    \I__5919\ : InMux
    port map (
            O => \N__32095\,
            I => \N__32079\
        );

    \I__5918\ : InMux
    port map (
            O => \N__32094\,
            I => \N__32079\
        );

    \I__5917\ : LocalMux
    port map (
            O => \N__32091\,
            I => \N__32074\
        );

    \I__5916\ : LocalMux
    port map (
            O => \N__32088\,
            I => \N__32074\
        );

    \I__5915\ : CascadeMux
    port map (
            O => \N__32087\,
            I => \N__32071\
        );

    \I__5914\ : Span4Mux_h
    port map (
            O => \N__32084\,
            I => \N__32064\
        );

    \I__5913\ : LocalMux
    port map (
            O => \N__32079\,
            I => \N__32061\
        );

    \I__5912\ : Sp12to4
    port map (
            O => \N__32074\,
            I => \N__32058\
        );

    \I__5911\ : InMux
    port map (
            O => \N__32071\,
            I => \N__32055\
        );

    \I__5910\ : InMux
    port map (
            O => \N__32070\,
            I => \N__32052\
        );

    \I__5909\ : InMux
    port map (
            O => \N__32069\,
            I => \N__32045\
        );

    \I__5908\ : InMux
    port map (
            O => \N__32068\,
            I => \N__32045\
        );

    \I__5907\ : InMux
    port map (
            O => \N__32067\,
            I => \N__32045\
        );

    \I__5906\ : Odrv4
    port map (
            O => \N__32064\,
            I => acadc_rst
        );

    \I__5905\ : Odrv4
    port map (
            O => \N__32061\,
            I => acadc_rst
        );

    \I__5904\ : Odrv12
    port map (
            O => \N__32058\,
            I => acadc_rst
        );

    \I__5903\ : LocalMux
    port map (
            O => \N__32055\,
            I => acadc_rst
        );

    \I__5902\ : LocalMux
    port map (
            O => \N__32052\,
            I => acadc_rst
        );

    \I__5901\ : LocalMux
    port map (
            O => \N__32045\,
            I => acadc_rst
        );

    \I__5900\ : InMux
    port map (
            O => \N__32032\,
            I => \N__32029\
        );

    \I__5899\ : LocalMux
    port map (
            O => \N__32029\,
            I => \N__32026\
        );

    \I__5898\ : Span4Mux_v
    port map (
            O => \N__32026\,
            I => \N__32023\
        );

    \I__5897\ : Span4Mux_h
    port map (
            O => \N__32023\,
            I => \N__32020\
        );

    \I__5896\ : Odrv4
    port map (
            O => \N__32020\,
            I => buf_data_iac_15
        );

    \I__5895\ : InMux
    port map (
            O => \N__32017\,
            I => \N__32013\
        );

    \I__5894\ : InMux
    port map (
            O => \N__32016\,
            I => \N__32009\
        );

    \I__5893\ : LocalMux
    port map (
            O => \N__32013\,
            I => \N__32006\
        );

    \I__5892\ : InMux
    port map (
            O => \N__32012\,
            I => \N__32003\
        );

    \I__5891\ : LocalMux
    port map (
            O => \N__32009\,
            I => \N__31998\
        );

    \I__5890\ : Span4Mux_v
    port map (
            O => \N__32006\,
            I => \N__31998\
        );

    \I__5889\ : LocalMux
    port map (
            O => \N__32003\,
            I => \N__31995\
        );

    \I__5888\ : Odrv4
    port map (
            O => \N__31998\,
            I => buf_dds1_2
        );

    \I__5887\ : Odrv4
    port map (
            O => \N__31995\,
            I => buf_dds1_2
        );

    \I__5886\ : InMux
    port map (
            O => \N__31990\,
            I => \N__31987\
        );

    \I__5885\ : LocalMux
    port map (
            O => \N__31987\,
            I => \N__31983\
        );

    \I__5884\ : InMux
    port map (
            O => \N__31986\,
            I => \N__31980\
        );

    \I__5883\ : Span4Mux_v
    port map (
            O => \N__31983\,
            I => \N__31976\
        );

    \I__5882\ : LocalMux
    port map (
            O => \N__31980\,
            I => \N__31973\
        );

    \I__5881\ : InMux
    port map (
            O => \N__31979\,
            I => \N__31970\
        );

    \I__5880\ : Span4Mux_h
    port map (
            O => \N__31976\,
            I => \N__31965\
        );

    \I__5879\ : Span4Mux_h
    port map (
            O => \N__31973\,
            I => \N__31965\
        );

    \I__5878\ : LocalMux
    port map (
            O => \N__31970\,
            I => buf_adcdata_iac_15
        );

    \I__5877\ : Odrv4
    port map (
            O => \N__31965\,
            I => buf_adcdata_iac_15
        );

    \I__5876\ : InMux
    port map (
            O => \N__31960\,
            I => \N__31957\
        );

    \I__5875\ : LocalMux
    port map (
            O => \N__31957\,
            I => \N__31954\
        );

    \I__5874\ : Span12Mux_v
    port map (
            O => \N__31954\,
            I => \N__31951\
        );

    \I__5873\ : Odrv12
    port map (
            O => \N__31951\,
            I => n21961
        );

    \I__5872\ : CascadeMux
    port map (
            O => \N__31948\,
            I => \n16_adj_1621_cascade_\
        );

    \I__5871\ : InMux
    port map (
            O => \N__31945\,
            I => \N__31942\
        );

    \I__5870\ : LocalMux
    port map (
            O => \N__31942\,
            I => \N__31939\
        );

    \I__5869\ : Span4Mux_v
    port map (
            O => \N__31939\,
            I => \N__31936\
        );

    \I__5868\ : Odrv4
    port map (
            O => \N__31936\,
            I => n16_adj_1504
        );

    \I__5867\ : InMux
    port map (
            O => \N__31933\,
            I => \N__31928\
        );

    \I__5866\ : InMux
    port map (
            O => \N__31932\,
            I => \N__31925\
        );

    \I__5865\ : CascadeMux
    port map (
            O => \N__31931\,
            I => \N__31922\
        );

    \I__5864\ : LocalMux
    port map (
            O => \N__31928\,
            I => \N__31917\
        );

    \I__5863\ : LocalMux
    port map (
            O => \N__31925\,
            I => \N__31917\
        );

    \I__5862\ : InMux
    port map (
            O => \N__31922\,
            I => \N__31914\
        );

    \I__5861\ : Span4Mux_h
    port map (
            O => \N__31917\,
            I => \N__31911\
        );

    \I__5860\ : LocalMux
    port map (
            O => \N__31914\,
            I => buf_dds1_1
        );

    \I__5859\ : Odrv4
    port map (
            O => \N__31911\,
            I => buf_dds1_1
        );

    \I__5858\ : InMux
    port map (
            O => \N__31906\,
            I => \N__31899\
        );

    \I__5857\ : InMux
    port map (
            O => \N__31905\,
            I => \N__31899\
        );

    \I__5856\ : InMux
    port map (
            O => \N__31904\,
            I => \N__31896\
        );

    \I__5855\ : LocalMux
    port map (
            O => \N__31899\,
            I => \acadc_skipCount_6\
        );

    \I__5854\ : LocalMux
    port map (
            O => \N__31896\,
            I => \acadc_skipCount_6\
        );

    \I__5853\ : InMux
    port map (
            O => \N__31891\,
            I => \N__31888\
        );

    \I__5852\ : LocalMux
    port map (
            O => \N__31888\,
            I => n17
        );

    \I__5851\ : InMux
    port map (
            O => \N__31885\,
            I => \N__31879\
        );

    \I__5850\ : InMux
    port map (
            O => \N__31884\,
            I => \N__31876\
        );

    \I__5849\ : InMux
    port map (
            O => \N__31883\,
            I => \N__31873\
        );

    \I__5848\ : InMux
    port map (
            O => \N__31882\,
            I => \N__31870\
        );

    \I__5847\ : LocalMux
    port map (
            O => \N__31879\,
            I => acadc_dtrig_v
        );

    \I__5846\ : LocalMux
    port map (
            O => \N__31876\,
            I => acadc_dtrig_v
        );

    \I__5845\ : LocalMux
    port map (
            O => \N__31873\,
            I => acadc_dtrig_v
        );

    \I__5844\ : LocalMux
    port map (
            O => \N__31870\,
            I => acadc_dtrig_v
        );

    \I__5843\ : InMux
    port map (
            O => \N__31861\,
            I => \N__31855\
        );

    \I__5842\ : InMux
    port map (
            O => \N__31860\,
            I => \N__31852\
        );

    \I__5841\ : InMux
    port map (
            O => \N__31859\,
            I => \N__31847\
        );

    \I__5840\ : InMux
    port map (
            O => \N__31858\,
            I => \N__31847\
        );

    \I__5839\ : LocalMux
    port map (
            O => \N__31855\,
            I => acadc_dtrig_i
        );

    \I__5838\ : LocalMux
    port map (
            O => \N__31852\,
            I => acadc_dtrig_i
        );

    \I__5837\ : LocalMux
    port map (
            O => \N__31847\,
            I => acadc_dtrig_i
        );

    \I__5836\ : CascadeMux
    port map (
            O => \N__31840\,
            I => \iac_raw_buf_N_728_cascade_\
        );

    \I__5835\ : InMux
    port map (
            O => \N__31837\,
            I => \N__31834\
        );

    \I__5834\ : LocalMux
    port map (
            O => \N__31834\,
            I => \N__31831\
        );

    \I__5833\ : Odrv4
    port map (
            O => \N__31831\,
            I => n21997
        );

    \I__5832\ : InMux
    port map (
            O => \N__31828\,
            I => \N__31824\
        );

    \I__5831\ : InMux
    port map (
            O => \N__31827\,
            I => \N__31821\
        );

    \I__5830\ : LocalMux
    port map (
            O => \N__31824\,
            I => \N__31815\
        );

    \I__5829\ : LocalMux
    port map (
            O => \N__31821\,
            I => \N__31815\
        );

    \I__5828\ : InMux
    port map (
            O => \N__31820\,
            I => \N__31812\
        );

    \I__5827\ : Span4Mux_h
    port map (
            O => \N__31815\,
            I => \N__31809\
        );

    \I__5826\ : LocalMux
    port map (
            O => \N__31812\,
            I => buf_dds1_3
        );

    \I__5825\ : Odrv4
    port map (
            O => \N__31809\,
            I => buf_dds1_3
        );

    \I__5824\ : InMux
    port map (
            O => \N__31804\,
            I => \N__31801\
        );

    \I__5823\ : LocalMux
    port map (
            O => \N__31801\,
            I => \N__31798\
        );

    \I__5822\ : Span12Mux_h
    port map (
            O => \N__31798\,
            I => \N__31795\
        );

    \I__5821\ : Odrv12
    port map (
            O => \N__31795\,
            I => n20624
        );

    \I__5820\ : CascadeMux
    port map (
            O => \N__31792\,
            I => \n12353_cascade_\
        );

    \I__5819\ : CascadeMux
    port map (
            O => \N__31789\,
            I => \N__31786\
        );

    \I__5818\ : InMux
    port map (
            O => \N__31786\,
            I => \N__31783\
        );

    \I__5817\ : LocalMux
    port map (
            O => \N__31783\,
            I => \N__31780\
        );

    \I__5816\ : Odrv4
    port map (
            O => \N__31780\,
            I => n35
        );

    \I__5815\ : SRMux
    port map (
            O => \N__31777\,
            I => \N__31773\
        );

    \I__5814\ : SRMux
    port map (
            O => \N__31776\,
            I => \N__31770\
        );

    \I__5813\ : LocalMux
    port map (
            O => \N__31773\,
            I => \N__31763\
        );

    \I__5812\ : LocalMux
    port map (
            O => \N__31770\,
            I => \N__31760\
        );

    \I__5811\ : SRMux
    port map (
            O => \N__31769\,
            I => \N__31757\
        );

    \I__5810\ : SRMux
    port map (
            O => \N__31768\,
            I => \N__31754\
        );

    \I__5809\ : SRMux
    port map (
            O => \N__31767\,
            I => \N__31747\
        );

    \I__5808\ : SRMux
    port map (
            O => \N__31766\,
            I => \N__31744\
        );

    \I__5807\ : Span4Mux_h
    port map (
            O => \N__31763\,
            I => \N__31741\
        );

    \I__5806\ : Span4Mux_v
    port map (
            O => \N__31760\,
            I => \N__31736\
        );

    \I__5805\ : LocalMux
    port map (
            O => \N__31757\,
            I => \N__31736\
        );

    \I__5804\ : LocalMux
    port map (
            O => \N__31754\,
            I => \N__31733\
        );

    \I__5803\ : SRMux
    port map (
            O => \N__31753\,
            I => \N__31730\
        );

    \I__5802\ : SRMux
    port map (
            O => \N__31752\,
            I => \N__31727\
        );

    \I__5801\ : SRMux
    port map (
            O => \N__31751\,
            I => \N__31723\
        );

    \I__5800\ : SRMux
    port map (
            O => \N__31750\,
            I => \N__31720\
        );

    \I__5799\ : LocalMux
    port map (
            O => \N__31747\,
            I => \N__31716\
        );

    \I__5798\ : LocalMux
    port map (
            O => \N__31744\,
            I => \N__31713\
        );

    \I__5797\ : Span4Mux_v
    port map (
            O => \N__31741\,
            I => \N__31708\
        );

    \I__5796\ : Span4Mux_h
    port map (
            O => \N__31736\,
            I => \N__31708\
        );

    \I__5795\ : Span4Mux_v
    port map (
            O => \N__31733\,
            I => \N__31703\
        );

    \I__5794\ : LocalMux
    port map (
            O => \N__31730\,
            I => \N__31703\
        );

    \I__5793\ : LocalMux
    port map (
            O => \N__31727\,
            I => \N__31700\
        );

    \I__5792\ : SRMux
    port map (
            O => \N__31726\,
            I => \N__31697\
        );

    \I__5791\ : LocalMux
    port map (
            O => \N__31723\,
            I => \N__31694\
        );

    \I__5790\ : LocalMux
    port map (
            O => \N__31720\,
            I => \N__31691\
        );

    \I__5789\ : SRMux
    port map (
            O => \N__31719\,
            I => \N__31688\
        );

    \I__5788\ : Span4Mux_v
    port map (
            O => \N__31716\,
            I => \N__31685\
        );

    \I__5787\ : Span4Mux_h
    port map (
            O => \N__31713\,
            I => \N__31682\
        );

    \I__5786\ : Span4Mux_v
    port map (
            O => \N__31708\,
            I => \N__31677\
        );

    \I__5785\ : Span4Mux_h
    port map (
            O => \N__31703\,
            I => \N__31677\
        );

    \I__5784\ : Span4Mux_v
    port map (
            O => \N__31700\,
            I => \N__31672\
        );

    \I__5783\ : LocalMux
    port map (
            O => \N__31697\,
            I => \N__31672\
        );

    \I__5782\ : Span4Mux_v
    port map (
            O => \N__31694\,
            I => \N__31665\
        );

    \I__5781\ : Span4Mux_v
    port map (
            O => \N__31691\,
            I => \N__31665\
        );

    \I__5780\ : LocalMux
    port map (
            O => \N__31688\,
            I => \N__31665\
        );

    \I__5779\ : Span4Mux_h
    port map (
            O => \N__31685\,
            I => \N__31662\
        );

    \I__5778\ : Span4Mux_h
    port map (
            O => \N__31682\,
            I => \N__31659\
        );

    \I__5777\ : Span4Mux_v
    port map (
            O => \N__31677\,
            I => \N__31654\
        );

    \I__5776\ : Span4Mux_h
    port map (
            O => \N__31672\,
            I => \N__31654\
        );

    \I__5775\ : Span4Mux_h
    port map (
            O => \N__31665\,
            I => \N__31651\
        );

    \I__5774\ : Span4Mux_h
    port map (
            O => \N__31662\,
            I => \N__31648\
        );

    \I__5773\ : Span4Mux_h
    port map (
            O => \N__31659\,
            I => \N__31641\
        );

    \I__5772\ : Span4Mux_h
    port map (
            O => \N__31654\,
            I => \N__31641\
        );

    \I__5771\ : Span4Mux_h
    port map (
            O => \N__31651\,
            I => \N__31641\
        );

    \I__5770\ : Odrv4
    port map (
            O => \N__31648\,
            I => \iac_raw_buf_N_726\
        );

    \I__5769\ : Odrv4
    port map (
            O => \N__31641\,
            I => \iac_raw_buf_N_726\
        );

    \I__5768\ : CascadeMux
    port map (
            O => \N__31636\,
            I => \N__31633\
        );

    \I__5767\ : CascadeBuf
    port map (
            O => \N__31633\,
            I => \N__31630\
        );

    \I__5766\ : CascadeMux
    port map (
            O => \N__31630\,
            I => \N__31627\
        );

    \I__5765\ : CascadeBuf
    port map (
            O => \N__31627\,
            I => \N__31624\
        );

    \I__5764\ : CascadeMux
    port map (
            O => \N__31624\,
            I => \N__31621\
        );

    \I__5763\ : CascadeBuf
    port map (
            O => \N__31621\,
            I => \N__31618\
        );

    \I__5762\ : CascadeMux
    port map (
            O => \N__31618\,
            I => \N__31615\
        );

    \I__5761\ : CascadeBuf
    port map (
            O => \N__31615\,
            I => \N__31612\
        );

    \I__5760\ : CascadeMux
    port map (
            O => \N__31612\,
            I => \N__31609\
        );

    \I__5759\ : CascadeBuf
    port map (
            O => \N__31609\,
            I => \N__31606\
        );

    \I__5758\ : CascadeMux
    port map (
            O => \N__31606\,
            I => \N__31603\
        );

    \I__5757\ : CascadeBuf
    port map (
            O => \N__31603\,
            I => \N__31600\
        );

    \I__5756\ : CascadeMux
    port map (
            O => \N__31600\,
            I => \N__31597\
        );

    \I__5755\ : CascadeBuf
    port map (
            O => \N__31597\,
            I => \N__31594\
        );

    \I__5754\ : CascadeMux
    port map (
            O => \N__31594\,
            I => \N__31591\
        );

    \I__5753\ : CascadeBuf
    port map (
            O => \N__31591\,
            I => \N__31588\
        );

    \I__5752\ : CascadeMux
    port map (
            O => \N__31588\,
            I => \N__31584\
        );

    \I__5751\ : CascadeMux
    port map (
            O => \N__31587\,
            I => \N__31581\
        );

    \I__5750\ : CascadeBuf
    port map (
            O => \N__31584\,
            I => \N__31578\
        );

    \I__5749\ : CascadeBuf
    port map (
            O => \N__31581\,
            I => \N__31575\
        );

    \I__5748\ : CascadeMux
    port map (
            O => \N__31578\,
            I => \N__31572\
        );

    \I__5747\ : CascadeMux
    port map (
            O => \N__31575\,
            I => \N__31569\
        );

    \I__5746\ : InMux
    port map (
            O => \N__31572\,
            I => \N__31566\
        );

    \I__5745\ : InMux
    port map (
            O => \N__31569\,
            I => \N__31563\
        );

    \I__5744\ : LocalMux
    port map (
            O => \N__31566\,
            I => \N__31560\
        );

    \I__5743\ : LocalMux
    port map (
            O => \N__31563\,
            I => \N__31557\
        );

    \I__5742\ : Span4Mux_h
    port map (
            O => \N__31560\,
            I => \N__31554\
        );

    \I__5741\ : Span4Mux_v
    port map (
            O => \N__31557\,
            I => \N__31551\
        );

    \I__5740\ : Span4Mux_h
    port map (
            O => \N__31554\,
            I => \N__31548\
        );

    \I__5739\ : Sp12to4
    port map (
            O => \N__31551\,
            I => \N__31545\
        );

    \I__5738\ : Span4Mux_v
    port map (
            O => \N__31548\,
            I => \N__31542\
        );

    \I__5737\ : Odrv12
    port map (
            O => \N__31545\,
            I => \data_index_9_N_212_0\
        );

    \I__5736\ : Odrv4
    port map (
            O => \N__31542\,
            I => \data_index_9_N_212_0\
        );

    \I__5735\ : InMux
    port map (
            O => \N__31537\,
            I => \N__31534\
        );

    \I__5734\ : LocalMux
    port map (
            O => \N__31534\,
            I => \N__31530\
        );

    \I__5733\ : InMux
    port map (
            O => \N__31533\,
            I => \N__31526\
        );

    \I__5732\ : Span4Mux_h
    port map (
            O => \N__31530\,
            I => \N__31523\
        );

    \I__5731\ : InMux
    port map (
            O => \N__31529\,
            I => \N__31520\
        );

    \I__5730\ : LocalMux
    port map (
            O => \N__31526\,
            I => \acadc_skipCount_8\
        );

    \I__5729\ : Odrv4
    port map (
            O => \N__31523\,
            I => \acadc_skipCount_8\
        );

    \I__5728\ : LocalMux
    port map (
            O => \N__31520\,
            I => \acadc_skipCount_8\
        );

    \I__5727\ : CascadeMux
    port map (
            O => \N__31513\,
            I => \n20_cascade_\
        );

    \I__5726\ : InMux
    port map (
            O => \N__31510\,
            I => \N__31507\
        );

    \I__5725\ : LocalMux
    port map (
            O => \N__31507\,
            I => \N__31504\
        );

    \I__5724\ : Odrv4
    port map (
            O => \N__31504\,
            I => n14_adj_1498
        );

    \I__5723\ : InMux
    port map (
            O => \N__31501\,
            I => \N__31498\
        );

    \I__5722\ : LocalMux
    port map (
            O => \N__31498\,
            I => \N__31495\
        );

    \I__5721\ : Odrv4
    port map (
            O => \N__31495\,
            I => n18_adj_1587
        );

    \I__5720\ : CascadeMux
    port map (
            O => \N__31492\,
            I => \n26_adj_1604_cascade_\
        );

    \I__5719\ : InMux
    port map (
            O => \N__31489\,
            I => \N__31483\
        );

    \I__5718\ : InMux
    port map (
            O => \N__31488\,
            I => \N__31483\
        );

    \I__5717\ : LocalMux
    port map (
            O => \N__31483\,
            I => \N__31480\
        );

    \I__5716\ : Odrv4
    port map (
            O => \N__31480\,
            I => n31
        );

    \I__5715\ : CascadeMux
    port map (
            O => \N__31477\,
            I => \N__31474\
        );

    \I__5714\ : CascadeBuf
    port map (
            O => \N__31474\,
            I => \N__31471\
        );

    \I__5713\ : CascadeMux
    port map (
            O => \N__31471\,
            I => \N__31468\
        );

    \I__5712\ : CascadeBuf
    port map (
            O => \N__31468\,
            I => \N__31465\
        );

    \I__5711\ : CascadeMux
    port map (
            O => \N__31465\,
            I => \N__31462\
        );

    \I__5710\ : CascadeBuf
    port map (
            O => \N__31462\,
            I => \N__31459\
        );

    \I__5709\ : CascadeMux
    port map (
            O => \N__31459\,
            I => \N__31456\
        );

    \I__5708\ : CascadeBuf
    port map (
            O => \N__31456\,
            I => \N__31453\
        );

    \I__5707\ : CascadeMux
    port map (
            O => \N__31453\,
            I => \N__31450\
        );

    \I__5706\ : CascadeBuf
    port map (
            O => \N__31450\,
            I => \N__31447\
        );

    \I__5705\ : CascadeMux
    port map (
            O => \N__31447\,
            I => \N__31444\
        );

    \I__5704\ : CascadeBuf
    port map (
            O => \N__31444\,
            I => \N__31441\
        );

    \I__5703\ : CascadeMux
    port map (
            O => \N__31441\,
            I => \N__31438\
        );

    \I__5702\ : CascadeBuf
    port map (
            O => \N__31438\,
            I => \N__31435\
        );

    \I__5701\ : CascadeMux
    port map (
            O => \N__31435\,
            I => \N__31431\
        );

    \I__5700\ : CascadeMux
    port map (
            O => \N__31434\,
            I => \N__31428\
        );

    \I__5699\ : CascadeBuf
    port map (
            O => \N__31431\,
            I => \N__31425\
        );

    \I__5698\ : CascadeBuf
    port map (
            O => \N__31428\,
            I => \N__31422\
        );

    \I__5697\ : CascadeMux
    port map (
            O => \N__31425\,
            I => \N__31419\
        );

    \I__5696\ : CascadeMux
    port map (
            O => \N__31422\,
            I => \N__31416\
        );

    \I__5695\ : CascadeBuf
    port map (
            O => \N__31419\,
            I => \N__31413\
        );

    \I__5694\ : InMux
    port map (
            O => \N__31416\,
            I => \N__31410\
        );

    \I__5693\ : CascadeMux
    port map (
            O => \N__31413\,
            I => \N__31407\
        );

    \I__5692\ : LocalMux
    port map (
            O => \N__31410\,
            I => \N__31404\
        );

    \I__5691\ : InMux
    port map (
            O => \N__31407\,
            I => \N__31401\
        );

    \I__5690\ : Span4Mux_v
    port map (
            O => \N__31404\,
            I => \N__31398\
        );

    \I__5689\ : LocalMux
    port map (
            O => \N__31401\,
            I => \N__31395\
        );

    \I__5688\ : Span4Mux_h
    port map (
            O => \N__31398\,
            I => \N__31392\
        );

    \I__5687\ : Span4Mux_v
    port map (
            O => \N__31395\,
            I => \N__31389\
        );

    \I__5686\ : Span4Mux_h
    port map (
            O => \N__31392\,
            I => \N__31384\
        );

    \I__5685\ : Span4Mux_h
    port map (
            O => \N__31389\,
            I => \N__31384\
        );

    \I__5684\ : Odrv4
    port map (
            O => \N__31384\,
            I => \data_index_9_N_212_3\
        );

    \I__5683\ : CascadeMux
    port map (
            O => \N__31381\,
            I => \N__31378\
        );

    \I__5682\ : InMux
    port map (
            O => \N__31378\,
            I => \N__31373\
        );

    \I__5681\ : InMux
    port map (
            O => \N__31377\,
            I => \N__31370\
        );

    \I__5680\ : InMux
    port map (
            O => \N__31376\,
            I => \N__31367\
        );

    \I__5679\ : LocalMux
    port map (
            O => \N__31373\,
            I => \N__31364\
        );

    \I__5678\ : LocalMux
    port map (
            O => \N__31370\,
            I => \acadc_skipCount_5\
        );

    \I__5677\ : LocalMux
    port map (
            O => \N__31367\,
            I => \acadc_skipCount_5\
        );

    \I__5676\ : Odrv4
    port map (
            O => \N__31364\,
            I => \acadc_skipCount_5\
        );

    \I__5675\ : InMux
    port map (
            O => \N__31357\,
            I => \N__31353\
        );

    \I__5674\ : InMux
    port map (
            O => \N__31356\,
            I => \N__31350\
        );

    \I__5673\ : LocalMux
    port map (
            O => \N__31353\,
            I => \N__31347\
        );

    \I__5672\ : LocalMux
    port map (
            O => \N__31350\,
            I => data_idxvec_13
        );

    \I__5671\ : Odrv4
    port map (
            O => \N__31347\,
            I => data_idxvec_13
        );

    \I__5670\ : InMux
    port map (
            O => \N__31342\,
            I => n19347
        );

    \I__5669\ : CascadeMux
    port map (
            O => \N__31339\,
            I => \N__31336\
        );

    \I__5668\ : InMux
    port map (
            O => \N__31336\,
            I => \N__31333\
        );

    \I__5667\ : LocalMux
    port map (
            O => \N__31333\,
            I => \N__31329\
        );

    \I__5666\ : CascadeMux
    port map (
            O => \N__31332\,
            I => \N__31326\
        );

    \I__5665\ : Span4Mux_h
    port map (
            O => \N__31329\,
            I => \N__31323\
        );

    \I__5664\ : InMux
    port map (
            O => \N__31326\,
            I => \N__31320\
        );

    \I__5663\ : Span4Mux_v
    port map (
            O => \N__31323\,
            I => \N__31317\
        );

    \I__5662\ : LocalMux
    port map (
            O => \N__31320\,
            I => data_idxvec_14
        );

    \I__5661\ : Odrv4
    port map (
            O => \N__31317\,
            I => data_idxvec_14
        );

    \I__5660\ : InMux
    port map (
            O => \N__31312\,
            I => n19348
        );

    \I__5659\ : InMux
    port map (
            O => \N__31309\,
            I => n19349
        );

    \I__5658\ : InMux
    port map (
            O => \N__31306\,
            I => \N__31303\
        );

    \I__5657\ : LocalMux
    port map (
            O => \N__31303\,
            I => \N__31299\
        );

    \I__5656\ : InMux
    port map (
            O => \N__31302\,
            I => \N__31296\
        );

    \I__5655\ : Span4Mux_h
    port map (
            O => \N__31299\,
            I => \N__31293\
        );

    \I__5654\ : LocalMux
    port map (
            O => \N__31296\,
            I => data_idxvec_15
        );

    \I__5653\ : Odrv4
    port map (
            O => \N__31293\,
            I => data_idxvec_15
        );

    \I__5652\ : InMux
    port map (
            O => \N__31288\,
            I => \N__31284\
        );

    \I__5651\ : InMux
    port map (
            O => \N__31287\,
            I => \N__31281\
        );

    \I__5650\ : LocalMux
    port map (
            O => \N__31284\,
            I => \N__31278\
        );

    \I__5649\ : LocalMux
    port map (
            O => \N__31281\,
            I => data_idxvec_5
        );

    \I__5648\ : Odrv4
    port map (
            O => \N__31278\,
            I => data_idxvec_5
        );

    \I__5647\ : CascadeMux
    port map (
            O => \N__31273\,
            I => \n26_adj_1486_cascade_\
        );

    \I__5646\ : CascadeMux
    port map (
            O => \N__31270\,
            I => \n22177_cascade_\
        );

    \I__5645\ : InMux
    port map (
            O => \N__31267\,
            I => \N__31264\
        );

    \I__5644\ : LocalMux
    port map (
            O => \N__31264\,
            I => \N__31261\
        );

    \I__5643\ : Span4Mux_v
    port map (
            O => \N__31261\,
            I => \N__31258\
        );

    \I__5642\ : Odrv4
    port map (
            O => \N__31258\,
            I => n22120
        );

    \I__5641\ : CascadeMux
    port map (
            O => \N__31255\,
            I => \n22180_cascade_\
        );

    \I__5640\ : CascadeMux
    port map (
            O => \N__31252\,
            I => \n30_adj_1485_cascade_\
        );

    \I__5639\ : InMux
    port map (
            O => \N__31249\,
            I => \N__31246\
        );

    \I__5638\ : LocalMux
    port map (
            O => \N__31246\,
            I => \N__31243\
        );

    \I__5637\ : Span4Mux_h
    port map (
            O => \N__31243\,
            I => \N__31240\
        );

    \I__5636\ : Span4Mux_h
    port map (
            O => \N__31240\,
            I => \N__31237\
        );

    \I__5635\ : Odrv4
    port map (
            O => \N__31237\,
            I => buf_data_iac_13
        );

    \I__5634\ : InMux
    port map (
            O => \N__31234\,
            I => \N__31231\
        );

    \I__5633\ : LocalMux
    port map (
            O => \N__31231\,
            I => n21036
        );

    \I__5632\ : InMux
    port map (
            O => \N__31228\,
            I => n19338
        );

    \I__5631\ : InMux
    port map (
            O => \N__31225\,
            I => n19339
        );

    \I__5630\ : InMux
    port map (
            O => \N__31222\,
            I => \N__31218\
        );

    \I__5629\ : InMux
    port map (
            O => \N__31221\,
            I => \N__31215\
        );

    \I__5628\ : LocalMux
    port map (
            O => \N__31218\,
            I => \N__31212\
        );

    \I__5627\ : LocalMux
    port map (
            O => \N__31215\,
            I => data_idxvec_6
        );

    \I__5626\ : Odrv4
    port map (
            O => \N__31212\,
            I => data_idxvec_6
        );

    \I__5625\ : InMux
    port map (
            O => \N__31207\,
            I => n19340
        );

    \I__5624\ : InMux
    port map (
            O => \N__31204\,
            I => n19341
        );

    \I__5623\ : InMux
    port map (
            O => \N__31201\,
            I => \bfn_12_13_0_\
        );

    \I__5622\ : InMux
    port map (
            O => \N__31198\,
            I => \N__31195\
        );

    \I__5621\ : LocalMux
    port map (
            O => \N__31195\,
            I => \N__31191\
        );

    \I__5620\ : InMux
    port map (
            O => \N__31194\,
            I => \N__31188\
        );

    \I__5619\ : Span4Mux_v
    port map (
            O => \N__31191\,
            I => \N__31185\
        );

    \I__5618\ : LocalMux
    port map (
            O => \N__31188\,
            I => data_idxvec_9
        );

    \I__5617\ : Odrv4
    port map (
            O => \N__31185\,
            I => data_idxvec_9
        );

    \I__5616\ : InMux
    port map (
            O => \N__31180\,
            I => n19343
        );

    \I__5615\ : CascadeMux
    port map (
            O => \N__31177\,
            I => \N__31173\
        );

    \I__5614\ : InMux
    port map (
            O => \N__31176\,
            I => \N__31170\
        );

    \I__5613\ : InMux
    port map (
            O => \N__31173\,
            I => \N__31167\
        );

    \I__5612\ : LocalMux
    port map (
            O => \N__31170\,
            I => \N__31164\
        );

    \I__5611\ : LocalMux
    port map (
            O => \N__31167\,
            I => \N__31159\
        );

    \I__5610\ : Span4Mux_v
    port map (
            O => \N__31164\,
            I => \N__31159\
        );

    \I__5609\ : Odrv4
    port map (
            O => \N__31159\,
            I => data_idxvec_10
        );

    \I__5608\ : InMux
    port map (
            O => \N__31156\,
            I => n19344
        );

    \I__5607\ : InMux
    port map (
            O => \N__31153\,
            I => n19345
        );

    \I__5606\ : CascadeMux
    port map (
            O => \N__31150\,
            I => \N__31147\
        );

    \I__5605\ : InMux
    port map (
            O => \N__31147\,
            I => \N__31143\
        );

    \I__5604\ : CascadeMux
    port map (
            O => \N__31146\,
            I => \N__31140\
        );

    \I__5603\ : LocalMux
    port map (
            O => \N__31143\,
            I => \N__31137\
        );

    \I__5602\ : InMux
    port map (
            O => \N__31140\,
            I => \N__31134\
        );

    \I__5601\ : Span4Mux_h
    port map (
            O => \N__31137\,
            I => \N__31131\
        );

    \I__5600\ : LocalMux
    port map (
            O => \N__31134\,
            I => data_idxvec_12
        );

    \I__5599\ : Odrv4
    port map (
            O => \N__31131\,
            I => data_idxvec_12
        );

    \I__5598\ : InMux
    port map (
            O => \N__31126\,
            I => n19346
        );

    \I__5597\ : InMux
    port map (
            O => \N__31123\,
            I => \N__31120\
        );

    \I__5596\ : LocalMux
    port map (
            O => \N__31120\,
            I => \N__31117\
        );

    \I__5595\ : Span4Mux_h
    port map (
            O => \N__31117\,
            I => \N__31114\
        );

    \I__5594\ : Span4Mux_v
    port map (
            O => \N__31114\,
            I => \N__31111\
        );

    \I__5593\ : Span4Mux_h
    port map (
            O => \N__31111\,
            I => \N__31108\
        );

    \I__5592\ : Odrv4
    port map (
            O => \N__31108\,
            I => buf_data_vac_13
        );

    \I__5591\ : InMux
    port map (
            O => \N__31105\,
            I => \N__31102\
        );

    \I__5590\ : LocalMux
    port map (
            O => \N__31102\,
            I => \N__31099\
        );

    \I__5589\ : Span4Mux_h
    port map (
            O => \N__31099\,
            I => \N__31096\
        );

    \I__5588\ : Span4Mux_v
    port map (
            O => \N__31096\,
            I => \N__31093\
        );

    \I__5587\ : Span4Mux_h
    port map (
            O => \N__31093\,
            I => \N__31090\
        );

    \I__5586\ : Odrv4
    port map (
            O => \N__31090\,
            I => buf_data_vac_12
        );

    \I__5585\ : InMux
    port map (
            O => \N__31087\,
            I => \N__31084\
        );

    \I__5584\ : LocalMux
    port map (
            O => \N__31084\,
            I => \N__31081\
        );

    \I__5583\ : Span4Mux_h
    port map (
            O => \N__31081\,
            I => \N__31078\
        );

    \I__5582\ : Span4Mux_h
    port map (
            O => \N__31078\,
            I => \N__31075\
        );

    \I__5581\ : Span4Mux_v
    port map (
            O => \N__31075\,
            I => \N__31072\
        );

    \I__5580\ : Odrv4
    port map (
            O => \N__31072\,
            I => buf_data_vac_11
        );

    \I__5579\ : InMux
    port map (
            O => \N__31069\,
            I => \N__31066\
        );

    \I__5578\ : LocalMux
    port map (
            O => \N__31066\,
            I => \N__31063\
        );

    \I__5577\ : Span4Mux_v
    port map (
            O => \N__31063\,
            I => \N__31060\
        );

    \I__5576\ : Span4Mux_v
    port map (
            O => \N__31060\,
            I => \N__31057\
        );

    \I__5575\ : Span4Mux_h
    port map (
            O => \N__31057\,
            I => \N__31054\
        );

    \I__5574\ : Span4Mux_h
    port map (
            O => \N__31054\,
            I => \N__31051\
        );

    \I__5573\ : Odrv4
    port map (
            O => \N__31051\,
            I => buf_data_vac_10
        );

    \I__5572\ : InMux
    port map (
            O => \N__31048\,
            I => \N__31045\
        );

    \I__5571\ : LocalMux
    port map (
            O => \N__31045\,
            I => \N__31042\
        );

    \I__5570\ : Span4Mux_h
    port map (
            O => \N__31042\,
            I => \N__31039\
        );

    \I__5569\ : Span4Mux_v
    port map (
            O => \N__31039\,
            I => \N__31036\
        );

    \I__5568\ : Span4Mux_v
    port map (
            O => \N__31036\,
            I => \N__31033\
        );

    \I__5567\ : Span4Mux_h
    port map (
            O => \N__31033\,
            I => \N__31030\
        );

    \I__5566\ : Odrv4
    port map (
            O => \N__31030\,
            I => buf_data_vac_9
        );

    \I__5565\ : InMux
    port map (
            O => \N__31027\,
            I => \N__31024\
        );

    \I__5564\ : LocalMux
    port map (
            O => \N__31024\,
            I => \N__31021\
        );

    \I__5563\ : Span4Mux_h
    port map (
            O => \N__31021\,
            I => \N__31018\
        );

    \I__5562\ : Span4Mux_h
    port map (
            O => \N__31018\,
            I => \N__31015\
        );

    \I__5561\ : Odrv4
    port map (
            O => \N__31015\,
            I => n14_adj_1516
        );

    \I__5560\ : InMux
    port map (
            O => \N__31012\,
            I => \bfn_12_12_0_\
        );

    \I__5559\ : InMux
    port map (
            O => \N__31009\,
            I => n19335
        );

    \I__5558\ : InMux
    port map (
            O => \N__31006\,
            I => n19336
        );

    \I__5557\ : InMux
    port map (
            O => \N__31003\,
            I => n19337
        );

    \I__5556\ : InMux
    port map (
            O => \N__31000\,
            I => \N__30994\
        );

    \I__5555\ : InMux
    port map (
            O => \N__30999\,
            I => \N__30994\
        );

    \I__5554\ : LocalMux
    port map (
            O => \N__30994\,
            I => \N__30986\
        );

    \I__5553\ : CascadeMux
    port map (
            O => \N__30993\,
            I => \N__30983\
        );

    \I__5552\ : InMux
    port map (
            O => \N__30992\,
            I => \N__30980\
        );

    \I__5551\ : InMux
    port map (
            O => \N__30991\,
            I => \N__30977\
        );

    \I__5550\ : InMux
    port map (
            O => \N__30990\,
            I => \N__30972\
        );

    \I__5549\ : InMux
    port map (
            O => \N__30989\,
            I => \N__30972\
        );

    \I__5548\ : Sp12to4
    port map (
            O => \N__30986\,
            I => \N__30969\
        );

    \I__5547\ : InMux
    port map (
            O => \N__30983\,
            I => \N__30966\
        );

    \I__5546\ : LocalMux
    port map (
            O => \N__30980\,
            I => \N__30959\
        );

    \I__5545\ : LocalMux
    port map (
            O => \N__30977\,
            I => \N__30959\
        );

    \I__5544\ : LocalMux
    port map (
            O => \N__30972\,
            I => \N__30959\
        );

    \I__5543\ : Span12Mux_v
    port map (
            O => \N__30969\,
            I => \N__30956\
        );

    \I__5542\ : LocalMux
    port map (
            O => \N__30966\,
            I => \N__30953\
        );

    \I__5541\ : Span4Mux_h
    port map (
            O => \N__30959\,
            I => \N__30950\
        );

    \I__5540\ : Odrv12
    port map (
            O => \N__30956\,
            I => n14490
        );

    \I__5539\ : Odrv4
    port map (
            O => \N__30953\,
            I => n14490
        );

    \I__5538\ : Odrv4
    port map (
            O => \N__30950\,
            I => n14490
        );

    \I__5537\ : InMux
    port map (
            O => \N__30943\,
            I => \N__30940\
        );

    \I__5536\ : LocalMux
    port map (
            O => \N__30940\,
            I => \N__30936\
        );

    \I__5535\ : InMux
    port map (
            O => \N__30939\,
            I => \N__30933\
        );

    \I__5534\ : Span4Mux_h
    port map (
            O => \N__30936\,
            I => \N__30925\
        );

    \I__5533\ : LocalMux
    port map (
            O => \N__30933\,
            I => \N__30922\
        );

    \I__5532\ : InMux
    port map (
            O => \N__30932\,
            I => \N__30917\
        );

    \I__5531\ : InMux
    port map (
            O => \N__30931\,
            I => \N__30917\
        );

    \I__5530\ : InMux
    port map (
            O => \N__30930\,
            I => \N__30912\
        );

    \I__5529\ : InMux
    port map (
            O => \N__30929\,
            I => \N__30912\
        );

    \I__5528\ : InMux
    port map (
            O => \N__30928\,
            I => \N__30909\
        );

    \I__5527\ : Odrv4
    port map (
            O => \N__30925\,
            I => n11882
        );

    \I__5526\ : Odrv4
    port map (
            O => \N__30922\,
            I => n11882
        );

    \I__5525\ : LocalMux
    port map (
            O => \N__30917\,
            I => n11882
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__30912\,
            I => n11882
        );

    \I__5523\ : LocalMux
    port map (
            O => \N__30909\,
            I => n11882
        );

    \I__5522\ : InMux
    port map (
            O => \N__30898\,
            I => \N__30895\
        );

    \I__5521\ : LocalMux
    port map (
            O => \N__30895\,
            I => \N__30892\
        );

    \I__5520\ : Span4Mux_v
    port map (
            O => \N__30892\,
            I => \N__30889\
        );

    \I__5519\ : Span4Mux_h
    port map (
            O => \N__30889\,
            I => \N__30886\
        );

    \I__5518\ : Odrv4
    port map (
            O => \N__30886\,
            I => buf_data_iac_0
        );

    \I__5517\ : InMux
    port map (
            O => \N__30883\,
            I => \N__30880\
        );

    \I__5516\ : LocalMux
    port map (
            O => \N__30880\,
            I => \N__30877\
        );

    \I__5515\ : Span4Mux_v
    port map (
            O => \N__30877\,
            I => \N__30874\
        );

    \I__5514\ : Odrv4
    port map (
            O => \N__30874\,
            I => n22_adj_1476
        );

    \I__5513\ : InMux
    port map (
            O => \N__30871\,
            I => \N__30868\
        );

    \I__5512\ : LocalMux
    port map (
            O => \N__30868\,
            I => \N__30865\
        );

    \I__5511\ : Span4Mux_h
    port map (
            O => \N__30865\,
            I => \N__30862\
        );

    \I__5510\ : Span4Mux_v
    port map (
            O => \N__30862\,
            I => \N__30859\
        );

    \I__5509\ : Span4Mux_v
    port map (
            O => \N__30859\,
            I => \N__30856\
        );

    \I__5508\ : Span4Mux_h
    port map (
            O => \N__30856\,
            I => \N__30853\
        );

    \I__5507\ : Odrv4
    port map (
            O => \N__30853\,
            I => buf_data_vac_8
        );

    \I__5506\ : InMux
    port map (
            O => \N__30850\,
            I => \N__30847\
        );

    \I__5505\ : LocalMux
    port map (
            O => \N__30847\,
            I => \N__30844\
        );

    \I__5504\ : Span4Mux_h
    port map (
            O => \N__30844\,
            I => \N__30841\
        );

    \I__5503\ : Span4Mux_h
    port map (
            O => \N__30841\,
            I => \N__30838\
        );

    \I__5502\ : Span4Mux_h
    port map (
            O => \N__30838\,
            I => \N__30835\
        );

    \I__5501\ : Odrv4
    port map (
            O => \N__30835\,
            I => buf_data_vac_15
        );

    \I__5500\ : InMux
    port map (
            O => \N__30832\,
            I => \N__30829\
        );

    \I__5499\ : LocalMux
    port map (
            O => \N__30829\,
            I => \N__30826\
        );

    \I__5498\ : Span4Mux_v
    port map (
            O => \N__30826\,
            I => \N__30823\
        );

    \I__5497\ : Span4Mux_h
    port map (
            O => \N__30823\,
            I => \N__30820\
        );

    \I__5496\ : Span4Mux_h
    port map (
            O => \N__30820\,
            I => \N__30817\
        );

    \I__5495\ : Odrv4
    port map (
            O => \N__30817\,
            I => buf_data_vac_14
        );

    \I__5494\ : InMux
    port map (
            O => \N__30814\,
            I => \N__30811\
        );

    \I__5493\ : LocalMux
    port map (
            O => \N__30811\,
            I => \N__30807\
        );

    \I__5492\ : InMux
    port map (
            O => \N__30810\,
            I => \N__30804\
        );

    \I__5491\ : Span4Mux_v
    port map (
            O => \N__30807\,
            I => \N__30800\
        );

    \I__5490\ : LocalMux
    port map (
            O => \N__30804\,
            I => \N__30797\
        );

    \I__5489\ : InMux
    port map (
            O => \N__30803\,
            I => \N__30794\
        );

    \I__5488\ : Span4Mux_h
    port map (
            O => \N__30800\,
            I => \N__30791\
        );

    \I__5487\ : Span4Mux_h
    port map (
            O => \N__30797\,
            I => \N__30788\
        );

    \I__5486\ : LocalMux
    port map (
            O => \N__30794\,
            I => \N__30785\
        );

    \I__5485\ : Odrv4
    port map (
            O => \N__30791\,
            I => comm_buf_0_7
        );

    \I__5484\ : Odrv4
    port map (
            O => \N__30788\,
            I => comm_buf_0_7
        );

    \I__5483\ : Odrv4
    port map (
            O => \N__30785\,
            I => comm_buf_0_7
        );

    \I__5482\ : InMux
    port map (
            O => \N__30778\,
            I => \N__30775\
        );

    \I__5481\ : LocalMux
    port map (
            O => \N__30775\,
            I => \ADC_VDC.n10\
        );

    \I__5480\ : InMux
    port map (
            O => \N__30772\,
            I => \N__30767\
        );

    \I__5479\ : InMux
    port map (
            O => \N__30771\,
            I => \N__30764\
        );

    \I__5478\ : InMux
    port map (
            O => \N__30770\,
            I => \N__30761\
        );

    \I__5477\ : LocalMux
    port map (
            O => \N__30767\,
            I => \ADC_VDC.n15\
        );

    \I__5476\ : LocalMux
    port map (
            O => \N__30764\,
            I => \ADC_VDC.n15\
        );

    \I__5475\ : LocalMux
    port map (
            O => \N__30761\,
            I => \ADC_VDC.n15\
        );

    \I__5474\ : InMux
    port map (
            O => \N__30754\,
            I => \N__30751\
        );

    \I__5473\ : LocalMux
    port map (
            O => \N__30751\,
            I => \N__30748\
        );

    \I__5472\ : Odrv4
    port map (
            O => \N__30748\,
            I => \ADC_VDC.n19_adj_1405\
        );

    \I__5471\ : CascadeMux
    port map (
            O => \N__30745\,
            I => \N__30741\
        );

    \I__5470\ : InMux
    port map (
            O => \N__30744\,
            I => \N__30736\
        );

    \I__5469\ : InMux
    port map (
            O => \N__30741\,
            I => \N__30729\
        );

    \I__5468\ : InMux
    port map (
            O => \N__30740\,
            I => \N__30729\
        );

    \I__5467\ : InMux
    port map (
            O => \N__30739\,
            I => \N__30729\
        );

    \I__5466\ : LocalMux
    port map (
            O => \N__30736\,
            I => wdtick_cnt_0
        );

    \I__5465\ : LocalMux
    port map (
            O => \N__30729\,
            I => wdtick_cnt_0
        );

    \I__5464\ : InMux
    port map (
            O => \N__30724\,
            I => \N__30718\
        );

    \I__5463\ : InMux
    port map (
            O => \N__30723\,
            I => \N__30711\
        );

    \I__5462\ : InMux
    port map (
            O => \N__30722\,
            I => \N__30711\
        );

    \I__5461\ : InMux
    port map (
            O => \N__30721\,
            I => \N__30711\
        );

    \I__5460\ : LocalMux
    port map (
            O => \N__30718\,
            I => wdtick_cnt_1
        );

    \I__5459\ : LocalMux
    port map (
            O => \N__30711\,
            I => wdtick_cnt_1
        );

    \I__5458\ : CascadeMux
    port map (
            O => \N__30706\,
            I => \N__30703\
        );

    \I__5457\ : InMux
    port map (
            O => \N__30703\,
            I => \N__30698\
        );

    \I__5456\ : InMux
    port map (
            O => \N__30702\,
            I => \N__30693\
        );

    \I__5455\ : InMux
    port map (
            O => \N__30701\,
            I => \N__30693\
        );

    \I__5454\ : LocalMux
    port map (
            O => \N__30698\,
            I => wdtick_cnt_2
        );

    \I__5453\ : LocalMux
    port map (
            O => \N__30693\,
            I => wdtick_cnt_2
        );

    \I__5452\ : CascadeMux
    port map (
            O => \N__30688\,
            I => \ADC_VDC.n20490_cascade_\
        );

    \I__5451\ : CascadeMux
    port map (
            O => \N__30685\,
            I => \ADC_VDC.n11251_cascade_\
        );

    \I__5450\ : CascadeMux
    port map (
            O => \N__30682\,
            I => \ADC_VDC.n20523_cascade_\
        );

    \I__5449\ : InMux
    port map (
            O => \N__30679\,
            I => \N__30676\
        );

    \I__5448\ : LocalMux
    port map (
            O => \N__30676\,
            I => \N__30673\
        );

    \I__5447\ : Span4Mux_h
    port map (
            O => \N__30673\,
            I => \N__30670\
        );

    \I__5446\ : Odrv4
    port map (
            O => \N__30670\,
            I => \ADC_VDC.n21178\
        );

    \I__5445\ : InMux
    port map (
            O => \N__30667\,
            I => \N__30664\
        );

    \I__5444\ : LocalMux
    port map (
            O => \N__30664\,
            I => \N__30660\
        );

    \I__5443\ : InMux
    port map (
            O => \N__30663\,
            I => \N__30657\
        );

    \I__5442\ : Span4Mux_h
    port map (
            O => \N__30660\,
            I => \N__30654\
        );

    \I__5441\ : LocalMux
    port map (
            O => \N__30657\,
            I => \ADC_VDC.n20490\
        );

    \I__5440\ : Odrv4
    port map (
            O => \N__30654\,
            I => \ADC_VDC.n20490\
        );

    \I__5439\ : InMux
    port map (
            O => \N__30649\,
            I => \N__30646\
        );

    \I__5438\ : LocalMux
    port map (
            O => \N__30646\,
            I => \N__30643\
        );

    \I__5437\ : Span4Mux_h
    port map (
            O => \N__30643\,
            I => \N__30640\
        );

    \I__5436\ : Odrv4
    port map (
            O => \N__30640\,
            I => \ADC_VDC.n21025\
        );

    \I__5435\ : InMux
    port map (
            O => \N__30637\,
            I => \N__30633\
        );

    \I__5434\ : InMux
    port map (
            O => \N__30636\,
            I => \N__30630\
        );

    \I__5433\ : LocalMux
    port map (
            O => \N__30633\,
            I => \ADC_VDC.n7_adj_1403\
        );

    \I__5432\ : LocalMux
    port map (
            O => \N__30630\,
            I => \ADC_VDC.n7_adj_1403\
        );

    \I__5431\ : InMux
    port map (
            O => \N__30625\,
            I => \N__30616\
        );

    \I__5430\ : InMux
    port map (
            O => \N__30624\,
            I => \N__30616\
        );

    \I__5429\ : InMux
    port map (
            O => \N__30623\,
            I => \N__30616\
        );

    \I__5428\ : LocalMux
    port map (
            O => \N__30616\,
            I => \ADC_VDC.n20712\
        );

    \I__5427\ : InMux
    port map (
            O => \N__30613\,
            I => \N__30610\
        );

    \I__5426\ : LocalMux
    port map (
            O => \N__30610\,
            I => \N__30607\
        );

    \I__5425\ : Span4Mux_v
    port map (
            O => \N__30607\,
            I => \N__30604\
        );

    \I__5424\ : Odrv4
    port map (
            O => \N__30604\,
            I => \ADC_VDC.n11662\
        );

    \I__5423\ : InMux
    port map (
            O => \N__30601\,
            I => \N__30598\
        );

    \I__5422\ : LocalMux
    port map (
            O => \N__30598\,
            I => \ADC_VDC.n21028\
        );

    \I__5421\ : InMux
    port map (
            O => \N__30595\,
            I => \N__30591\
        );

    \I__5420\ : InMux
    port map (
            O => \N__30594\,
            I => \N__30588\
        );

    \I__5419\ : LocalMux
    port map (
            O => \N__30591\,
            I => \ADC_VDC.genclk.t0off_14\
        );

    \I__5418\ : LocalMux
    port map (
            O => \N__30588\,
            I => \ADC_VDC.genclk.t0off_14\
        );

    \I__5417\ : CascadeMux
    port map (
            O => \N__30583\,
            I => \N__30580\
        );

    \I__5416\ : InMux
    port map (
            O => \N__30580\,
            I => \N__30576\
        );

    \I__5415\ : InMux
    port map (
            O => \N__30579\,
            I => \N__30573\
        );

    \I__5414\ : LocalMux
    port map (
            O => \N__30576\,
            I => \ADC_VDC.genclk.t0off_9\
        );

    \I__5413\ : LocalMux
    port map (
            O => \N__30573\,
            I => \ADC_VDC.genclk.t0off_9\
        );

    \I__5412\ : CascadeMux
    port map (
            O => \N__30568\,
            I => \N__30564\
        );

    \I__5411\ : InMux
    port map (
            O => \N__30567\,
            I => \N__30561\
        );

    \I__5410\ : InMux
    port map (
            O => \N__30564\,
            I => \N__30558\
        );

    \I__5409\ : LocalMux
    port map (
            O => \N__30561\,
            I => \ADC_VDC.genclk.t0off_15\
        );

    \I__5408\ : LocalMux
    port map (
            O => \N__30558\,
            I => \ADC_VDC.genclk.t0off_15\
        );

    \I__5407\ : CascadeMux
    port map (
            O => \N__30553\,
            I => \N__30550\
        );

    \I__5406\ : InMux
    port map (
            O => \N__30550\,
            I => \N__30546\
        );

    \I__5405\ : InMux
    port map (
            O => \N__30549\,
            I => \N__30543\
        );

    \I__5404\ : LocalMux
    port map (
            O => \N__30546\,
            I => \ADC_VDC.genclk.t0off_11\
        );

    \I__5403\ : LocalMux
    port map (
            O => \N__30543\,
            I => \ADC_VDC.genclk.t0off_11\
        );

    \I__5402\ : InMux
    port map (
            O => \N__30538\,
            I => \N__30535\
        );

    \I__5401\ : LocalMux
    port map (
            O => \N__30535\,
            I => \ADC_VDC.genclk.n28\
        );

    \I__5400\ : CEMux
    port map (
            O => \N__30532\,
            I => \N__30529\
        );

    \I__5399\ : LocalMux
    port map (
            O => \N__30529\,
            I => \N__30525\
        );

    \I__5398\ : CEMux
    port map (
            O => \N__30528\,
            I => \N__30522\
        );

    \I__5397\ : Span4Mux_h
    port map (
            O => \N__30525\,
            I => \N__30519\
        );

    \I__5396\ : LocalMux
    port map (
            O => \N__30522\,
            I => \N__30516\
        );

    \I__5395\ : Odrv4
    port map (
            O => \N__30519\,
            I => \ADC_VDC.genclk.n11721\
        );

    \I__5394\ : Odrv4
    port map (
            O => \N__30516\,
            I => \ADC_VDC.genclk.n11721\
        );

    \I__5393\ : CascadeMux
    port map (
            O => \N__30511\,
            I => \ADC_VDC.n10112_cascade_\
        );

    \I__5392\ : CEMux
    port map (
            O => \N__30508\,
            I => \N__30505\
        );

    \I__5391\ : LocalMux
    port map (
            O => \N__30505\,
            I => \N__30502\
        );

    \I__5390\ : Odrv4
    port map (
            O => \N__30502\,
            I => \ADC_VDC.n12793\
        );

    \I__5389\ : CEMux
    port map (
            O => \N__30499\,
            I => \N__30496\
        );

    \I__5388\ : LocalMux
    port map (
            O => \N__30496\,
            I => \ADC_VDC.n17\
        );

    \I__5387\ : SRMux
    port map (
            O => \N__30493\,
            I => \N__30490\
        );

    \I__5386\ : LocalMux
    port map (
            O => \N__30490\,
            I => \N__30487\
        );

    \I__5385\ : Span4Mux_h
    port map (
            O => \N__30487\,
            I => \N__30484\
        );

    \I__5384\ : Odrv4
    port map (
            O => \N__30484\,
            I => \ADC_VDC.n4\
        );

    \I__5383\ : InMux
    port map (
            O => \N__30481\,
            I => \N__30478\
        );

    \I__5382\ : LocalMux
    port map (
            O => \N__30478\,
            I => \ADC_VDC.n12\
        );

    \I__5381\ : InMux
    port map (
            O => \N__30475\,
            I => \N__30472\
        );

    \I__5380\ : LocalMux
    port map (
            O => \N__30472\,
            I => \ADC_VDC.n72\
        );

    \I__5379\ : InMux
    port map (
            O => \N__30469\,
            I => \N__30466\
        );

    \I__5378\ : LocalMux
    port map (
            O => \N__30466\,
            I => \ADC_VDC.n20710\
        );

    \I__5377\ : CascadeMux
    port map (
            O => \N__30463\,
            I => \N__30458\
        );

    \I__5376\ : CascadeMux
    port map (
            O => \N__30462\,
            I => \N__30455\
        );

    \I__5375\ : InMux
    port map (
            O => \N__30461\,
            I => \N__30451\
        );

    \I__5374\ : InMux
    port map (
            O => \N__30458\,
            I => \N__30448\
        );

    \I__5373\ : InMux
    port map (
            O => \N__30455\,
            I => \N__30443\
        );

    \I__5372\ : InMux
    port map (
            O => \N__30454\,
            I => \N__30443\
        );

    \I__5371\ : LocalMux
    port map (
            O => \N__30451\,
            I => \N__30439\
        );

    \I__5370\ : LocalMux
    port map (
            O => \N__30448\,
            I => \N__30436\
        );

    \I__5369\ : LocalMux
    port map (
            O => \N__30443\,
            I => \N__30433\
        );

    \I__5368\ : InMux
    port map (
            O => \N__30442\,
            I => \N__30430\
        );

    \I__5367\ : Span4Mux_v
    port map (
            O => \N__30439\,
            I => \N__30427\
        );

    \I__5366\ : Span4Mux_v
    port map (
            O => \N__30436\,
            I => \N__30422\
        );

    \I__5365\ : Span4Mux_h
    port map (
            O => \N__30433\,
            I => \N__30422\
        );

    \I__5364\ : LocalMux
    port map (
            O => \N__30430\,
            I => eis_start
        );

    \I__5363\ : Odrv4
    port map (
            O => \N__30427\,
            I => eis_start
        );

    \I__5362\ : Odrv4
    port map (
            O => \N__30422\,
            I => eis_start
        );

    \I__5361\ : InMux
    port map (
            O => \N__30415\,
            I => \N__30412\
        );

    \I__5360\ : LocalMux
    port map (
            O => \N__30412\,
            I => n17357
        );

    \I__5359\ : CascadeMux
    port map (
            O => \N__30409\,
            I => \n11_adj_1620_cascade_\
        );

    \I__5358\ : CEMux
    port map (
            O => \N__30406\,
            I => \N__30403\
        );

    \I__5357\ : LocalMux
    port map (
            O => \N__30403\,
            I => \N__30400\
        );

    \I__5356\ : Span4Mux_v
    port map (
            O => \N__30400\,
            I => \N__30397\
        );

    \I__5355\ : Odrv4
    port map (
            O => \N__30397\,
            I => n11730
        );

    \I__5354\ : CascadeMux
    port map (
            O => \N__30394\,
            I => \N__30391\
        );

    \I__5353\ : InMux
    port map (
            O => \N__30391\,
            I => \N__30387\
        );

    \I__5352\ : InMux
    port map (
            O => \N__30390\,
            I => \N__30384\
        );

    \I__5351\ : LocalMux
    port map (
            O => \N__30387\,
            I => \ADC_VDC.genclk.t0off_6\
        );

    \I__5350\ : LocalMux
    port map (
            O => \N__30384\,
            I => \ADC_VDC.genclk.t0off_6\
        );

    \I__5349\ : InMux
    port map (
            O => \N__30379\,
            I => \N__30375\
        );

    \I__5348\ : InMux
    port map (
            O => \N__30378\,
            I => \N__30372\
        );

    \I__5347\ : LocalMux
    port map (
            O => \N__30375\,
            I => \ADC_VDC.genclk.t0off_1\
        );

    \I__5346\ : LocalMux
    port map (
            O => \N__30372\,
            I => \ADC_VDC.genclk.t0off_1\
        );

    \I__5345\ : CascadeMux
    port map (
            O => \N__30367\,
            I => \N__30363\
        );

    \I__5344\ : CascadeMux
    port map (
            O => \N__30366\,
            I => \N__30360\
        );

    \I__5343\ : InMux
    port map (
            O => \N__30363\,
            I => \N__30357\
        );

    \I__5342\ : InMux
    port map (
            O => \N__30360\,
            I => \N__30354\
        );

    \I__5341\ : LocalMux
    port map (
            O => \N__30357\,
            I => \ADC_VDC.genclk.t0off_4\
        );

    \I__5340\ : LocalMux
    port map (
            O => \N__30354\,
            I => \ADC_VDC.genclk.t0off_4\
        );

    \I__5339\ : InMux
    port map (
            O => \N__30349\,
            I => \N__30345\
        );

    \I__5338\ : InMux
    port map (
            O => \N__30348\,
            I => \N__30342\
        );

    \I__5337\ : LocalMux
    port map (
            O => \N__30345\,
            I => \ADC_VDC.genclk.t0off_0\
        );

    \I__5336\ : LocalMux
    port map (
            O => \N__30342\,
            I => \ADC_VDC.genclk.t0off_0\
        );

    \I__5335\ : CascadeMux
    port map (
            O => \N__30337\,
            I => \ADC_VDC.genclk.n21169_cascade_\
        );

    \I__5334\ : InMux
    port map (
            O => \N__30334\,
            I => \N__30330\
        );

    \I__5333\ : InMux
    port map (
            O => \N__30333\,
            I => \N__30327\
        );

    \I__5332\ : LocalMux
    port map (
            O => \N__30330\,
            I => \ADC_VDC.genclk.t0off_12\
        );

    \I__5331\ : LocalMux
    port map (
            O => \N__30327\,
            I => \ADC_VDC.genclk.t0off_12\
        );

    \I__5330\ : CascadeMux
    port map (
            O => \N__30322\,
            I => \N__30319\
        );

    \I__5329\ : InMux
    port map (
            O => \N__30319\,
            I => \N__30315\
        );

    \I__5328\ : InMux
    port map (
            O => \N__30318\,
            I => \N__30312\
        );

    \I__5327\ : LocalMux
    port map (
            O => \N__30315\,
            I => \ADC_VDC.genclk.t0off_2\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__30312\,
            I => \ADC_VDC.genclk.t0off_2\
        );

    \I__5325\ : CascadeMux
    port map (
            O => \N__30307\,
            I => \N__30303\
        );

    \I__5324\ : InMux
    port map (
            O => \N__30306\,
            I => \N__30300\
        );

    \I__5323\ : InMux
    port map (
            O => \N__30303\,
            I => \N__30297\
        );

    \I__5322\ : LocalMux
    port map (
            O => \N__30300\,
            I => \ADC_VDC.genclk.t0off_7\
        );

    \I__5321\ : LocalMux
    port map (
            O => \N__30297\,
            I => \ADC_VDC.genclk.t0off_7\
        );

    \I__5320\ : InMux
    port map (
            O => \N__30292\,
            I => \N__30288\
        );

    \I__5319\ : InMux
    port map (
            O => \N__30291\,
            I => \N__30285\
        );

    \I__5318\ : LocalMux
    port map (
            O => \N__30288\,
            I => \ADC_VDC.genclk.t0off_10\
        );

    \I__5317\ : LocalMux
    port map (
            O => \N__30285\,
            I => \ADC_VDC.genclk.t0off_10\
        );

    \I__5316\ : InMux
    port map (
            O => \N__30280\,
            I => \N__30277\
        );

    \I__5315\ : LocalMux
    port map (
            O => \N__30277\,
            I => \ADC_VDC.genclk.n27\
        );

    \I__5314\ : CascadeMux
    port map (
            O => \N__30274\,
            I => \N__30271\
        );

    \I__5313\ : InMux
    port map (
            O => \N__30271\,
            I => \N__30267\
        );

    \I__5312\ : InMux
    port map (
            O => \N__30270\,
            I => \N__30264\
        );

    \I__5311\ : LocalMux
    port map (
            O => \N__30267\,
            I => \ADC_VDC.genclk.t0off_13\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__30264\,
            I => \ADC_VDC.genclk.t0off_13\
        );

    \I__5309\ : InMux
    port map (
            O => \N__30259\,
            I => \N__30255\
        );

    \I__5308\ : InMux
    port map (
            O => \N__30258\,
            I => \N__30252\
        );

    \I__5307\ : LocalMux
    port map (
            O => \N__30255\,
            I => \ADC_VDC.genclk.t0off_8\
        );

    \I__5306\ : LocalMux
    port map (
            O => \N__30252\,
            I => \ADC_VDC.genclk.t0off_8\
        );

    \I__5305\ : CascadeMux
    port map (
            O => \N__30247\,
            I => \N__30243\
        );

    \I__5304\ : InMux
    port map (
            O => \N__30246\,
            I => \N__30240\
        );

    \I__5303\ : InMux
    port map (
            O => \N__30243\,
            I => \N__30237\
        );

    \I__5302\ : LocalMux
    port map (
            O => \N__30240\,
            I => \ADC_VDC.genclk.t0off_5\
        );

    \I__5301\ : LocalMux
    port map (
            O => \N__30237\,
            I => \ADC_VDC.genclk.t0off_5\
        );

    \I__5300\ : InMux
    port map (
            O => \N__30232\,
            I => \N__30228\
        );

    \I__5299\ : InMux
    port map (
            O => \N__30231\,
            I => \N__30225\
        );

    \I__5298\ : LocalMux
    port map (
            O => \N__30228\,
            I => \ADC_VDC.genclk.t0off_3\
        );

    \I__5297\ : LocalMux
    port map (
            O => \N__30225\,
            I => \ADC_VDC.genclk.t0off_3\
        );

    \I__5296\ : InMux
    port map (
            O => \N__30220\,
            I => \N__30217\
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__30217\,
            I => \N__30214\
        );

    \I__5294\ : Sp12to4
    port map (
            O => \N__30214\,
            I => \N__30211\
        );

    \I__5293\ : Odrv12
    port map (
            O => \N__30211\,
            I => \ADC_VDC.genclk.n26\
        );

    \I__5292\ : CascadeMux
    port map (
            O => \N__30208\,
            I => \n4_adj_1473_cascade_\
        );

    \I__5291\ : InMux
    port map (
            O => \N__30205\,
            I => \N__30200\
        );

    \I__5290\ : InMux
    port map (
            O => \N__30204\,
            I => \N__30197\
        );

    \I__5289\ : InMux
    port map (
            O => \N__30203\,
            I => \N__30194\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__30200\,
            I => \acadc_skipCount_13\
        );

    \I__5287\ : LocalMux
    port map (
            O => \N__30197\,
            I => \acadc_skipCount_13\
        );

    \I__5286\ : LocalMux
    port map (
            O => \N__30194\,
            I => \acadc_skipCount_13\
        );

    \I__5285\ : InMux
    port map (
            O => \N__30187\,
            I => \N__30182\
        );

    \I__5284\ : InMux
    port map (
            O => \N__30186\,
            I => \N__30179\
        );

    \I__5283\ : InMux
    port map (
            O => \N__30185\,
            I => \N__30176\
        );

    \I__5282\ : LocalMux
    port map (
            O => \N__30182\,
            I => \N__30173\
        );

    \I__5281\ : LocalMux
    port map (
            O => \N__30179\,
            I => \N__30170\
        );

    \I__5280\ : LocalMux
    port map (
            O => \N__30176\,
            I => buf_dds1_10
        );

    \I__5279\ : Odrv4
    port map (
            O => \N__30173\,
            I => buf_dds1_10
        );

    \I__5278\ : Odrv4
    port map (
            O => \N__30170\,
            I => buf_dds1_10
        );

    \I__5277\ : InMux
    port map (
            O => \N__30163\,
            I => \N__30160\
        );

    \I__5276\ : LocalMux
    port map (
            O => \N__30160\,
            I => n22147
        );

    \I__5275\ : InMux
    port map (
            O => \N__30157\,
            I => \N__30154\
        );

    \I__5274\ : LocalMux
    port map (
            O => \N__30154\,
            I => \N__30151\
        );

    \I__5273\ : Span4Mux_v
    port map (
            O => \N__30151\,
            I => \N__30148\
        );

    \I__5272\ : Odrv4
    port map (
            O => \N__30148\,
            I => n22150
        );

    \I__5271\ : CascadeMux
    port map (
            O => \N__30145\,
            I => \n20690_cascade_\
        );

    \I__5270\ : InMux
    port map (
            O => \N__30142\,
            I => \N__30134\
        );

    \I__5269\ : InMux
    port map (
            O => \N__30141\,
            I => \N__30134\
        );

    \I__5268\ : InMux
    port map (
            O => \N__30140\,
            I => \N__30128\
        );

    \I__5267\ : InMux
    port map (
            O => \N__30139\,
            I => \N__30128\
        );

    \I__5266\ : LocalMux
    port map (
            O => \N__30134\,
            I => \N__30125\
        );

    \I__5265\ : InMux
    port map (
            O => \N__30133\,
            I => \N__30122\
        );

    \I__5264\ : LocalMux
    port map (
            O => \N__30128\,
            I => \N__30119\
        );

    \I__5263\ : Span4Mux_h
    port map (
            O => \N__30125\,
            I => \N__30116\
        );

    \I__5262\ : LocalMux
    port map (
            O => \N__30122\,
            I => \N__30111\
        );

    \I__5261\ : Span4Mux_v
    port map (
            O => \N__30119\,
            I => \N__30111\
        );

    \I__5260\ : Odrv4
    port map (
            O => \N__30116\,
            I => acadc_trig
        );

    \I__5259\ : Odrv4
    port map (
            O => \N__30111\,
            I => acadc_trig
        );

    \I__5258\ : InMux
    port map (
            O => \N__30106\,
            I => \N__30103\
        );

    \I__5257\ : LocalMux
    port map (
            O => \N__30103\,
            I => n20529
        );

    \I__5256\ : InMux
    port map (
            O => \N__30100\,
            I => \N__30096\
        );

    \I__5255\ : CascadeMux
    port map (
            O => \N__30099\,
            I => \N__30093\
        );

    \I__5254\ : LocalMux
    port map (
            O => \N__30096\,
            I => \N__30090\
        );

    \I__5253\ : InMux
    port map (
            O => \N__30093\,
            I => \N__30087\
        );

    \I__5252\ : Span4Mux_h
    port map (
            O => \N__30090\,
            I => \N__30084\
        );

    \I__5251\ : LocalMux
    port map (
            O => \N__30087\,
            I => eis_end
        );

    \I__5250\ : Odrv4
    port map (
            O => \N__30084\,
            I => eis_end
        );

    \I__5249\ : InMux
    port map (
            O => \N__30079\,
            I => \N__30075\
        );

    \I__5248\ : InMux
    port map (
            O => \N__30078\,
            I => \N__30072\
        );

    \I__5247\ : LocalMux
    port map (
            O => \N__30075\,
            I => \N__30069\
        );

    \I__5246\ : LocalMux
    port map (
            O => \N__30072\,
            I => \N__30064\
        );

    \I__5245\ : Span4Mux_v
    port map (
            O => \N__30069\,
            I => \N__30064\
        );

    \I__5244\ : Span4Mux_h
    port map (
            O => \N__30064\,
            I => \N__30061\
        );

    \I__5243\ : Odrv4
    port map (
            O => \N__30061\,
            I => n8_adj_1536
        );

    \I__5242\ : IoInMux
    port map (
            O => \N__30058\,
            I => \N__30055\
        );

    \I__5241\ : LocalMux
    port map (
            O => \N__30055\,
            I => \N__30052\
        );

    \I__5240\ : Span4Mux_s2_h
    port map (
            O => \N__30052\,
            I => \N__30049\
        );

    \I__5239\ : Sp12to4
    port map (
            O => \N__30049\,
            I => \N__30046\
        );

    \I__5238\ : Span12Mux_v
    port map (
            O => \N__30046\,
            I => \N__30042\
        );

    \I__5237\ : InMux
    port map (
            O => \N__30045\,
            I => \N__30038\
        );

    \I__5236\ : Span12Mux_h
    port map (
            O => \N__30042\,
            I => \N__30035\
        );

    \I__5235\ : InMux
    port map (
            O => \N__30041\,
            I => \N__30032\
        );

    \I__5234\ : LocalMux
    port map (
            O => \N__30038\,
            I => \N__30029\
        );

    \I__5233\ : Odrv12
    port map (
            O => \N__30035\,
            I => \AMPV_POW\
        );

    \I__5232\ : LocalMux
    port map (
            O => \N__30032\,
            I => \AMPV_POW\
        );

    \I__5231\ : Odrv4
    port map (
            O => \N__30029\,
            I => \AMPV_POW\
        );

    \I__5230\ : InMux
    port map (
            O => \N__30022\,
            I => \N__30018\
        );

    \I__5229\ : InMux
    port map (
            O => \N__30021\,
            I => \N__30015\
        );

    \I__5228\ : LocalMux
    port map (
            O => \N__30018\,
            I => \N__30009\
        );

    \I__5227\ : LocalMux
    port map (
            O => \N__30015\,
            I => \N__30006\
        );

    \I__5226\ : CascadeMux
    port map (
            O => \N__30014\,
            I => \N__30000\
        );

    \I__5225\ : CascadeMux
    port map (
            O => \N__30013\,
            I => \N__29996\
        );

    \I__5224\ : CascadeMux
    port map (
            O => \N__30012\,
            I => \N__29991\
        );

    \I__5223\ : Span4Mux_h
    port map (
            O => \N__30009\,
            I => \N__29987\
        );

    \I__5222\ : Span4Mux_h
    port map (
            O => \N__30006\,
            I => \N__29984\
        );

    \I__5221\ : InMux
    port map (
            O => \N__30005\,
            I => \N__29981\
        );

    \I__5220\ : InMux
    port map (
            O => \N__30004\,
            I => \N__29974\
        );

    \I__5219\ : InMux
    port map (
            O => \N__30003\,
            I => \N__29974\
        );

    \I__5218\ : InMux
    port map (
            O => \N__30000\,
            I => \N__29974\
        );

    \I__5217\ : InMux
    port map (
            O => \N__29999\,
            I => \N__29961\
        );

    \I__5216\ : InMux
    port map (
            O => \N__29996\,
            I => \N__29961\
        );

    \I__5215\ : InMux
    port map (
            O => \N__29995\,
            I => \N__29961\
        );

    \I__5214\ : InMux
    port map (
            O => \N__29994\,
            I => \N__29961\
        );

    \I__5213\ : InMux
    port map (
            O => \N__29991\,
            I => \N__29961\
        );

    \I__5212\ : InMux
    port map (
            O => \N__29990\,
            I => \N__29961\
        );

    \I__5211\ : Odrv4
    port map (
            O => \N__29987\,
            I => \DTRIG_N_910\
        );

    \I__5210\ : Odrv4
    port map (
            O => \N__29984\,
            I => \DTRIG_N_910\
        );

    \I__5209\ : LocalMux
    port map (
            O => \N__29981\,
            I => \DTRIG_N_910\
        );

    \I__5208\ : LocalMux
    port map (
            O => \N__29974\,
            I => \DTRIG_N_910\
        );

    \I__5207\ : LocalMux
    port map (
            O => \N__29961\,
            I => \DTRIG_N_910\
        );

    \I__5206\ : InMux
    port map (
            O => \N__29950\,
            I => \N__29946\
        );

    \I__5205\ : InMux
    port map (
            O => \N__29949\,
            I => \N__29943\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__29946\,
            I => \N__29940\
        );

    \I__5203\ : LocalMux
    port map (
            O => \N__29943\,
            I => \N__29937\
        );

    \I__5202\ : Span4Mux_h
    port map (
            O => \N__29940\,
            I => \N__29924\
        );

    \I__5201\ : Span4Mux_v
    port map (
            O => \N__29937\,
            I => \N__29921\
        );

    \I__5200\ : InMux
    port map (
            O => \N__29936\,
            I => \N__29918\
        );

    \I__5199\ : InMux
    port map (
            O => \N__29935\,
            I => \N__29909\
        );

    \I__5198\ : InMux
    port map (
            O => \N__29934\,
            I => \N__29909\
        );

    \I__5197\ : InMux
    port map (
            O => \N__29933\,
            I => \N__29909\
        );

    \I__5196\ : InMux
    port map (
            O => \N__29932\,
            I => \N__29909\
        );

    \I__5195\ : InMux
    port map (
            O => \N__29931\,
            I => \N__29898\
        );

    \I__5194\ : InMux
    port map (
            O => \N__29930\,
            I => \N__29898\
        );

    \I__5193\ : InMux
    port map (
            O => \N__29929\,
            I => \N__29898\
        );

    \I__5192\ : InMux
    port map (
            O => \N__29928\,
            I => \N__29898\
        );

    \I__5191\ : InMux
    port map (
            O => \N__29927\,
            I => \N__29898\
        );

    \I__5190\ : Odrv4
    port map (
            O => \N__29924\,
            I => adc_state_1
        );

    \I__5189\ : Odrv4
    port map (
            O => \N__29921\,
            I => adc_state_1
        );

    \I__5188\ : LocalMux
    port map (
            O => \N__29918\,
            I => adc_state_1
        );

    \I__5187\ : LocalMux
    port map (
            O => \N__29909\,
            I => adc_state_1
        );

    \I__5186\ : LocalMux
    port map (
            O => \N__29898\,
            I => adc_state_1
        );

    \I__5185\ : InMux
    port map (
            O => \N__29887\,
            I => \N__29883\
        );

    \I__5184\ : InMux
    port map (
            O => \N__29886\,
            I => \N__29880\
        );

    \I__5183\ : LocalMux
    port map (
            O => \N__29883\,
            I => \N__29876\
        );

    \I__5182\ : LocalMux
    port map (
            O => \N__29880\,
            I => \N__29873\
        );

    \I__5181\ : InMux
    port map (
            O => \N__29879\,
            I => \N__29870\
        );

    \I__5180\ : Odrv4
    port map (
            O => \N__29876\,
            I => n10503
        );

    \I__5179\ : Odrv4
    port map (
            O => \N__29873\,
            I => n10503
        );

    \I__5178\ : LocalMux
    port map (
            O => \N__29870\,
            I => n10503
        );

    \I__5177\ : InMux
    port map (
            O => \N__29863\,
            I => \N__29859\
        );

    \I__5176\ : InMux
    port map (
            O => \N__29862\,
            I => \N__29851\
        );

    \I__5175\ : LocalMux
    port map (
            O => \N__29859\,
            I => \N__29848\
        );

    \I__5174\ : CascadeMux
    port map (
            O => \N__29858\,
            I => \N__29842\
        );

    \I__5173\ : CascadeMux
    port map (
            O => \N__29857\,
            I => \N__29838\
        );

    \I__5172\ : InMux
    port map (
            O => \N__29856\,
            I => \N__29830\
        );

    \I__5171\ : InMux
    port map (
            O => \N__29855\,
            I => \N__29830\
        );

    \I__5170\ : InMux
    port map (
            O => \N__29854\,
            I => \N__29830\
        );

    \I__5169\ : LocalMux
    port map (
            O => \N__29851\,
            I => \N__29827\
        );

    \I__5168\ : Span4Mux_v
    port map (
            O => \N__29848\,
            I => \N__29824\
        );

    \I__5167\ : InMux
    port map (
            O => \N__29847\,
            I => \N__29819\
        );

    \I__5166\ : InMux
    port map (
            O => \N__29846\,
            I => \N__29819\
        );

    \I__5165\ : InMux
    port map (
            O => \N__29845\,
            I => \N__29808\
        );

    \I__5164\ : InMux
    port map (
            O => \N__29842\,
            I => \N__29808\
        );

    \I__5163\ : InMux
    port map (
            O => \N__29841\,
            I => \N__29808\
        );

    \I__5162\ : InMux
    port map (
            O => \N__29838\,
            I => \N__29808\
        );

    \I__5161\ : InMux
    port map (
            O => \N__29837\,
            I => \N__29808\
        );

    \I__5160\ : LocalMux
    port map (
            O => \N__29830\,
            I => \N__29805\
        );

    \I__5159\ : Odrv12
    port map (
            O => \N__29827\,
            I => \DTRIG_N_910_adj_1444\
        );

    \I__5158\ : Odrv4
    port map (
            O => \N__29824\,
            I => \DTRIG_N_910_adj_1444\
        );

    \I__5157\ : LocalMux
    port map (
            O => \N__29819\,
            I => \DTRIG_N_910_adj_1444\
        );

    \I__5156\ : LocalMux
    port map (
            O => \N__29808\,
            I => \DTRIG_N_910_adj_1444\
        );

    \I__5155\ : Odrv12
    port map (
            O => \N__29805\,
            I => \DTRIG_N_910_adj_1444\
        );

    \I__5154\ : InMux
    port map (
            O => \N__29794\,
            I => \N__29788\
        );

    \I__5153\ : CascadeMux
    port map (
            O => \N__29793\,
            I => \N__29784\
        );

    \I__5152\ : InMux
    port map (
            O => \N__29792\,
            I => \N__29776\
        );

    \I__5151\ : InMux
    port map (
            O => \N__29791\,
            I => \N__29776\
        );

    \I__5150\ : LocalMux
    port map (
            O => \N__29788\,
            I => \N__29773\
        );

    \I__5149\ : InMux
    port map (
            O => \N__29787\,
            I => \N__29768\
        );

    \I__5148\ : InMux
    port map (
            O => \N__29784\,
            I => \N__29768\
        );

    \I__5147\ : InMux
    port map (
            O => \N__29783\,
            I => \N__29757\
        );

    \I__5146\ : InMux
    port map (
            O => \N__29782\,
            I => \N__29757\
        );

    \I__5145\ : InMux
    port map (
            O => \N__29781\,
            I => \N__29757\
        );

    \I__5144\ : LocalMux
    port map (
            O => \N__29776\,
            I => \N__29754\
        );

    \I__5143\ : Span4Mux_h
    port map (
            O => \N__29773\,
            I => \N__29749\
        );

    \I__5142\ : LocalMux
    port map (
            O => \N__29768\,
            I => \N__29749\
        );

    \I__5141\ : InMux
    port map (
            O => \N__29767\,
            I => \N__29742\
        );

    \I__5140\ : InMux
    port map (
            O => \N__29766\,
            I => \N__29742\
        );

    \I__5139\ : InMux
    port map (
            O => \N__29765\,
            I => \N__29742\
        );

    \I__5138\ : InMux
    port map (
            O => \N__29764\,
            I => \N__29739\
        );

    \I__5137\ : LocalMux
    port map (
            O => \N__29757\,
            I => \N__29736\
        );

    \I__5136\ : Odrv4
    port map (
            O => \N__29754\,
            I => adc_state_1_adj_1410
        );

    \I__5135\ : Odrv4
    port map (
            O => \N__29749\,
            I => adc_state_1_adj_1410
        );

    \I__5134\ : LocalMux
    port map (
            O => \N__29742\,
            I => adc_state_1_adj_1410
        );

    \I__5133\ : LocalMux
    port map (
            O => \N__29739\,
            I => adc_state_1_adj_1410
        );

    \I__5132\ : Odrv4
    port map (
            O => \N__29736\,
            I => adc_state_1_adj_1410
        );

    \I__5131\ : IoInMux
    port map (
            O => \N__29725\,
            I => \N__29722\
        );

    \I__5130\ : LocalMux
    port map (
            O => \N__29722\,
            I => \N__29719\
        );

    \I__5129\ : Span4Mux_s2_h
    port map (
            O => \N__29719\,
            I => \N__29716\
        );

    \I__5128\ : Sp12to4
    port map (
            O => \N__29716\,
            I => \N__29712\
        );

    \I__5127\ : InMux
    port map (
            O => \N__29715\,
            I => \N__29709\
        );

    \I__5126\ : Span12Mux_v
    port map (
            O => \N__29712\,
            I => \N__29706\
        );

    \I__5125\ : LocalMux
    port map (
            O => \N__29709\,
            I => \N__29702\
        );

    \I__5124\ : Span12Mux_h
    port map (
            O => \N__29706\,
            I => \N__29699\
        );

    \I__5123\ : InMux
    port map (
            O => \N__29705\,
            I => \N__29696\
        );

    \I__5122\ : Span4Mux_v
    port map (
            O => \N__29702\,
            I => \N__29693\
        );

    \I__5121\ : Odrv12
    port map (
            O => \N__29699\,
            I => \VAC_OSR1\
        );

    \I__5120\ : LocalMux
    port map (
            O => \N__29696\,
            I => \VAC_OSR1\
        );

    \I__5119\ : Odrv4
    port map (
            O => \N__29693\,
            I => \VAC_OSR1\
        );

    \I__5118\ : CascadeMux
    port map (
            O => \N__29686\,
            I => \n21940_cascade_\
        );

    \I__5117\ : CascadeMux
    port map (
            O => \N__29683\,
            I => \n30_adj_1490_cascade_\
        );

    \I__5116\ : InMux
    port map (
            O => \N__29680\,
            I => \N__29677\
        );

    \I__5115\ : LocalMux
    port map (
            O => \N__29677\,
            I => n26_adj_1495
        );

    \I__5114\ : CascadeMux
    port map (
            O => \N__29674\,
            I => \N__29671\
        );

    \I__5113\ : InMux
    port map (
            O => \N__29671\,
            I => \N__29668\
        );

    \I__5112\ : LocalMux
    port map (
            O => \N__29668\,
            I => \N__29665\
        );

    \I__5111\ : Span4Mux_h
    port map (
            O => \N__29665\,
            I => \N__29662\
        );

    \I__5110\ : Odrv4
    port map (
            O => \N__29662\,
            I => n21109
        );

    \I__5109\ : CascadeMux
    port map (
            O => \N__29659\,
            I => \n22111_cascade_\
        );

    \I__5108\ : InMux
    port map (
            O => \N__29656\,
            I => \N__29653\
        );

    \I__5107\ : LocalMux
    port map (
            O => \N__29653\,
            I => n22114
        );

    \I__5106\ : CascadeMux
    port map (
            O => \N__29650\,
            I => \n16539_cascade_\
        );

    \I__5105\ : CascadeMux
    port map (
            O => \N__29647\,
            I => \n17_adj_1601_cascade_\
        );

    \I__5104\ : InMux
    port map (
            O => \N__29644\,
            I => \N__29641\
        );

    \I__5103\ : LocalMux
    port map (
            O => \N__29641\,
            I => n16547
        );

    \I__5102\ : CascadeMux
    port map (
            O => \N__29638\,
            I => \n16547_cascade_\
        );

    \I__5101\ : CascadeMux
    port map (
            O => \N__29635\,
            I => \n13_cascade_\
        );

    \I__5100\ : InMux
    port map (
            O => \N__29632\,
            I => \N__29629\
        );

    \I__5099\ : LocalMux
    port map (
            O => \N__29629\,
            I => \N__29626\
        );

    \I__5098\ : Span12Mux_h
    port map (
            O => \N__29626\,
            I => \N__29623\
        );

    \I__5097\ : Odrv12
    port map (
            O => \N__29623\,
            I => n19_adj_1482
        );

    \I__5096\ : CascadeMux
    port map (
            O => \N__29620\,
            I => \N__29617\
        );

    \I__5095\ : InMux
    port map (
            O => \N__29617\,
            I => \N__29614\
        );

    \I__5094\ : LocalMux
    port map (
            O => \N__29614\,
            I => \N__29611\
        );

    \I__5093\ : Span4Mux_h
    port map (
            O => \N__29611\,
            I => \N__29608\
        );

    \I__5092\ : Span4Mux_h
    port map (
            O => \N__29608\,
            I => \N__29604\
        );

    \I__5091\ : CascadeMux
    port map (
            O => \N__29607\,
            I => \N__29601\
        );

    \I__5090\ : Span4Mux_v
    port map (
            O => \N__29604\,
            I => \N__29598\
        );

    \I__5089\ : InMux
    port map (
            O => \N__29601\,
            I => \N__29595\
        );

    \I__5088\ : Odrv4
    port map (
            O => \N__29598\,
            I => \buf_readRTD_6\
        );

    \I__5087\ : LocalMux
    port map (
            O => \N__29595\,
            I => \buf_readRTD_6\
        );

    \I__5086\ : CascadeMux
    port map (
            O => \N__29590\,
            I => \n21937_cascade_\
        );

    \I__5085\ : InMux
    port map (
            O => \N__29587\,
            I => \N__29583\
        );

    \I__5084\ : InMux
    port map (
            O => \N__29586\,
            I => \N__29580\
        );

    \I__5083\ : LocalMux
    port map (
            O => \N__29583\,
            I => \N__29577\
        );

    \I__5082\ : LocalMux
    port map (
            O => \N__29580\,
            I => \N__29573\
        );

    \I__5081\ : Span4Mux_h
    port map (
            O => \N__29577\,
            I => \N__29570\
        );

    \I__5080\ : InMux
    port map (
            O => \N__29576\,
            I => \N__29567\
        );

    \I__5079\ : Span4Mux_h
    port map (
            O => \N__29573\,
            I => \N__29562\
        );

    \I__5078\ : Span4Mux_h
    port map (
            O => \N__29570\,
            I => \N__29562\
        );

    \I__5077\ : LocalMux
    port map (
            O => \N__29567\,
            I => buf_adcdata_iac_14
        );

    \I__5076\ : Odrv4
    port map (
            O => \N__29562\,
            I => buf_adcdata_iac_14
        );

    \I__5075\ : InMux
    port map (
            O => \N__29557\,
            I => \N__29552\
        );

    \I__5074\ : InMux
    port map (
            O => \N__29556\,
            I => \N__29549\
        );

    \I__5073\ : InMux
    port map (
            O => \N__29555\,
            I => \N__29546\
        );

    \I__5072\ : LocalMux
    port map (
            O => \N__29552\,
            I => \N__29543\
        );

    \I__5071\ : LocalMux
    port map (
            O => \N__29549\,
            I => buf_dds1_11
        );

    \I__5070\ : LocalMux
    port map (
            O => \N__29546\,
            I => buf_dds1_11
        );

    \I__5069\ : Odrv4
    port map (
            O => \N__29543\,
            I => buf_dds1_11
        );

    \I__5068\ : InMux
    port map (
            O => \N__29536\,
            I => \N__29533\
        );

    \I__5067\ : LocalMux
    port map (
            O => \N__29533\,
            I => \N__29530\
        );

    \I__5066\ : Span12Mux_v
    port map (
            O => \N__29530\,
            I => \N__29527\
        );

    \I__5065\ : Odrv12
    port map (
            O => \N__29527\,
            I => n22075
        );

    \I__5064\ : InMux
    port map (
            O => \N__29524\,
            I => \N__29521\
        );

    \I__5063\ : LocalMux
    port map (
            O => \N__29521\,
            I => \N__29518\
        );

    \I__5062\ : Span4Mux_h
    port map (
            O => \N__29518\,
            I => \N__29515\
        );

    \I__5061\ : Span4Mux_h
    port map (
            O => \N__29515\,
            I => \N__29512\
        );

    \I__5060\ : Odrv4
    port map (
            O => \N__29512\,
            I => n22078
        );

    \I__5059\ : InMux
    port map (
            O => \N__29509\,
            I => \N__29505\
        );

    \I__5058\ : InMux
    port map (
            O => \N__29508\,
            I => \N__29502\
        );

    \I__5057\ : LocalMux
    port map (
            O => \N__29505\,
            I => \N__29499\
        );

    \I__5056\ : LocalMux
    port map (
            O => \N__29502\,
            I => \N__29493\
        );

    \I__5055\ : Span4Mux_v
    port map (
            O => \N__29499\,
            I => \N__29493\
        );

    \I__5054\ : InMux
    port map (
            O => \N__29498\,
            I => \N__29490\
        );

    \I__5053\ : Span4Mux_v
    port map (
            O => \N__29493\,
            I => \N__29487\
        );

    \I__5052\ : LocalMux
    port map (
            O => \N__29490\,
            I => buf_dds1_5
        );

    \I__5051\ : Odrv4
    port map (
            O => \N__29487\,
            I => buf_dds1_5
        );

    \I__5050\ : InMux
    port map (
            O => \N__29482\,
            I => \N__29479\
        );

    \I__5049\ : LocalMux
    port map (
            O => \N__29479\,
            I => n7
        );

    \I__5048\ : InMux
    port map (
            O => \N__29476\,
            I => \N__29459\
        );

    \I__5047\ : InMux
    port map (
            O => \N__29475\,
            I => \N__29459\
        );

    \I__5046\ : InMux
    port map (
            O => \N__29474\,
            I => \N__29459\
        );

    \I__5045\ : InMux
    port map (
            O => \N__29473\,
            I => \N__29459\
        );

    \I__5044\ : InMux
    port map (
            O => \N__29472\,
            I => \N__29459\
        );

    \I__5043\ : InMux
    port map (
            O => \N__29471\,
            I => \N__29454\
        );

    \I__5042\ : InMux
    port map (
            O => \N__29470\,
            I => \N__29454\
        );

    \I__5041\ : LocalMux
    port map (
            O => \N__29459\,
            I => n12214
        );

    \I__5040\ : LocalMux
    port map (
            O => \N__29454\,
            I => n12214
        );

    \I__5039\ : InMux
    port map (
            O => \N__29449\,
            I => \N__29440\
        );

    \I__5038\ : InMux
    port map (
            O => \N__29448\,
            I => \N__29440\
        );

    \I__5037\ : InMux
    port map (
            O => \N__29447\,
            I => \N__29440\
        );

    \I__5036\ : LocalMux
    port map (
            O => \N__29440\,
            I => comm_cmd_4
        );

    \I__5035\ : CascadeMux
    port map (
            O => \N__29437\,
            I => \N__29433\
        );

    \I__5034\ : InMux
    port map (
            O => \N__29436\,
            I => \N__29425\
        );

    \I__5033\ : InMux
    port map (
            O => \N__29433\,
            I => \N__29425\
        );

    \I__5032\ : InMux
    port map (
            O => \N__29432\,
            I => \N__29425\
        );

    \I__5031\ : LocalMux
    port map (
            O => \N__29425\,
            I => comm_cmd_6
        );

    \I__5030\ : InMux
    port map (
            O => \N__29422\,
            I => \N__29417\
        );

    \I__5029\ : InMux
    port map (
            O => \N__29421\,
            I => \N__29412\
        );

    \I__5028\ : InMux
    port map (
            O => \N__29420\,
            I => \N__29412\
        );

    \I__5027\ : LocalMux
    port map (
            O => \N__29417\,
            I => comm_cmd_5
        );

    \I__5026\ : LocalMux
    port map (
            O => \N__29412\,
            I => comm_cmd_5
        );

    \I__5025\ : CascadeMux
    port map (
            O => \N__29407\,
            I => \n8_adj_1522_cascade_\
        );

    \I__5024\ : CascadeMux
    port map (
            O => \N__29404\,
            I => \n12214_cascade_\
        );

    \I__5023\ : InMux
    port map (
            O => \N__29401\,
            I => \N__29398\
        );

    \I__5022\ : LocalMux
    port map (
            O => \N__29398\,
            I => \N__29394\
        );

    \I__5021\ : InMux
    port map (
            O => \N__29397\,
            I => \N__29390\
        );

    \I__5020\ : Span4Mux_v
    port map (
            O => \N__29394\,
            I => \N__29387\
        );

    \I__5019\ : InMux
    port map (
            O => \N__29393\,
            I => \N__29384\
        );

    \I__5018\ : LocalMux
    port map (
            O => \N__29390\,
            I => buf_dds1_13
        );

    \I__5017\ : Odrv4
    port map (
            O => \N__29387\,
            I => buf_dds1_13
        );

    \I__5016\ : LocalMux
    port map (
            O => \N__29384\,
            I => buf_dds1_13
        );

    \I__5015\ : InMux
    port map (
            O => \N__29377\,
            I => \N__29374\
        );

    \I__5014\ : LocalMux
    port map (
            O => \N__29374\,
            I => \N__29371\
        );

    \I__5013\ : Span4Mux_v
    port map (
            O => \N__29371\,
            I => \N__29368\
        );

    \I__5012\ : Span4Mux_h
    port map (
            O => \N__29368\,
            I => \N__29365\
        );

    \I__5011\ : Span4Mux_v
    port map (
            O => \N__29365\,
            I => \N__29362\
        );

    \I__5010\ : Span4Mux_v
    port map (
            O => \N__29362\,
            I => \N__29359\
        );

    \I__5009\ : Odrv4
    port map (
            O => \N__29359\,
            I => \THERMOSTAT\
        );

    \I__5008\ : InMux
    port map (
            O => \N__29356\,
            I => \N__29353\
        );

    \I__5007\ : LocalMux
    port map (
            O => \N__29353\,
            I => \N__29350\
        );

    \I__5006\ : Odrv4
    port map (
            O => \N__29350\,
            I => buf_control_7
        );

    \I__5005\ : CascadeMux
    port map (
            O => \N__29347\,
            I => \n21050_cascade_\
        );

    \I__5004\ : CEMux
    port map (
            O => \N__29344\,
            I => \N__29341\
        );

    \I__5003\ : LocalMux
    port map (
            O => \N__29341\,
            I => \N__29338\
        );

    \I__5002\ : Span4Mux_h
    port map (
            O => \N__29338\,
            I => \N__29335\
        );

    \I__5001\ : Span4Mux_h
    port map (
            O => \N__29335\,
            I => \N__29332\
        );

    \I__5000\ : Odrv4
    port map (
            O => \N__29332\,
            I => n11905
        );

    \I__4999\ : CascadeMux
    port map (
            O => \N__29329\,
            I => \N__29326\
        );

    \I__4998\ : InMux
    port map (
            O => \N__29326\,
            I => \N__29322\
        );

    \I__4997\ : CascadeMux
    port map (
            O => \N__29325\,
            I => \N__29319\
        );

    \I__4996\ : LocalMux
    port map (
            O => \N__29322\,
            I => \N__29314\
        );

    \I__4995\ : InMux
    port map (
            O => \N__29319\,
            I => \N__29311\
        );

    \I__4994\ : CascadeMux
    port map (
            O => \N__29318\,
            I => \N__29308\
        );

    \I__4993\ : InMux
    port map (
            O => \N__29317\,
            I => \N__29305\
        );

    \I__4992\ : Sp12to4
    port map (
            O => \N__29314\,
            I => \N__29300\
        );

    \I__4991\ : LocalMux
    port map (
            O => \N__29311\,
            I => \N__29300\
        );

    \I__4990\ : InMux
    port map (
            O => \N__29308\,
            I => \N__29297\
        );

    \I__4989\ : LocalMux
    port map (
            O => \N__29305\,
            I => \N__29293\
        );

    \I__4988\ : Span12Mux_v
    port map (
            O => \N__29300\,
            I => \N__29288\
        );

    \I__4987\ : LocalMux
    port map (
            O => \N__29297\,
            I => \N__29288\
        );

    \I__4986\ : InMux
    port map (
            O => \N__29296\,
            I => \N__29285\
        );

    \I__4985\ : Span4Mux_v
    port map (
            O => \N__29293\,
            I => \N__29282\
        );

    \I__4984\ : Odrv12
    port map (
            O => \N__29288\,
            I => \buf_cfgRTD_6\
        );

    \I__4983\ : LocalMux
    port map (
            O => \N__29285\,
            I => \buf_cfgRTD_6\
        );

    \I__4982\ : Odrv4
    port map (
            O => \N__29282\,
            I => \buf_cfgRTD_6\
        );

    \I__4981\ : CascadeMux
    port map (
            O => \N__29275\,
            I => \n11882_cascade_\
        );

    \I__4980\ : InMux
    port map (
            O => \N__29272\,
            I => \N__29268\
        );

    \I__4979\ : InMux
    port map (
            O => \N__29271\,
            I => \N__29265\
        );

    \I__4978\ : LocalMux
    port map (
            O => \N__29268\,
            I => \ADC_VDC.avg_cnt_7\
        );

    \I__4977\ : LocalMux
    port map (
            O => \N__29265\,
            I => \ADC_VDC.avg_cnt_7\
        );

    \I__4976\ : InMux
    port map (
            O => \N__29260\,
            I => \ADC_VDC.n19405\
        );

    \I__4975\ : CascadeMux
    port map (
            O => \N__29257\,
            I => \N__29254\
        );

    \I__4974\ : InMux
    port map (
            O => \N__29254\,
            I => \N__29250\
        );

    \I__4973\ : InMux
    port map (
            O => \N__29253\,
            I => \N__29247\
        );

    \I__4972\ : LocalMux
    port map (
            O => \N__29250\,
            I => \N__29244\
        );

    \I__4971\ : LocalMux
    port map (
            O => \N__29247\,
            I => \ADC_VDC.avg_cnt_8\
        );

    \I__4970\ : Odrv12
    port map (
            O => \N__29244\,
            I => \ADC_VDC.avg_cnt_8\
        );

    \I__4969\ : InMux
    port map (
            O => \N__29239\,
            I => \bfn_11_8_0_\
        );

    \I__4968\ : InMux
    port map (
            O => \N__29236\,
            I => \N__29232\
        );

    \I__4967\ : InMux
    port map (
            O => \N__29235\,
            I => \N__29229\
        );

    \I__4966\ : LocalMux
    port map (
            O => \N__29232\,
            I => \ADC_VDC.avg_cnt_9\
        );

    \I__4965\ : LocalMux
    port map (
            O => \N__29229\,
            I => \ADC_VDC.avg_cnt_9\
        );

    \I__4964\ : InMux
    port map (
            O => \N__29224\,
            I => \ADC_VDC.n19407\
        );

    \I__4963\ : InMux
    port map (
            O => \N__29221\,
            I => \N__29217\
        );

    \I__4962\ : InMux
    port map (
            O => \N__29220\,
            I => \N__29214\
        );

    \I__4961\ : LocalMux
    port map (
            O => \N__29217\,
            I => \ADC_VDC.avg_cnt_10\
        );

    \I__4960\ : LocalMux
    port map (
            O => \N__29214\,
            I => \ADC_VDC.avg_cnt_10\
        );

    \I__4959\ : InMux
    port map (
            O => \N__29209\,
            I => \ADC_VDC.n19408\
        );

    \I__4958\ : InMux
    port map (
            O => \N__29206\,
            I => \ADC_VDC.n19409\
        );

    \I__4957\ : InMux
    port map (
            O => \N__29203\,
            I => \N__29199\
        );

    \I__4956\ : InMux
    port map (
            O => \N__29202\,
            I => \N__29196\
        );

    \I__4955\ : LocalMux
    port map (
            O => \N__29199\,
            I => \ADC_VDC.avg_cnt_11\
        );

    \I__4954\ : LocalMux
    port map (
            O => \N__29196\,
            I => \ADC_VDC.avg_cnt_11\
        );

    \I__4953\ : CEMux
    port map (
            O => \N__29191\,
            I => \N__29187\
        );

    \I__4952\ : CEMux
    port map (
            O => \N__29190\,
            I => \N__29183\
        );

    \I__4951\ : LocalMux
    port map (
            O => \N__29187\,
            I => \N__29180\
        );

    \I__4950\ : CEMux
    port map (
            O => \N__29186\,
            I => \N__29174\
        );

    \I__4949\ : LocalMux
    port map (
            O => \N__29183\,
            I => \N__29169\
        );

    \I__4948\ : Span4Mux_v
    port map (
            O => \N__29180\,
            I => \N__29169\
        );

    \I__4947\ : CEMux
    port map (
            O => \N__29179\,
            I => \N__29166\
        );

    \I__4946\ : CEMux
    port map (
            O => \N__29178\,
            I => \N__29163\
        );

    \I__4945\ : CEMux
    port map (
            O => \N__29177\,
            I => \N__29159\
        );

    \I__4944\ : LocalMux
    port map (
            O => \N__29174\,
            I => \N__29152\
        );

    \I__4943\ : Span4Mux_v
    port map (
            O => \N__29169\,
            I => \N__29152\
        );

    \I__4942\ : LocalMux
    port map (
            O => \N__29166\,
            I => \N__29152\
        );

    \I__4941\ : LocalMux
    port map (
            O => \N__29163\,
            I => \N__29149\
        );

    \I__4940\ : CEMux
    port map (
            O => \N__29162\,
            I => \N__29146\
        );

    \I__4939\ : LocalMux
    port map (
            O => \N__29159\,
            I => \N__29143\
        );

    \I__4938\ : Span4Mux_v
    port map (
            O => \N__29152\,
            I => \N__29140\
        );

    \I__4937\ : Span4Mux_v
    port map (
            O => \N__29149\,
            I => \N__29135\
        );

    \I__4936\ : LocalMux
    port map (
            O => \N__29146\,
            I => \N__29135\
        );

    \I__4935\ : Span4Mux_h
    port map (
            O => \N__29143\,
            I => \N__29131\
        );

    \I__4934\ : Span4Mux_h
    port map (
            O => \N__29140\,
            I => \N__29128\
        );

    \I__4933\ : Span4Mux_h
    port map (
            O => \N__29135\,
            I => \N__29125\
        );

    \I__4932\ : InMux
    port map (
            O => \N__29134\,
            I => \N__29122\
        );

    \I__4931\ : Odrv4
    port map (
            O => \N__29131\,
            I => \ADC_VDC.n13060\
        );

    \I__4930\ : Odrv4
    port map (
            O => \N__29128\,
            I => \ADC_VDC.n13060\
        );

    \I__4929\ : Odrv4
    port map (
            O => \N__29125\,
            I => \ADC_VDC.n13060\
        );

    \I__4928\ : LocalMux
    port map (
            O => \N__29122\,
            I => \ADC_VDC.n13060\
        );

    \I__4927\ : SRMux
    port map (
            O => \N__29113\,
            I => \N__29110\
        );

    \I__4926\ : LocalMux
    port map (
            O => \N__29110\,
            I => \N__29105\
        );

    \I__4925\ : SRMux
    port map (
            O => \N__29109\,
            I => \N__29100\
        );

    \I__4924\ : SRMux
    port map (
            O => \N__29108\,
            I => \N__29096\
        );

    \I__4923\ : Span4Mux_v
    port map (
            O => \N__29105\,
            I => \N__29092\
        );

    \I__4922\ : SRMux
    port map (
            O => \N__29104\,
            I => \N__29089\
        );

    \I__4921\ : SRMux
    port map (
            O => \N__29103\,
            I => \N__29086\
        );

    \I__4920\ : LocalMux
    port map (
            O => \N__29100\,
            I => \N__29083\
        );

    \I__4919\ : SRMux
    port map (
            O => \N__29099\,
            I => \N__29080\
        );

    \I__4918\ : LocalMux
    port map (
            O => \N__29096\,
            I => \N__29077\
        );

    \I__4917\ : SRMux
    port map (
            O => \N__29095\,
            I => \N__29074\
        );

    \I__4916\ : Span4Mux_v
    port map (
            O => \N__29092\,
            I => \N__29069\
        );

    \I__4915\ : LocalMux
    port map (
            O => \N__29089\,
            I => \N__29069\
        );

    \I__4914\ : LocalMux
    port map (
            O => \N__29086\,
            I => \N__29066\
        );

    \I__4913\ : Span4Mux_h
    port map (
            O => \N__29083\,
            I => \N__29061\
        );

    \I__4912\ : LocalMux
    port map (
            O => \N__29080\,
            I => \N__29061\
        );

    \I__4911\ : Span4Mux_h
    port map (
            O => \N__29077\,
            I => \N__29056\
        );

    \I__4910\ : LocalMux
    port map (
            O => \N__29074\,
            I => \N__29056\
        );

    \I__4909\ : Span4Mux_v
    port map (
            O => \N__29069\,
            I => \N__29051\
        );

    \I__4908\ : Span4Mux_h
    port map (
            O => \N__29066\,
            I => \N__29051\
        );

    \I__4907\ : Span4Mux_v
    port map (
            O => \N__29061\,
            I => \N__29048\
        );

    \I__4906\ : Span4Mux_v
    port map (
            O => \N__29056\,
            I => \N__29045\
        );

    \I__4905\ : Span4Mux_v
    port map (
            O => \N__29051\,
            I => \N__29042\
        );

    \I__4904\ : Odrv4
    port map (
            O => \N__29048\,
            I => \ADC_VDC.n14900\
        );

    \I__4903\ : Odrv4
    port map (
            O => \N__29045\,
            I => \ADC_VDC.n14900\
        );

    \I__4902\ : Odrv4
    port map (
            O => \N__29042\,
            I => \ADC_VDC.n14900\
        );

    \I__4901\ : CascadeMux
    port map (
            O => \N__29035\,
            I => \n23_adj_1510_cascade_\
        );

    \I__4900\ : InMux
    port map (
            O => \N__29032\,
            I => \N__29029\
        );

    \I__4899\ : LocalMux
    port map (
            O => \N__29029\,
            I => \N__29026\
        );

    \I__4898\ : Span4Mux_v
    port map (
            O => \N__29026\,
            I => \N__29023\
        );

    \I__4897\ : Span4Mux_h
    port map (
            O => \N__29023\,
            I => \N__29020\
        );

    \I__4896\ : Odrv4
    port map (
            O => \N__29020\,
            I => n20833
        );

    \I__4895\ : InMux
    port map (
            O => \N__29017\,
            I => \N__29014\
        );

    \I__4894\ : LocalMux
    port map (
            O => \N__29014\,
            I => \N__29011\
        );

    \I__4893\ : Span4Mux_v
    port map (
            O => \N__29011\,
            I => \N__29008\
        );

    \I__4892\ : Span4Mux_h
    port map (
            O => \N__29008\,
            I => \N__29005\
        );

    \I__4891\ : Span4Mux_h
    port map (
            O => \N__29005\,
            I => \N__29002\
        );

    \I__4890\ : Odrv4
    port map (
            O => \N__29002\,
            I => buf_data_iac_20
        );

    \I__4889\ : CascadeMux
    port map (
            O => \N__28999\,
            I => \N__28996\
        );

    \I__4888\ : InMux
    port map (
            O => \N__28996\,
            I => \N__28993\
        );

    \I__4887\ : LocalMux
    port map (
            O => \N__28993\,
            I => \N__28990\
        );

    \I__4886\ : Span4Mux_h
    port map (
            O => \N__28990\,
            I => \N__28987\
        );

    \I__4885\ : Span4Mux_v
    port map (
            O => \N__28987\,
            I => \N__28984\
        );

    \I__4884\ : Odrv4
    port map (
            O => \N__28984\,
            I => n20810
        );

    \I__4883\ : InMux
    port map (
            O => \N__28981\,
            I => \N__28968\
        );

    \I__4882\ : InMux
    port map (
            O => \N__28980\,
            I => \N__28968\
        );

    \I__4881\ : InMux
    port map (
            O => \N__28979\,
            I => \N__28955\
        );

    \I__4880\ : InMux
    port map (
            O => \N__28978\,
            I => \N__28955\
        );

    \I__4879\ : InMux
    port map (
            O => \N__28977\,
            I => \N__28955\
        );

    \I__4878\ : InMux
    port map (
            O => \N__28976\,
            I => \N__28955\
        );

    \I__4877\ : InMux
    port map (
            O => \N__28975\,
            I => \N__28955\
        );

    \I__4876\ : InMux
    port map (
            O => \N__28974\,
            I => \N__28955\
        );

    \I__4875\ : SRMux
    port map (
            O => \N__28973\,
            I => \N__28944\
        );

    \I__4874\ : LocalMux
    port map (
            O => \N__28968\,
            I => \N__28937\
        );

    \I__4873\ : LocalMux
    port map (
            O => \N__28955\,
            I => \N__28934\
        );

    \I__4872\ : InMux
    port map (
            O => \N__28954\,
            I => \N__28931\
        );

    \I__4871\ : InMux
    port map (
            O => \N__28953\,
            I => \N__28916\
        );

    \I__4870\ : InMux
    port map (
            O => \N__28952\,
            I => \N__28916\
        );

    \I__4869\ : InMux
    port map (
            O => \N__28951\,
            I => \N__28916\
        );

    \I__4868\ : InMux
    port map (
            O => \N__28950\,
            I => \N__28916\
        );

    \I__4867\ : InMux
    port map (
            O => \N__28949\,
            I => \N__28916\
        );

    \I__4866\ : InMux
    port map (
            O => \N__28948\,
            I => \N__28916\
        );

    \I__4865\ : InMux
    port map (
            O => \N__28947\,
            I => \N__28916\
        );

    \I__4864\ : LocalMux
    port map (
            O => \N__28944\,
            I => \N__28913\
        );

    \I__4863\ : InMux
    port map (
            O => \N__28943\,
            I => \N__28910\
        );

    \I__4862\ : CascadeMux
    port map (
            O => \N__28942\,
            I => \N__28904\
        );

    \I__4861\ : InMux
    port map (
            O => \N__28941\,
            I => \N__28899\
        );

    \I__4860\ : InMux
    port map (
            O => \N__28940\,
            I => \N__28899\
        );

    \I__4859\ : Span4Mux_v
    port map (
            O => \N__28937\,
            I => \N__28892\
        );

    \I__4858\ : Span4Mux_v
    port map (
            O => \N__28934\,
            I => \N__28892\
        );

    \I__4857\ : LocalMux
    port map (
            O => \N__28931\,
            I => \N__28892\
        );

    \I__4856\ : LocalMux
    port map (
            O => \N__28916\,
            I => \N__28889\
        );

    \I__4855\ : Span4Mux_h
    port map (
            O => \N__28913\,
            I => \N__28884\
        );

    \I__4854\ : LocalMux
    port map (
            O => \N__28910\,
            I => \N__28884\
        );

    \I__4853\ : InMux
    port map (
            O => \N__28909\,
            I => \N__28881\
        );

    \I__4852\ : CascadeMux
    port map (
            O => \N__28908\,
            I => \N__28877\
        );

    \I__4851\ : CEMux
    port map (
            O => \N__28907\,
            I => \N__28873\
        );

    \I__4850\ : InMux
    port map (
            O => \N__28904\,
            I => \N__28870\
        );

    \I__4849\ : LocalMux
    port map (
            O => \N__28899\,
            I => \N__28867\
        );

    \I__4848\ : Span4Mux_v
    port map (
            O => \N__28892\,
            I => \N__28860\
        );

    \I__4847\ : Span4Mux_v
    port map (
            O => \N__28889\,
            I => \N__28860\
        );

    \I__4846\ : Span4Mux_v
    port map (
            O => \N__28884\,
            I => \N__28855\
        );

    \I__4845\ : LocalMux
    port map (
            O => \N__28881\,
            I => \N__28855\
        );

    \I__4844\ : InMux
    port map (
            O => \N__28880\,
            I => \N__28852\
        );

    \I__4843\ : InMux
    port map (
            O => \N__28877\,
            I => \N__28849\
        );

    \I__4842\ : InMux
    port map (
            O => \N__28876\,
            I => \N__28846\
        );

    \I__4841\ : LocalMux
    port map (
            O => \N__28873\,
            I => \N__28841\
        );

    \I__4840\ : LocalMux
    port map (
            O => \N__28870\,
            I => \N__28841\
        );

    \I__4839\ : Span4Mux_v
    port map (
            O => \N__28867\,
            I => \N__28838\
        );

    \I__4838\ : InMux
    port map (
            O => \N__28866\,
            I => \N__28833\
        );

    \I__4837\ : InMux
    port map (
            O => \N__28865\,
            I => \N__28833\
        );

    \I__4836\ : Span4Mux_v
    port map (
            O => \N__28860\,
            I => \N__28830\
        );

    \I__4835\ : Span4Mux_h
    port map (
            O => \N__28855\,
            I => \N__28827\
        );

    \I__4834\ : LocalMux
    port map (
            O => \N__28852\,
            I => dds_state_1_adj_1446
        );

    \I__4833\ : LocalMux
    port map (
            O => \N__28849\,
            I => dds_state_1_adj_1446
        );

    \I__4832\ : LocalMux
    port map (
            O => \N__28846\,
            I => dds_state_1_adj_1446
        );

    \I__4831\ : Odrv4
    port map (
            O => \N__28841\,
            I => dds_state_1_adj_1446
        );

    \I__4830\ : Odrv4
    port map (
            O => \N__28838\,
            I => dds_state_1_adj_1446
        );

    \I__4829\ : LocalMux
    port map (
            O => \N__28833\,
            I => dds_state_1_adj_1446
        );

    \I__4828\ : Odrv4
    port map (
            O => \N__28830\,
            I => dds_state_1_adj_1446
        );

    \I__4827\ : Odrv4
    port map (
            O => \N__28827\,
            I => dds_state_1_adj_1446
        );

    \I__4826\ : InMux
    port map (
            O => \N__28810\,
            I => \N__28788\
        );

    \I__4825\ : InMux
    port map (
            O => \N__28809\,
            I => \N__28788\
        );

    \I__4824\ : InMux
    port map (
            O => \N__28808\,
            I => \N__28788\
        );

    \I__4823\ : InMux
    port map (
            O => \N__28807\,
            I => \N__28777\
        );

    \I__4822\ : InMux
    port map (
            O => \N__28806\,
            I => \N__28777\
        );

    \I__4821\ : InMux
    port map (
            O => \N__28805\,
            I => \N__28777\
        );

    \I__4820\ : InMux
    port map (
            O => \N__28804\,
            I => \N__28777\
        );

    \I__4819\ : InMux
    port map (
            O => \N__28803\,
            I => \N__28777\
        );

    \I__4818\ : InMux
    port map (
            O => \N__28802\,
            I => \N__28756\
        );

    \I__4817\ : InMux
    port map (
            O => \N__28801\,
            I => \N__28756\
        );

    \I__4816\ : InMux
    port map (
            O => \N__28800\,
            I => \N__28756\
        );

    \I__4815\ : InMux
    port map (
            O => \N__28799\,
            I => \N__28756\
        );

    \I__4814\ : InMux
    port map (
            O => \N__28798\,
            I => \N__28756\
        );

    \I__4813\ : InMux
    port map (
            O => \N__28797\,
            I => \N__28756\
        );

    \I__4812\ : InMux
    port map (
            O => \N__28796\,
            I => \N__28756\
        );

    \I__4811\ : InMux
    port map (
            O => \N__28795\,
            I => \N__28756\
        );

    \I__4810\ : LocalMux
    port map (
            O => \N__28788\,
            I => \N__28751\
        );

    \I__4809\ : LocalMux
    port map (
            O => \N__28777\,
            I => \N__28751\
        );

    \I__4808\ : InMux
    port map (
            O => \N__28776\,
            I => \N__28743\
        );

    \I__4807\ : InMux
    port map (
            O => \N__28775\,
            I => \N__28740\
        );

    \I__4806\ : InMux
    port map (
            O => \N__28774\,
            I => \N__28737\
        );

    \I__4805\ : InMux
    port map (
            O => \N__28773\,
            I => \N__28733\
        );

    \I__4804\ : LocalMux
    port map (
            O => \N__28756\,
            I => \N__28728\
        );

    \I__4803\ : Span4Mux_v
    port map (
            O => \N__28751\,
            I => \N__28728\
        );

    \I__4802\ : InMux
    port map (
            O => \N__28750\,
            I => \N__28725\
        );

    \I__4801\ : InMux
    port map (
            O => \N__28749\,
            I => \N__28716\
        );

    \I__4800\ : InMux
    port map (
            O => \N__28748\,
            I => \N__28716\
        );

    \I__4799\ : InMux
    port map (
            O => \N__28747\,
            I => \N__28716\
        );

    \I__4798\ : InMux
    port map (
            O => \N__28746\,
            I => \N__28716\
        );

    \I__4797\ : LocalMux
    port map (
            O => \N__28743\,
            I => \N__28711\
        );

    \I__4796\ : LocalMux
    port map (
            O => \N__28740\,
            I => \N__28711\
        );

    \I__4795\ : LocalMux
    port map (
            O => \N__28737\,
            I => \N__28708\
        );

    \I__4794\ : InMux
    port map (
            O => \N__28736\,
            I => \N__28705\
        );

    \I__4793\ : LocalMux
    port map (
            O => \N__28733\,
            I => \N__28702\
        );

    \I__4792\ : Span4Mux_v
    port map (
            O => \N__28728\,
            I => \N__28699\
        );

    \I__4791\ : LocalMux
    port map (
            O => \N__28725\,
            I => \N__28694\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__28716\,
            I => \N__28694\
        );

    \I__4789\ : Span4Mux_v
    port map (
            O => \N__28711\,
            I => \N__28689\
        );

    \I__4788\ : Span4Mux_h
    port map (
            O => \N__28708\,
            I => \N__28689\
        );

    \I__4787\ : LocalMux
    port map (
            O => \N__28705\,
            I => dds_state_2_adj_1445
        );

    \I__4786\ : Odrv12
    port map (
            O => \N__28702\,
            I => dds_state_2_adj_1445
        );

    \I__4785\ : Odrv4
    port map (
            O => \N__28699\,
            I => dds_state_2_adj_1445
        );

    \I__4784\ : Odrv4
    port map (
            O => \N__28694\,
            I => dds_state_2_adj_1445
        );

    \I__4783\ : Odrv4
    port map (
            O => \N__28689\,
            I => dds_state_2_adj_1445
        );

    \I__4782\ : CascadeMux
    port map (
            O => \N__28678\,
            I => \N__28674\
        );

    \I__4781\ : CascadeMux
    port map (
            O => \N__28677\,
            I => \N__28671\
        );

    \I__4780\ : InMux
    port map (
            O => \N__28674\,
            I => \N__28668\
        );

    \I__4779\ : InMux
    port map (
            O => \N__28671\,
            I => \N__28665\
        );

    \I__4778\ : LocalMux
    port map (
            O => \N__28668\,
            I => \N__28661\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__28665\,
            I => \N__28658\
        );

    \I__4776\ : CascadeMux
    port map (
            O => \N__28664\,
            I => \N__28655\
        );

    \I__4775\ : Span4Mux_h
    port map (
            O => \N__28661\,
            I => \N__28649\
        );

    \I__4774\ : Span4Mux_v
    port map (
            O => \N__28658\,
            I => \N__28649\
        );

    \I__4773\ : InMux
    port map (
            O => \N__28655\,
            I => \N__28646\
        );

    \I__4772\ : CascadeMux
    port map (
            O => \N__28654\,
            I => \N__28643\
        );

    \I__4771\ : Span4Mux_v
    port map (
            O => \N__28649\,
            I => \N__28640\
        );

    \I__4770\ : LocalMux
    port map (
            O => \N__28646\,
            I => \N__28637\
        );

    \I__4769\ : InMux
    port map (
            O => \N__28643\,
            I => \N__28634\
        );

    \I__4768\ : Span4Mux_v
    port map (
            O => \N__28640\,
            I => \N__28631\
        );

    \I__4767\ : Span12Mux_h
    port map (
            O => \N__28637\,
            I => \N__28628\
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__28634\,
            I => trig_dds1
        );

    \I__4765\ : Odrv4
    port map (
            O => \N__28631\,
            I => trig_dds1
        );

    \I__4764\ : Odrv12
    port map (
            O => \N__28628\,
            I => trig_dds1
        );

    \I__4763\ : InMux
    port map (
            O => \N__28621\,
            I => \N__28618\
        );

    \I__4762\ : LocalMux
    port map (
            O => \N__28618\,
            I => \N__28614\
        );

    \I__4761\ : InMux
    port map (
            O => \N__28617\,
            I => \N__28608\
        );

    \I__4760\ : Span4Mux_h
    port map (
            O => \N__28614\,
            I => \N__28604\
        );

    \I__4759\ : InMux
    port map (
            O => \N__28613\,
            I => \N__28601\
        );

    \I__4758\ : InMux
    port map (
            O => \N__28612\,
            I => \N__28598\
        );

    \I__4757\ : InMux
    port map (
            O => \N__28611\,
            I => \N__28595\
        );

    \I__4756\ : LocalMux
    port map (
            O => \N__28608\,
            I => \N__28588\
        );

    \I__4755\ : InMux
    port map (
            O => \N__28607\,
            I => \N__28585\
        );

    \I__4754\ : Span4Mux_h
    port map (
            O => \N__28604\,
            I => \N__28582\
        );

    \I__4753\ : LocalMux
    port map (
            O => \N__28601\,
            I => \N__28575\
        );

    \I__4752\ : LocalMux
    port map (
            O => \N__28598\,
            I => \N__28575\
        );

    \I__4751\ : LocalMux
    port map (
            O => \N__28595\,
            I => \N__28575\
        );

    \I__4750\ : InMux
    port map (
            O => \N__28594\,
            I => \N__28566\
        );

    \I__4749\ : InMux
    port map (
            O => \N__28593\,
            I => \N__28566\
        );

    \I__4748\ : InMux
    port map (
            O => \N__28592\,
            I => \N__28566\
        );

    \I__4747\ : InMux
    port map (
            O => \N__28591\,
            I => \N__28566\
        );

    \I__4746\ : Odrv4
    port map (
            O => \N__28588\,
            I => dds_state_0_adj_1447
        );

    \I__4745\ : LocalMux
    port map (
            O => \N__28585\,
            I => dds_state_0_adj_1447
        );

    \I__4744\ : Odrv4
    port map (
            O => \N__28582\,
            I => dds_state_0_adj_1447
        );

    \I__4743\ : Odrv4
    port map (
            O => \N__28575\,
            I => dds_state_0_adj_1447
        );

    \I__4742\ : LocalMux
    port map (
            O => \N__28566\,
            I => dds_state_0_adj_1447
        );

    \I__4741\ : CEMux
    port map (
            O => \N__28555\,
            I => \N__28552\
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__28552\,
            I => \N__28548\
        );

    \I__4739\ : CEMux
    port map (
            O => \N__28551\,
            I => \N__28545\
        );

    \I__4738\ : Span4Mux_v
    port map (
            O => \N__28548\,
            I => \N__28540\
        );

    \I__4737\ : LocalMux
    port map (
            O => \N__28545\,
            I => \N__28540\
        );

    \I__4736\ : Span4Mux_v
    port map (
            O => \N__28540\,
            I => \N__28537\
        );

    \I__4735\ : Span4Mux_h
    port map (
            O => \N__28537\,
            I => \N__28534\
        );

    \I__4734\ : Odrv4
    port map (
            O => \N__28534\,
            I => \CLK_DDS.n12722\
        );

    \I__4733\ : InMux
    port map (
            O => \N__28531\,
            I => \N__28527\
        );

    \I__4732\ : InMux
    port map (
            O => \N__28530\,
            I => \N__28524\
        );

    \I__4731\ : LocalMux
    port map (
            O => \N__28527\,
            I => \ADC_VDC.avg_cnt_0\
        );

    \I__4730\ : LocalMux
    port map (
            O => \N__28524\,
            I => \ADC_VDC.avg_cnt_0\
        );

    \I__4729\ : InMux
    port map (
            O => \N__28519\,
            I => \bfn_11_7_0_\
        );

    \I__4728\ : CascadeMux
    port map (
            O => \N__28516\,
            I => \N__28512\
        );

    \I__4727\ : InMux
    port map (
            O => \N__28515\,
            I => \N__28509\
        );

    \I__4726\ : InMux
    port map (
            O => \N__28512\,
            I => \N__28506\
        );

    \I__4725\ : LocalMux
    port map (
            O => \N__28509\,
            I => \ADC_VDC.avg_cnt_1\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__28506\,
            I => \ADC_VDC.avg_cnt_1\
        );

    \I__4723\ : InMux
    port map (
            O => \N__28501\,
            I => \ADC_VDC.n19399\
        );

    \I__4722\ : InMux
    port map (
            O => \N__28498\,
            I => \N__28494\
        );

    \I__4721\ : InMux
    port map (
            O => \N__28497\,
            I => \N__28491\
        );

    \I__4720\ : LocalMux
    port map (
            O => \N__28494\,
            I => \ADC_VDC.avg_cnt_2\
        );

    \I__4719\ : LocalMux
    port map (
            O => \N__28491\,
            I => \ADC_VDC.avg_cnt_2\
        );

    \I__4718\ : InMux
    port map (
            O => \N__28486\,
            I => \ADC_VDC.n19400\
        );

    \I__4717\ : CascadeMux
    port map (
            O => \N__28483\,
            I => \N__28479\
        );

    \I__4716\ : InMux
    port map (
            O => \N__28482\,
            I => \N__28476\
        );

    \I__4715\ : InMux
    port map (
            O => \N__28479\,
            I => \N__28473\
        );

    \I__4714\ : LocalMux
    port map (
            O => \N__28476\,
            I => \ADC_VDC.avg_cnt_3\
        );

    \I__4713\ : LocalMux
    port map (
            O => \N__28473\,
            I => \ADC_VDC.avg_cnt_3\
        );

    \I__4712\ : InMux
    port map (
            O => \N__28468\,
            I => \ADC_VDC.n19401\
        );

    \I__4711\ : InMux
    port map (
            O => \N__28465\,
            I => \N__28461\
        );

    \I__4710\ : InMux
    port map (
            O => \N__28464\,
            I => \N__28458\
        );

    \I__4709\ : LocalMux
    port map (
            O => \N__28461\,
            I => \ADC_VDC.avg_cnt_4\
        );

    \I__4708\ : LocalMux
    port map (
            O => \N__28458\,
            I => \ADC_VDC.avg_cnt_4\
        );

    \I__4707\ : InMux
    port map (
            O => \N__28453\,
            I => \ADC_VDC.n19402\
        );

    \I__4706\ : InMux
    port map (
            O => \N__28450\,
            I => \N__28446\
        );

    \I__4705\ : InMux
    port map (
            O => \N__28449\,
            I => \N__28443\
        );

    \I__4704\ : LocalMux
    port map (
            O => \N__28446\,
            I => \ADC_VDC.avg_cnt_5\
        );

    \I__4703\ : LocalMux
    port map (
            O => \N__28443\,
            I => \ADC_VDC.avg_cnt_5\
        );

    \I__4702\ : InMux
    port map (
            O => \N__28438\,
            I => \ADC_VDC.n19403\
        );

    \I__4701\ : InMux
    port map (
            O => \N__28435\,
            I => \N__28431\
        );

    \I__4700\ : InMux
    port map (
            O => \N__28434\,
            I => \N__28428\
        );

    \I__4699\ : LocalMux
    port map (
            O => \N__28431\,
            I => \ADC_VDC.avg_cnt_6\
        );

    \I__4698\ : LocalMux
    port map (
            O => \N__28428\,
            I => \ADC_VDC.avg_cnt_6\
        );

    \I__4697\ : InMux
    port map (
            O => \N__28423\,
            I => \ADC_VDC.n19404\
        );

    \I__4696\ : InMux
    port map (
            O => \N__28420\,
            I => \N__28399\
        );

    \I__4695\ : InMux
    port map (
            O => \N__28419\,
            I => \N__28399\
        );

    \I__4694\ : InMux
    port map (
            O => \N__28418\,
            I => \N__28399\
        );

    \I__4693\ : InMux
    port map (
            O => \N__28417\,
            I => \N__28399\
        );

    \I__4692\ : InMux
    port map (
            O => \N__28416\,
            I => \N__28399\
        );

    \I__4691\ : InMux
    port map (
            O => \N__28415\,
            I => \N__28399\
        );

    \I__4690\ : InMux
    port map (
            O => \N__28414\,
            I => \N__28399\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__28399\,
            I => \N__28394\
        );

    \I__4688\ : CascadeMux
    port map (
            O => \N__28398\,
            I => \N__28391\
        );

    \I__4687\ : InMux
    port map (
            O => \N__28397\,
            I => \N__28385\
        );

    \I__4686\ : Span4Mux_v
    port map (
            O => \N__28394\,
            I => \N__28382\
        );

    \I__4685\ : InMux
    port map (
            O => \N__28391\,
            I => \N__28373\
        );

    \I__4684\ : InMux
    port map (
            O => \N__28390\,
            I => \N__28373\
        );

    \I__4683\ : InMux
    port map (
            O => \N__28389\,
            I => \N__28373\
        );

    \I__4682\ : InMux
    port map (
            O => \N__28388\,
            I => \N__28373\
        );

    \I__4681\ : LocalMux
    port map (
            O => \N__28385\,
            I => \N__28354\
        );

    \I__4680\ : Span4Mux_h
    port map (
            O => \N__28382\,
            I => \N__28354\
        );

    \I__4679\ : LocalMux
    port map (
            O => \N__28373\,
            I => \N__28354\
        );

    \I__4678\ : InMux
    port map (
            O => \N__28372\,
            I => \N__28337\
        );

    \I__4677\ : InMux
    port map (
            O => \N__28371\,
            I => \N__28337\
        );

    \I__4676\ : InMux
    port map (
            O => \N__28370\,
            I => \N__28337\
        );

    \I__4675\ : InMux
    port map (
            O => \N__28369\,
            I => \N__28337\
        );

    \I__4674\ : InMux
    port map (
            O => \N__28368\,
            I => \N__28337\
        );

    \I__4673\ : InMux
    port map (
            O => \N__28367\,
            I => \N__28337\
        );

    \I__4672\ : InMux
    port map (
            O => \N__28366\,
            I => \N__28337\
        );

    \I__4671\ : InMux
    port map (
            O => \N__28365\,
            I => \N__28337\
        );

    \I__4670\ : InMux
    port map (
            O => \N__28364\,
            I => \N__28330\
        );

    \I__4669\ : InMux
    port map (
            O => \N__28363\,
            I => \N__28330\
        );

    \I__4668\ : InMux
    port map (
            O => \N__28362\,
            I => \N__28330\
        );

    \I__4667\ : InMux
    port map (
            O => \N__28361\,
            I => \N__28327\
        );

    \I__4666\ : Span4Mux_v
    port map (
            O => \N__28354\,
            I => \N__28324\
        );

    \I__4665\ : LocalMux
    port map (
            O => \N__28337\,
            I => \N__28321\
        );

    \I__4664\ : LocalMux
    port map (
            O => \N__28330\,
            I => \N__28318\
        );

    \I__4663\ : LocalMux
    port map (
            O => \N__28327\,
            I => \N__28315\
        );

    \I__4662\ : Span4Mux_h
    port map (
            O => \N__28324\,
            I => \N__28312\
        );

    \I__4661\ : Span4Mux_v
    port map (
            O => \N__28321\,
            I => \N__28307\
        );

    \I__4660\ : Span4Mux_h
    port map (
            O => \N__28318\,
            I => \N__28307\
        );

    \I__4659\ : Odrv12
    port map (
            O => \N__28315\,
            I => n13073
        );

    \I__4658\ : Odrv4
    port map (
            O => \N__28312\,
            I => n13073
        );

    \I__4657\ : Odrv4
    port map (
            O => \N__28307\,
            I => n13073
        );

    \I__4656\ : CascadeMux
    port map (
            O => \N__28300\,
            I => \ADC_VDC.n20618_cascade_\
        );

    \I__4655\ : CEMux
    port map (
            O => \N__28297\,
            I => \N__28294\
        );

    \I__4654\ : LocalMux
    port map (
            O => \N__28294\,
            I => \N__28291\
        );

    \I__4653\ : Span4Mux_v
    port map (
            O => \N__28291\,
            I => \N__28288\
        );

    \I__4652\ : Odrv4
    port map (
            O => \N__28288\,
            I => \ADC_VDC.n47\
        );

    \I__4651\ : InMux
    port map (
            O => \N__28285\,
            I => \N__28282\
        );

    \I__4650\ : LocalMux
    port map (
            O => \N__28282\,
            I => \N__28279\
        );

    \I__4649\ : Odrv4
    port map (
            O => \N__28279\,
            I => \ADC_VDC.n20702\
        );

    \I__4648\ : InMux
    port map (
            O => \N__28276\,
            I => \N__28273\
        );

    \I__4647\ : LocalMux
    port map (
            O => \N__28273\,
            I => \N__28270\
        );

    \I__4646\ : Span4Mux_v
    port map (
            O => \N__28270\,
            I => \N__28267\
        );

    \I__4645\ : Odrv4
    port map (
            O => \N__28267\,
            I => \ADC_VDC.n20\
        );

    \I__4644\ : InMux
    port map (
            O => \N__28264\,
            I => \ADC_VDC.genclk.n19416\
        );

    \I__4643\ : InMux
    port map (
            O => \N__28261\,
            I => \bfn_11_4_0_\
        );

    \I__4642\ : InMux
    port map (
            O => \N__28258\,
            I => \ADC_VDC.genclk.n19418\
        );

    \I__4641\ : InMux
    port map (
            O => \N__28255\,
            I => \ADC_VDC.genclk.n19419\
        );

    \I__4640\ : InMux
    port map (
            O => \N__28252\,
            I => \ADC_VDC.genclk.n19420\
        );

    \I__4639\ : InMux
    port map (
            O => \N__28249\,
            I => \ADC_VDC.genclk.n19421\
        );

    \I__4638\ : InMux
    port map (
            O => \N__28246\,
            I => \ADC_VDC.genclk.n19422\
        );

    \I__4637\ : InMux
    port map (
            O => \N__28243\,
            I => \ADC_VDC.genclk.n19423\
        );

    \I__4636\ : InMux
    port map (
            O => \N__28240\,
            I => \ADC_VDC.genclk.n19424\
        );

    \I__4635\ : InMux
    port map (
            O => \N__28237\,
            I => \N__28234\
        );

    \I__4634\ : LocalMux
    port map (
            O => \N__28234\,
            I => \N__28231\
        );

    \I__4633\ : Span4Mux_h
    port map (
            O => \N__28231\,
            I => \N__28228\
        );

    \I__4632\ : Odrv4
    port map (
            O => \N__28228\,
            I => n16_adj_1489
        );

    \I__4631\ : IoInMux
    port map (
            O => \N__28225\,
            I => \N__28222\
        );

    \I__4630\ : LocalMux
    port map (
            O => \N__28222\,
            I => \N__28219\
        );

    \I__4629\ : IoSpan4Mux
    port map (
            O => \N__28219\,
            I => \N__28216\
        );

    \I__4628\ : Span4Mux_s3_v
    port map (
            O => \N__28216\,
            I => \N__28213\
        );

    \I__4627\ : Span4Mux_v
    port map (
            O => \N__28213\,
            I => \N__28208\
        );

    \I__4626\ : InMux
    port map (
            O => \N__28212\,
            I => \N__28205\
        );

    \I__4625\ : InMux
    port map (
            O => \N__28211\,
            I => \N__28202\
        );

    \I__4624\ : Odrv4
    port map (
            O => \N__28208\,
            I => \IAC_OSR0\
        );

    \I__4623\ : LocalMux
    port map (
            O => \N__28205\,
            I => \IAC_OSR0\
        );

    \I__4622\ : LocalMux
    port map (
            O => \N__28202\,
            I => \IAC_OSR0\
        );

    \I__4621\ : InMux
    port map (
            O => \N__28195\,
            I => \bfn_11_3_0_\
        );

    \I__4620\ : InMux
    port map (
            O => \N__28192\,
            I => \ADC_VDC.genclk.n19410\
        );

    \I__4619\ : InMux
    port map (
            O => \N__28189\,
            I => \ADC_VDC.genclk.n19411\
        );

    \I__4618\ : InMux
    port map (
            O => \N__28186\,
            I => \ADC_VDC.genclk.n19412\
        );

    \I__4617\ : InMux
    port map (
            O => \N__28183\,
            I => \ADC_VDC.genclk.n19413\
        );

    \I__4616\ : InMux
    port map (
            O => \N__28180\,
            I => \ADC_VDC.genclk.n19414\
        );

    \I__4615\ : InMux
    port map (
            O => \N__28177\,
            I => \ADC_VDC.genclk.n19415\
        );

    \I__4614\ : InMux
    port map (
            O => \N__28174\,
            I => \N__28171\
        );

    \I__4613\ : LocalMux
    port map (
            O => \N__28171\,
            I => \N__28168\
        );

    \I__4612\ : Span4Mux_v
    port map (
            O => \N__28168\,
            I => \N__28165\
        );

    \I__4611\ : Odrv4
    port map (
            O => \N__28165\,
            I => n23_adj_1513
        );

    \I__4610\ : CascadeMux
    port map (
            O => \N__28162\,
            I => \N__28158\
        );

    \I__4609\ : CascadeMux
    port map (
            O => \N__28161\,
            I => \N__28154\
        );

    \I__4608\ : InMux
    port map (
            O => \N__28158\,
            I => \N__28151\
        );

    \I__4607\ : InMux
    port map (
            O => \N__28157\,
            I => \N__28146\
        );

    \I__4606\ : InMux
    port map (
            O => \N__28154\,
            I => \N__28146\
        );

    \I__4605\ : LocalMux
    port map (
            O => \N__28151\,
            I => \N__28143\
        );

    \I__4604\ : LocalMux
    port map (
            O => \N__28146\,
            I => cmd_rdadctmp_28
        );

    \I__4603\ : Odrv4
    port map (
            O => \N__28143\,
            I => cmd_rdadctmp_28
        );

    \I__4602\ : InMux
    port map (
            O => \N__28138\,
            I => \N__28135\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__28135\,
            I => \N__28131\
        );

    \I__4600\ : CascadeMux
    port map (
            O => \N__28134\,
            I => \N__28128\
        );

    \I__4599\ : Span4Mux_h
    port map (
            O => \N__28131\,
            I => \N__28125\
        );

    \I__4598\ : InMux
    port map (
            O => \N__28128\,
            I => \N__28122\
        );

    \I__4597\ : Sp12to4
    port map (
            O => \N__28125\,
            I => \N__28118\
        );

    \I__4596\ : LocalMux
    port map (
            O => \N__28122\,
            I => \N__28115\
        );

    \I__4595\ : InMux
    port map (
            O => \N__28121\,
            I => \N__28112\
        );

    \I__4594\ : Span12Mux_v
    port map (
            O => \N__28118\,
            I => \N__28109\
        );

    \I__4593\ : Span4Mux_v
    port map (
            O => \N__28115\,
            I => \N__28106\
        );

    \I__4592\ : LocalMux
    port map (
            O => \N__28112\,
            I => buf_adcdata_iac_20
        );

    \I__4591\ : Odrv12
    port map (
            O => \N__28109\,
            I => buf_adcdata_iac_20
        );

    \I__4590\ : Odrv4
    port map (
            O => \N__28106\,
            I => buf_adcdata_iac_20
        );

    \I__4589\ : IoInMux
    port map (
            O => \N__28099\,
            I => \N__28096\
        );

    \I__4588\ : LocalMux
    port map (
            O => \N__28096\,
            I => \N__28093\
        );

    \I__4587\ : IoSpan4Mux
    port map (
            O => \N__28093\,
            I => \N__28090\
        );

    \I__4586\ : Span4Mux_s0_v
    port map (
            O => \N__28090\,
            I => \N__28087\
        );

    \I__4585\ : Span4Mux_v
    port map (
            O => \N__28087\,
            I => \N__28082\
        );

    \I__4584\ : CascadeMux
    port map (
            O => \N__28086\,
            I => \N__28079\
        );

    \I__4583\ : InMux
    port map (
            O => \N__28085\,
            I => \N__28076\
        );

    \I__4582\ : Span4Mux_v
    port map (
            O => \N__28082\,
            I => \N__28073\
        );

    \I__4581\ : InMux
    port map (
            O => \N__28079\,
            I => \N__28070\
        );

    \I__4580\ : LocalMux
    port map (
            O => \N__28076\,
            I => \N__28067\
        );

    \I__4579\ : Odrv4
    port map (
            O => \N__28073\,
            I => \IAC_FLT1\
        );

    \I__4578\ : LocalMux
    port map (
            O => \N__28070\,
            I => \IAC_FLT1\
        );

    \I__4577\ : Odrv4
    port map (
            O => \N__28067\,
            I => \IAC_FLT1\
        );

    \I__4576\ : IoInMux
    port map (
            O => \N__28060\,
            I => \N__28057\
        );

    \I__4575\ : LocalMux
    port map (
            O => \N__28057\,
            I => \N__28054\
        );

    \I__4574\ : Span4Mux_s1_v
    port map (
            O => \N__28054\,
            I => \N__28051\
        );

    \I__4573\ : Span4Mux_h
    port map (
            O => \N__28051\,
            I => \N__28047\
        );

    \I__4572\ : InMux
    port map (
            O => \N__28050\,
            I => \N__28043\
        );

    \I__4571\ : Span4Mux_v
    port map (
            O => \N__28047\,
            I => \N__28040\
        );

    \I__4570\ : InMux
    port map (
            O => \N__28046\,
            I => \N__28037\
        );

    \I__4569\ : LocalMux
    port map (
            O => \N__28043\,
            I => \N__28034\
        );

    \I__4568\ : Odrv4
    port map (
            O => \N__28040\,
            I => \IAC_OSR1\
        );

    \I__4567\ : LocalMux
    port map (
            O => \N__28037\,
            I => \IAC_OSR1\
        );

    \I__4566\ : Odrv4
    port map (
            O => \N__28034\,
            I => \IAC_OSR1\
        );

    \I__4565\ : IoInMux
    port map (
            O => \N__28027\,
            I => \N__28024\
        );

    \I__4564\ : LocalMux
    port map (
            O => \N__28024\,
            I => \N__28021\
        );

    \I__4563\ : IoSpan4Mux
    port map (
            O => \N__28021\,
            I => \N__28018\
        );

    \I__4562\ : Span4Mux_s1_v
    port map (
            O => \N__28018\,
            I => \N__28015\
        );

    \I__4561\ : Span4Mux_v
    port map (
            O => \N__28015\,
            I => \N__28010\
        );

    \I__4560\ : InMux
    port map (
            O => \N__28014\,
            I => \N__28007\
        );

    \I__4559\ : InMux
    port map (
            O => \N__28013\,
            I => \N__28004\
        );

    \I__4558\ : Odrv4
    port map (
            O => \N__28010\,
            I => \IAC_FLT0\
        );

    \I__4557\ : LocalMux
    port map (
            O => \N__28007\,
            I => \IAC_FLT0\
        );

    \I__4556\ : LocalMux
    port map (
            O => \N__28004\,
            I => \IAC_FLT0\
        );

    \I__4555\ : InMux
    port map (
            O => \N__27997\,
            I => \N__27994\
        );

    \I__4554\ : LocalMux
    port map (
            O => \N__27994\,
            I => \N__27989\
        );

    \I__4553\ : CascadeMux
    port map (
            O => \N__27993\,
            I => \N__27986\
        );

    \I__4552\ : CascadeMux
    port map (
            O => \N__27992\,
            I => \N__27983\
        );

    \I__4551\ : Span4Mux_v
    port map (
            O => \N__27989\,
            I => \N__27980\
        );

    \I__4550\ : InMux
    port map (
            O => \N__27986\,
            I => \N__27977\
        );

    \I__4549\ : InMux
    port map (
            O => \N__27983\,
            I => \N__27974\
        );

    \I__4548\ : Span4Mux_h
    port map (
            O => \N__27980\,
            I => \N__27971\
        );

    \I__4547\ : LocalMux
    port map (
            O => \N__27977\,
            I => buf_adcdata_iac_16
        );

    \I__4546\ : LocalMux
    port map (
            O => \N__27974\,
            I => buf_adcdata_iac_16
        );

    \I__4545\ : Odrv4
    port map (
            O => \N__27971\,
            I => buf_adcdata_iac_16
        );

    \I__4544\ : InMux
    port map (
            O => \N__27964\,
            I => \N__27960\
        );

    \I__4543\ : InMux
    port map (
            O => \N__27963\,
            I => \N__27956\
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__27960\,
            I => \N__27953\
        );

    \I__4541\ : InMux
    port map (
            O => \N__27959\,
            I => \N__27950\
        );

    \I__4540\ : LocalMux
    port map (
            O => \N__27956\,
            I => buf_dds1_8
        );

    \I__4539\ : Odrv12
    port map (
            O => \N__27953\,
            I => buf_dds1_8
        );

    \I__4538\ : LocalMux
    port map (
            O => \N__27950\,
            I => buf_dds1_8
        );

    \I__4537\ : CascadeMux
    port map (
            O => \N__27943\,
            I => \n22189_cascade_\
        );

    \I__4536\ : CascadeMux
    port map (
            O => \N__27940\,
            I => \N__27937\
        );

    \I__4535\ : InMux
    port map (
            O => \N__27937\,
            I => \N__27934\
        );

    \I__4534\ : LocalMux
    port map (
            O => \N__27934\,
            I => \N__27931\
        );

    \I__4533\ : Span4Mux_v
    port map (
            O => \N__27931\,
            I => \N__27928\
        );

    \I__4532\ : Span4Mux_v
    port map (
            O => \N__27928\,
            I => \N__27925\
        );

    \I__4531\ : Odrv4
    port map (
            O => \N__27925\,
            I => n20769
        );

    \I__4530\ : InMux
    port map (
            O => \N__27922\,
            I => \N__27917\
        );

    \I__4529\ : InMux
    port map (
            O => \N__27921\,
            I => \N__27914\
        );

    \I__4528\ : InMux
    port map (
            O => \N__27920\,
            I => \N__27911\
        );

    \I__4527\ : LocalMux
    port map (
            O => \N__27917\,
            I => \N__27908\
        );

    \I__4526\ : LocalMux
    port map (
            O => \N__27914\,
            I => buf_dds1_15
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__27911\,
            I => buf_dds1_15
        );

    \I__4524\ : Odrv4
    port map (
            O => \N__27908\,
            I => buf_dds1_15
        );

    \I__4523\ : InMux
    port map (
            O => \N__27901\,
            I => \N__27898\
        );

    \I__4522\ : LocalMux
    port map (
            O => \N__27898\,
            I => \N__27895\
        );

    \I__4521\ : Odrv4
    port map (
            O => \N__27895\,
            I => n22045
        );

    \I__4520\ : InMux
    port map (
            O => \N__27892\,
            I => \N__27889\
        );

    \I__4519\ : LocalMux
    port map (
            O => \N__27889\,
            I => \N__27886\
        );

    \I__4518\ : Span4Mux_h
    port map (
            O => \N__27886\,
            I => \N__27883\
        );

    \I__4517\ : Odrv4
    port map (
            O => \N__27883\,
            I => n22048
        );

    \I__4516\ : IoInMux
    port map (
            O => \N__27880\,
            I => \N__27877\
        );

    \I__4515\ : LocalMux
    port map (
            O => \N__27877\,
            I => \N__27874\
        );

    \I__4514\ : Span4Mux_s1_h
    port map (
            O => \N__27874\,
            I => \N__27870\
        );

    \I__4513\ : InMux
    port map (
            O => \N__27873\,
            I => \N__27867\
        );

    \I__4512\ : Sp12to4
    port map (
            O => \N__27870\,
            I => \N__27864\
        );

    \I__4511\ : LocalMux
    port map (
            O => \N__27867\,
            I => \N__27861\
        );

    \I__4510\ : Span12Mux_s5_v
    port map (
            O => \N__27864\,
            I => \N__27858\
        );

    \I__4509\ : Span4Mux_v
    port map (
            O => \N__27861\,
            I => \N__27854\
        );

    \I__4508\ : Span12Mux_h
    port map (
            O => \N__27858\,
            I => \N__27851\
        );

    \I__4507\ : InMux
    port map (
            O => \N__27857\,
            I => \N__27848\
        );

    \I__4506\ : Span4Mux_h
    port map (
            O => \N__27854\,
            I => \N__27845\
        );

    \I__4505\ : Odrv12
    port map (
            O => \N__27851\,
            I => \VAC_FLT0\
        );

    \I__4504\ : LocalMux
    port map (
            O => \N__27848\,
            I => \VAC_FLT0\
        );

    \I__4503\ : Odrv4
    port map (
            O => \N__27845\,
            I => \VAC_FLT0\
        );

    \I__4502\ : InMux
    port map (
            O => \N__27838\,
            I => \N__27835\
        );

    \I__4501\ : LocalMux
    port map (
            O => \N__27835\,
            I => \N__27832\
        );

    \I__4500\ : Span4Mux_h
    port map (
            O => \N__27832\,
            I => \N__27829\
        );

    \I__4499\ : Odrv4
    port map (
            O => \N__27829\,
            I => n16_adj_1480
        );

    \I__4498\ : InMux
    port map (
            O => \N__27826\,
            I => \N__27821\
        );

    \I__4497\ : InMux
    port map (
            O => \N__27825\,
            I => \N__27816\
        );

    \I__4496\ : InMux
    port map (
            O => \N__27824\,
            I => \N__27816\
        );

    \I__4495\ : LocalMux
    port map (
            O => \N__27821\,
            I => buf_dds1_0
        );

    \I__4494\ : LocalMux
    port map (
            O => \N__27816\,
            I => buf_dds1_0
        );

    \I__4493\ : InMux
    port map (
            O => \N__27811\,
            I => \N__27808\
        );

    \I__4492\ : LocalMux
    port map (
            O => \N__27808\,
            I => \N__27805\
        );

    \I__4491\ : Span4Mux_h
    port map (
            O => \N__27805\,
            I => \N__27802\
        );

    \I__4490\ : Span4Mux_v
    port map (
            O => \N__27802\,
            I => \N__27797\
        );

    \I__4489\ : CascadeMux
    port map (
            O => \N__27801\,
            I => \N__27794\
        );

    \I__4488\ : InMux
    port map (
            O => \N__27800\,
            I => \N__27791\
        );

    \I__4487\ : Span4Mux_v
    port map (
            O => \N__27797\,
            I => \N__27788\
        );

    \I__4486\ : InMux
    port map (
            O => \N__27794\,
            I => \N__27785\
        );

    \I__4485\ : LocalMux
    port map (
            O => \N__27791\,
            I => buf_adcdata_iac_18
        );

    \I__4484\ : Odrv4
    port map (
            O => \N__27788\,
            I => buf_adcdata_iac_18
        );

    \I__4483\ : LocalMux
    port map (
            O => \N__27785\,
            I => buf_adcdata_iac_18
        );

    \I__4482\ : CascadeMux
    port map (
            O => \N__27778\,
            I => \N__27774\
        );

    \I__4481\ : InMux
    port map (
            O => \N__27777\,
            I => \N__27770\
        );

    \I__4480\ : InMux
    port map (
            O => \N__27774\,
            I => \N__27767\
        );

    \I__4479\ : InMux
    port map (
            O => \N__27773\,
            I => \N__27764\
        );

    \I__4478\ : LocalMux
    port map (
            O => \N__27770\,
            I => cmd_rdadctmp_25
        );

    \I__4477\ : LocalMux
    port map (
            O => \N__27767\,
            I => cmd_rdadctmp_25
        );

    \I__4476\ : LocalMux
    port map (
            O => \N__27764\,
            I => cmd_rdadctmp_25
        );

    \I__4475\ : InMux
    port map (
            O => \N__27757\,
            I => \N__27753\
        );

    \I__4474\ : CascadeMux
    port map (
            O => \N__27756\,
            I => \N__27750\
        );

    \I__4473\ : LocalMux
    port map (
            O => \N__27753\,
            I => \N__27747\
        );

    \I__4472\ : InMux
    port map (
            O => \N__27750\,
            I => \N__27743\
        );

    \I__4471\ : Span4Mux_h
    port map (
            O => \N__27747\,
            I => \N__27740\
        );

    \I__4470\ : InMux
    port map (
            O => \N__27746\,
            I => \N__27737\
        );

    \I__4469\ : LocalMux
    port map (
            O => \N__27743\,
            I => cmd_rdadctmp_26
        );

    \I__4468\ : Odrv4
    port map (
            O => \N__27740\,
            I => cmd_rdadctmp_26
        );

    \I__4467\ : LocalMux
    port map (
            O => \N__27737\,
            I => cmd_rdadctmp_26
        );

    \I__4466\ : CascadeMux
    port map (
            O => \N__27730\,
            I => \N__27727\
        );

    \I__4465\ : InMux
    port map (
            O => \N__27727\,
            I => \N__27723\
        );

    \I__4464\ : InMux
    port map (
            O => \N__27726\,
            I => \N__27720\
        );

    \I__4463\ : LocalMux
    port map (
            O => \N__27723\,
            I => \N__27717\
        );

    \I__4462\ : LocalMux
    port map (
            O => \N__27720\,
            I => \N__27714\
        );

    \I__4461\ : Span4Mux_v
    port map (
            O => \N__27717\,
            I => \N__27709\
        );

    \I__4460\ : Span4Mux_h
    port map (
            O => \N__27714\,
            I => \N__27709\
        );

    \I__4459\ : Odrv4
    port map (
            O => \N__27709\,
            I => tmp_buf_15_adj_1448
        );

    \I__4458\ : CascadeMux
    port map (
            O => \N__27706\,
            I => \N__27703\
        );

    \I__4457\ : InMux
    port map (
            O => \N__27703\,
            I => \N__27700\
        );

    \I__4456\ : LocalMux
    port map (
            O => \N__27700\,
            I => \CLK_DDS.tmp_buf_0\
        );

    \I__4455\ : CascadeMux
    port map (
            O => \N__27697\,
            I => \N__27694\
        );

    \I__4454\ : InMux
    port map (
            O => \N__27694\,
            I => \N__27691\
        );

    \I__4453\ : LocalMux
    port map (
            O => \N__27691\,
            I => \CLK_DDS.tmp_buf_1\
        );

    \I__4452\ : CascadeMux
    port map (
            O => \N__27688\,
            I => \N__27685\
        );

    \I__4451\ : InMux
    port map (
            O => \N__27685\,
            I => \N__27682\
        );

    \I__4450\ : LocalMux
    port map (
            O => \N__27682\,
            I => \CLK_DDS.tmp_buf_2\
        );

    \I__4449\ : CascadeMux
    port map (
            O => \N__27679\,
            I => \N__27676\
        );

    \I__4448\ : InMux
    port map (
            O => \N__27676\,
            I => \N__27673\
        );

    \I__4447\ : LocalMux
    port map (
            O => \N__27673\,
            I => \N__27670\
        );

    \I__4446\ : Odrv4
    port map (
            O => \N__27670\,
            I => \CLK_DDS.tmp_buf_3\
        );

    \I__4445\ : CascadeMux
    port map (
            O => \N__27667\,
            I => \N__27664\
        );

    \I__4444\ : InMux
    port map (
            O => \N__27664\,
            I => \N__27661\
        );

    \I__4443\ : LocalMux
    port map (
            O => \N__27661\,
            I => \CLK_DDS.tmp_buf_4\
        );

    \I__4442\ : CascadeMux
    port map (
            O => \N__27658\,
            I => \N__27655\
        );

    \I__4441\ : InMux
    port map (
            O => \N__27655\,
            I => \N__27652\
        );

    \I__4440\ : LocalMux
    port map (
            O => \N__27652\,
            I => \CLK_DDS.tmp_buf_5\
        );

    \I__4439\ : CascadeMux
    port map (
            O => \N__27649\,
            I => \N__27646\
        );

    \I__4438\ : InMux
    port map (
            O => \N__27646\,
            I => \N__27643\
        );

    \I__4437\ : LocalMux
    port map (
            O => \N__27643\,
            I => \CLK_DDS.tmp_buf_6\
        );

    \I__4436\ : CascadeMux
    port map (
            O => \N__27640\,
            I => \N__27637\
        );

    \I__4435\ : InMux
    port map (
            O => \N__27637\,
            I => \N__27634\
        );

    \I__4434\ : LocalMux
    port map (
            O => \N__27634\,
            I => \N__27631\
        );

    \I__4433\ : Odrv12
    port map (
            O => \N__27631\,
            I => \CLK_DDS.tmp_buf_7\
        );

    \I__4432\ : CascadeMux
    port map (
            O => \N__27628\,
            I => \N__27625\
        );

    \I__4431\ : InMux
    port map (
            O => \N__27625\,
            I => \N__27622\
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__27622\,
            I => \CLK_DDS.tmp_buf_9\
        );

    \I__4429\ : InMux
    port map (
            O => \N__27619\,
            I => \N__27616\
        );

    \I__4428\ : LocalMux
    port map (
            O => \N__27616\,
            I => \CLK_DDS.tmp_buf_8\
        );

    \I__4427\ : InMux
    port map (
            O => \N__27613\,
            I => \N__27610\
        );

    \I__4426\ : LocalMux
    port map (
            O => \N__27610\,
            I => \N__27605\
        );

    \I__4425\ : InMux
    port map (
            O => \N__27609\,
            I => \N__27602\
        );

    \I__4424\ : InMux
    port map (
            O => \N__27608\,
            I => \N__27599\
        );

    \I__4423\ : Span4Mux_v
    port map (
            O => \N__27605\,
            I => \N__27596\
        );

    \I__4422\ : LocalMux
    port map (
            O => \N__27602\,
            I => buf_dds1_14
        );

    \I__4421\ : LocalMux
    port map (
            O => \N__27599\,
            I => buf_dds1_14
        );

    \I__4420\ : Odrv4
    port map (
            O => \N__27596\,
            I => buf_dds1_14
        );

    \I__4419\ : InMux
    port map (
            O => \N__27589\,
            I => \N__27584\
        );

    \I__4418\ : InMux
    port map (
            O => \N__27588\,
            I => \N__27581\
        );

    \I__4417\ : InMux
    port map (
            O => \N__27587\,
            I => \N__27578\
        );

    \I__4416\ : LocalMux
    port map (
            O => \N__27584\,
            I => buf_dds1_12
        );

    \I__4415\ : LocalMux
    port map (
            O => \N__27581\,
            I => buf_dds1_12
        );

    \I__4414\ : LocalMux
    port map (
            O => \N__27578\,
            I => buf_dds1_12
        );

    \I__4413\ : InMux
    port map (
            O => \N__27571\,
            I => \N__27567\
        );

    \I__4412\ : CascadeMux
    port map (
            O => \N__27570\,
            I => \N__27563\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__27567\,
            I => \N__27560\
        );

    \I__4410\ : InMux
    port map (
            O => \N__27566\,
            I => \N__27557\
        );

    \I__4409\ : InMux
    port map (
            O => \N__27563\,
            I => \N__27554\
        );

    \I__4408\ : Span4Mux_h
    port map (
            O => \N__27560\,
            I => \N__27551\
        );

    \I__4407\ : LocalMux
    port map (
            O => \N__27557\,
            I => buf_dds1_9
        );

    \I__4406\ : LocalMux
    port map (
            O => \N__27554\,
            I => buf_dds1_9
        );

    \I__4405\ : Odrv4
    port map (
            O => \N__27551\,
            I => buf_dds1_9
        );

    \I__4404\ : CascadeMux
    port map (
            O => \N__27544\,
            I => \n22036_cascade_\
        );

    \I__4403\ : InMux
    port map (
            O => \N__27541\,
            I => \N__27538\
        );

    \I__4402\ : LocalMux
    port map (
            O => \N__27538\,
            I => \N__27535\
        );

    \I__4401\ : Span4Mux_h
    port map (
            O => \N__27535\,
            I => \N__27532\
        );

    \I__4400\ : Odrv4
    port map (
            O => \N__27532\,
            I => n22156
        );

    \I__4399\ : InMux
    port map (
            O => \N__27529\,
            I => \N__27526\
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__27526\,
            I => n21910
        );

    \I__4397\ : CascadeMux
    port map (
            O => \N__27523\,
            I => \n20823_cascade_\
        );

    \I__4396\ : CascadeMux
    port map (
            O => \N__27520\,
            I => \n30_adj_1514_cascade_\
        );

    \I__4395\ : CEMux
    port map (
            O => \N__27517\,
            I => \N__27514\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__27514\,
            I => \N__27509\
        );

    \I__4393\ : CEMux
    port map (
            O => \N__27513\,
            I => \N__27506\
        );

    \I__4392\ : CEMux
    port map (
            O => \N__27512\,
            I => \N__27501\
        );

    \I__4391\ : Span4Mux_h
    port map (
            O => \N__27509\,
            I => \N__27496\
        );

    \I__4390\ : LocalMux
    port map (
            O => \N__27506\,
            I => \N__27496\
        );

    \I__4389\ : CEMux
    port map (
            O => \N__27505\,
            I => \N__27493\
        );

    \I__4388\ : CEMux
    port map (
            O => \N__27504\,
            I => \N__27490\
        );

    \I__4387\ : LocalMux
    port map (
            O => \N__27501\,
            I => \N__27487\
        );

    \I__4386\ : Span4Mux_h
    port map (
            O => \N__27496\,
            I => \N__27484\
        );

    \I__4385\ : LocalMux
    port map (
            O => \N__27493\,
            I => \N__27481\
        );

    \I__4384\ : LocalMux
    port map (
            O => \N__27490\,
            I => \N__27478\
        );

    \I__4383\ : Odrv4
    port map (
            O => \N__27487\,
            I => n11941
        );

    \I__4382\ : Odrv4
    port map (
            O => \N__27484\,
            I => n11941
        );

    \I__4381\ : Odrv12
    port map (
            O => \N__27481\,
            I => n11941
        );

    \I__4380\ : Odrv12
    port map (
            O => \N__27478\,
            I => n11941
        );

    \I__4379\ : SRMux
    port map (
            O => \N__27469\,
            I => \N__27466\
        );

    \I__4378\ : LocalMux
    port map (
            O => \N__27466\,
            I => \N__27461\
        );

    \I__4377\ : SRMux
    port map (
            O => \N__27465\,
            I => \N__27458\
        );

    \I__4376\ : SRMux
    port map (
            O => \N__27464\,
            I => \N__27455\
        );

    \I__4375\ : Span4Mux_v
    port map (
            O => \N__27461\,
            I => \N__27448\
        );

    \I__4374\ : LocalMux
    port map (
            O => \N__27458\,
            I => \N__27448\
        );

    \I__4373\ : LocalMux
    port map (
            O => \N__27455\,
            I => \N__27445\
        );

    \I__4372\ : SRMux
    port map (
            O => \N__27454\,
            I => \N__27442\
        );

    \I__4371\ : SRMux
    port map (
            O => \N__27453\,
            I => \N__27439\
        );

    \I__4370\ : Span4Mux_h
    port map (
            O => \N__27448\,
            I => \N__27436\
        );

    \I__4369\ : Span4Mux_h
    port map (
            O => \N__27445\,
            I => \N__27433\
        );

    \I__4368\ : LocalMux
    port map (
            O => \N__27442\,
            I => \N__27430\
        );

    \I__4367\ : LocalMux
    port map (
            O => \N__27439\,
            I => \N__27427\
        );

    \I__4366\ : Odrv4
    port map (
            O => \N__27436\,
            I => n14735
        );

    \I__4365\ : Odrv4
    port map (
            O => \N__27433\,
            I => n14735
        );

    \I__4364\ : Odrv12
    port map (
            O => \N__27430\,
            I => n14735
        );

    \I__4363\ : Odrv12
    port map (
            O => \N__27427\,
            I => n14735
        );

    \I__4362\ : CascadeMux
    port map (
            O => \N__27418\,
            I => \N__27415\
        );

    \I__4361\ : InMux
    port map (
            O => \N__27415\,
            I => \N__27412\
        );

    \I__4360\ : LocalMux
    port map (
            O => \N__27412\,
            I => \CLK_DDS.tmp_buf_10\
        );

    \I__4359\ : CascadeMux
    port map (
            O => \N__27409\,
            I => \N__27406\
        );

    \I__4358\ : InMux
    port map (
            O => \N__27406\,
            I => \N__27403\
        );

    \I__4357\ : LocalMux
    port map (
            O => \N__27403\,
            I => \CLK_DDS.tmp_buf_11\
        );

    \I__4356\ : CascadeMux
    port map (
            O => \N__27400\,
            I => \N__27397\
        );

    \I__4355\ : InMux
    port map (
            O => \N__27397\,
            I => \N__27394\
        );

    \I__4354\ : LocalMux
    port map (
            O => \N__27394\,
            I => \CLK_DDS.tmp_buf_12\
        );

    \I__4353\ : CascadeMux
    port map (
            O => \N__27391\,
            I => \N__27388\
        );

    \I__4352\ : InMux
    port map (
            O => \N__27388\,
            I => \N__27385\
        );

    \I__4351\ : LocalMux
    port map (
            O => \N__27385\,
            I => \CLK_DDS.tmp_buf_13\
        );

    \I__4350\ : CascadeMux
    port map (
            O => \N__27382\,
            I => \N__27379\
        );

    \I__4349\ : InMux
    port map (
            O => \N__27379\,
            I => \N__27376\
        );

    \I__4348\ : LocalMux
    port map (
            O => \N__27376\,
            I => \CLK_DDS.tmp_buf_14\
        );

    \I__4347\ : InMux
    port map (
            O => \N__27373\,
            I => \N__27370\
        );

    \I__4346\ : LocalMux
    port map (
            O => \N__27370\,
            I => \N__27367\
        );

    \I__4345\ : Span4Mux_h
    port map (
            O => \N__27367\,
            I => \N__27364\
        );

    \I__4344\ : Span4Mux_h
    port map (
            O => \N__27364\,
            I => \N__27361\
        );

    \I__4343\ : Odrv4
    port map (
            O => \N__27361\,
            I => buf_data_iac_18
        );

    \I__4342\ : CascadeMux
    port map (
            O => \N__27358\,
            I => \n20794_cascade_\
        );

    \I__4341\ : InMux
    port map (
            O => \N__27355\,
            I => \N__27352\
        );

    \I__4340\ : LocalMux
    port map (
            O => \N__27352\,
            I => n21922
        );

    \I__4339\ : CascadeMux
    port map (
            O => \N__27349\,
            I => \n20796_cascade_\
        );

    \I__4338\ : InMux
    port map (
            O => \N__27346\,
            I => \N__27343\
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__27343\,
            I => \N__27340\
        );

    \I__4336\ : Span4Mux_h
    port map (
            O => \N__27340\,
            I => \N__27337\
        );

    \I__4335\ : Odrv4
    port map (
            O => \N__27337\,
            I => n21934
        );

    \I__4334\ : CascadeMux
    port map (
            O => \N__27334\,
            I => \n22213_cascade_\
        );

    \I__4333\ : CascadeMux
    port map (
            O => \N__27331\,
            I => \n22216_cascade_\
        );

    \I__4332\ : InMux
    port map (
            O => \N__27328\,
            I => \N__27325\
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__27325\,
            I => \N__27322\
        );

    \I__4330\ : Span4Mux_h
    port map (
            O => \N__27322\,
            I => \N__27319\
        );

    \I__4329\ : Span4Mux_h
    port map (
            O => \N__27319\,
            I => \N__27316\
        );

    \I__4328\ : Odrv4
    port map (
            O => \N__27316\,
            I => n20937
        );

    \I__4327\ : CascadeMux
    port map (
            O => \N__27313\,
            I => \N__27310\
        );

    \I__4326\ : InMux
    port map (
            O => \N__27310\,
            I => \N__27307\
        );

    \I__4325\ : LocalMux
    port map (
            O => \N__27307\,
            I => n20936
        );

    \I__4324\ : CascadeMux
    port map (
            O => \N__27304\,
            I => \n21907_cascade_\
        );

    \I__4323\ : InMux
    port map (
            O => \N__27301\,
            I => \N__27297\
        );

    \I__4322\ : CascadeMux
    port map (
            O => \N__27300\,
            I => \N__27294\
        );

    \I__4321\ : LocalMux
    port map (
            O => \N__27297\,
            I => \N__27291\
        );

    \I__4320\ : InMux
    port map (
            O => \N__27294\,
            I => \N__27288\
        );

    \I__4319\ : Span12Mux_h
    port map (
            O => \N__27291\,
            I => \N__27284\
        );

    \I__4318\ : LocalMux
    port map (
            O => \N__27288\,
            I => \N__27281\
        );

    \I__4317\ : InMux
    port map (
            O => \N__27287\,
            I => \N__27278\
        );

    \I__4316\ : Span12Mux_v
    port map (
            O => \N__27284\,
            I => \N__27275\
        );

    \I__4315\ : Span4Mux_h
    port map (
            O => \N__27281\,
            I => \N__27272\
        );

    \I__4314\ : LocalMux
    port map (
            O => \N__27278\,
            I => buf_adcdata_iac_21
        );

    \I__4313\ : Odrv12
    port map (
            O => \N__27275\,
            I => buf_adcdata_iac_21
        );

    \I__4312\ : Odrv4
    port map (
            O => \N__27272\,
            I => buf_adcdata_iac_21
        );

    \I__4311\ : CascadeMux
    port map (
            O => \N__27265\,
            I => \n22033_cascade_\
        );

    \I__4310\ : CascadeMux
    port map (
            O => \N__27262\,
            I => \n12_cascade_\
        );

    \I__4309\ : CEMux
    port map (
            O => \N__27259\,
            I => \N__27256\
        );

    \I__4308\ : LocalMux
    port map (
            O => \N__27256\,
            I => n12116
        );

    \I__4307\ : CascadeMux
    port map (
            O => \N__27253\,
            I => \n12116_cascade_\
        );

    \I__4306\ : SRMux
    port map (
            O => \N__27250\,
            I => \N__27247\
        );

    \I__4305\ : LocalMux
    port map (
            O => \N__27247\,
            I => \N__27244\
        );

    \I__4304\ : Span4Mux_h
    port map (
            O => \N__27244\,
            I => \N__27241\
        );

    \I__4303\ : Odrv4
    port map (
            O => \N__27241\,
            I => n14756
        );

    \I__4302\ : CascadeMux
    port map (
            O => \N__27238\,
            I => \n25_adj_1592_cascade_\
        );

    \I__4301\ : CascadeMux
    port map (
            O => \N__27235\,
            I => \n11944_cascade_\
        );

    \I__4300\ : CascadeMux
    port map (
            O => \N__27232\,
            I => \n11941_cascade_\
        );

    \I__4299\ : CascadeMux
    port map (
            O => \N__27229\,
            I => \n21919_cascade_\
        );

    \I__4298\ : InMux
    port map (
            O => \N__27226\,
            I => \N__27223\
        );

    \I__4297\ : LocalMux
    port map (
            O => \N__27223\,
            I => \N__27220\
        );

    \I__4296\ : Span4Mux_h
    port map (
            O => \N__27220\,
            I => \N__27217\
        );

    \I__4295\ : Span4Mux_v
    port map (
            O => \N__27217\,
            I => \N__27214\
        );

    \I__4294\ : Span4Mux_v
    port map (
            O => \N__27214\,
            I => \N__27211\
        );

    \I__4293\ : Odrv4
    port map (
            O => \N__27211\,
            I => buf_data_vac_23
        );

    \I__4292\ : InMux
    port map (
            O => \N__27208\,
            I => \N__27205\
        );

    \I__4291\ : LocalMux
    port map (
            O => \N__27205\,
            I => \N__27202\
        );

    \I__4290\ : Span4Mux_h
    port map (
            O => \N__27202\,
            I => \N__27199\
        );

    \I__4289\ : Span4Mux_h
    port map (
            O => \N__27199\,
            I => \N__27196\
        );

    \I__4288\ : Span4Mux_v
    port map (
            O => \N__27196\,
            I => \N__27193\
        );

    \I__4287\ : Odrv4
    port map (
            O => \N__27193\,
            I => buf_data_vac_22
        );

    \I__4286\ : CascadeMux
    port map (
            O => \N__27190\,
            I => \N__27187\
        );

    \I__4285\ : InMux
    port map (
            O => \N__27187\,
            I => \N__27184\
        );

    \I__4284\ : LocalMux
    port map (
            O => \N__27184\,
            I => \N__27181\
        );

    \I__4283\ : Span12Mux_h
    port map (
            O => \N__27181\,
            I => \N__27178\
        );

    \I__4282\ : Odrv12
    port map (
            O => \N__27178\,
            I => buf_data_vac_21
        );

    \I__4281\ : InMux
    port map (
            O => \N__27175\,
            I => \N__27172\
        );

    \I__4280\ : LocalMux
    port map (
            O => \N__27172\,
            I => \N__27169\
        );

    \I__4279\ : Span4Mux_h
    port map (
            O => \N__27169\,
            I => \N__27166\
        );

    \I__4278\ : Span4Mux_h
    port map (
            O => \N__27166\,
            I => \N__27163\
        );

    \I__4277\ : Span4Mux_v
    port map (
            O => \N__27163\,
            I => \N__27160\
        );

    \I__4276\ : Odrv4
    port map (
            O => \N__27160\,
            I => buf_data_vac_20
        );

    \I__4275\ : InMux
    port map (
            O => \N__27157\,
            I => \N__27154\
        );

    \I__4274\ : LocalMux
    port map (
            O => \N__27154\,
            I => \N__27151\
        );

    \I__4273\ : Odrv12
    port map (
            O => \N__27151\,
            I => buf_data_vac_19
        );

    \I__4272\ : InMux
    port map (
            O => \N__27148\,
            I => \N__27145\
        );

    \I__4271\ : LocalMux
    port map (
            O => \N__27145\,
            I => \N__27142\
        );

    \I__4270\ : Span4Mux_h
    port map (
            O => \N__27142\,
            I => \N__27139\
        );

    \I__4269\ : Span4Mux_h
    port map (
            O => \N__27139\,
            I => \N__27136\
        );

    \I__4268\ : Odrv4
    port map (
            O => \N__27136\,
            I => buf_data_vac_18
        );

    \I__4267\ : InMux
    port map (
            O => \N__27133\,
            I => \N__27130\
        );

    \I__4266\ : LocalMux
    port map (
            O => \N__27130\,
            I => \N__27127\
        );

    \I__4265\ : Span4Mux_v
    port map (
            O => \N__27127\,
            I => \N__27124\
        );

    \I__4264\ : Span4Mux_h
    port map (
            O => \N__27124\,
            I => \N__27121\
        );

    \I__4263\ : Odrv4
    port map (
            O => \N__27121\,
            I => buf_data_vac_17
        );

    \I__4262\ : CascadeMux
    port map (
            O => \N__27118\,
            I => \n21143_cascade_\
        );

    \I__4261\ : InMux
    port map (
            O => \N__27115\,
            I => \N__27111\
        );

    \I__4260\ : InMux
    port map (
            O => \N__27114\,
            I => \N__27108\
        );

    \I__4259\ : LocalMux
    port map (
            O => \N__27111\,
            I => cmd_rdadcbuf_18
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__27108\,
            I => cmd_rdadcbuf_18
        );

    \I__4257\ : InMux
    port map (
            O => \N__27103\,
            I => \N__27099\
        );

    \I__4256\ : InMux
    port map (
            O => \N__27102\,
            I => \N__27096\
        );

    \I__4255\ : LocalMux
    port map (
            O => \N__27099\,
            I => cmd_rdadcbuf_17
        );

    \I__4254\ : LocalMux
    port map (
            O => \N__27096\,
            I => cmd_rdadcbuf_17
        );

    \I__4253\ : CascadeMux
    port map (
            O => \N__27091\,
            I => \N__27088\
        );

    \I__4252\ : InMux
    port map (
            O => \N__27088\,
            I => \N__27084\
        );

    \I__4251\ : InMux
    port map (
            O => \N__27087\,
            I => \N__27081\
        );

    \I__4250\ : LocalMux
    port map (
            O => \N__27084\,
            I => cmd_rdadcbuf_16
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__27081\,
            I => cmd_rdadcbuf_16
        );

    \I__4248\ : InMux
    port map (
            O => \N__27076\,
            I => \N__27073\
        );

    \I__4247\ : LocalMux
    port map (
            O => \N__27073\,
            I => \N__27070\
        );

    \I__4246\ : Odrv12
    port map (
            O => \N__27070\,
            I => \ADC_VDC.n18394\
        );

    \I__4245\ : InMux
    port map (
            O => \N__27067\,
            I => \N__27064\
        );

    \I__4244\ : LocalMux
    port map (
            O => \N__27064\,
            I => \N__27061\
        );

    \I__4243\ : Odrv4
    port map (
            O => \N__27061\,
            I => \ADC_VDC.cmd_rdadcbuf_35_N_1130_34\
        );

    \I__4242\ : CascadeMux
    port map (
            O => \N__27058\,
            I => \ADC_VDC.n21106_cascade_\
        );

    \I__4241\ : InMux
    port map (
            O => \N__27055\,
            I => \N__27052\
        );

    \I__4240\ : LocalMux
    port map (
            O => \N__27052\,
            I => \N__27049\
        );

    \I__4239\ : Span4Mux_h
    port map (
            O => \N__27049\,
            I => \N__27044\
        );

    \I__4238\ : InMux
    port map (
            O => \N__27048\,
            I => \N__27041\
        );

    \I__4237\ : InMux
    port map (
            O => \N__27047\,
            I => \N__27038\
        );

    \I__4236\ : Odrv4
    port map (
            O => \N__27044\,
            I => cmd_rdadcbuf_34
        );

    \I__4235\ : LocalMux
    port map (
            O => \N__27041\,
            I => cmd_rdadcbuf_34
        );

    \I__4234\ : LocalMux
    port map (
            O => \N__27038\,
            I => cmd_rdadcbuf_34
        );

    \I__4233\ : CEMux
    port map (
            O => \N__27031\,
            I => \N__27028\
        );

    \I__4232\ : LocalMux
    port map (
            O => \N__27028\,
            I => \N__27025\
        );

    \I__4231\ : Odrv4
    port map (
            O => \N__27025\,
            I => \ADC_VDC.n13020\
        );

    \I__4230\ : InMux
    port map (
            O => \N__27022\,
            I => \N__27019\
        );

    \I__4229\ : LocalMux
    port map (
            O => \N__27019\,
            I => \N__27016\
        );

    \I__4228\ : Odrv12
    port map (
            O => \N__27016\,
            I => \ADC_VDC.n21\
        );

    \I__4227\ : InMux
    port map (
            O => \N__27013\,
            I => \N__27010\
        );

    \I__4226\ : LocalMux
    port map (
            O => \N__27010\,
            I => \N__27007\
        );

    \I__4225\ : Odrv12
    port map (
            O => \N__27007\,
            I => \ADC_VDC.n19\
        );

    \I__4224\ : InMux
    port map (
            O => \N__27004\,
            I => \N__27001\
        );

    \I__4223\ : LocalMux
    port map (
            O => \N__27001\,
            I => \N__26998\
        );

    \I__4222\ : Span4Mux_h
    port map (
            O => \N__26998\,
            I => \N__26995\
        );

    \I__4221\ : Span4Mux_h
    port map (
            O => \N__26995\,
            I => \N__26992\
        );

    \I__4220\ : Odrv4
    port map (
            O => \N__26992\,
            I => buf_data_vac_16
        );

    \I__4219\ : InMux
    port map (
            O => \N__26989\,
            I => \N__26985\
        );

    \I__4218\ : CascadeMux
    port map (
            O => \N__26988\,
            I => \N__26981\
        );

    \I__4217\ : LocalMux
    port map (
            O => \N__26985\,
            I => \N__26978\
        );

    \I__4216\ : CascadeMux
    port map (
            O => \N__26984\,
            I => \N__26975\
        );

    \I__4215\ : InMux
    port map (
            O => \N__26981\,
            I => \N__26972\
        );

    \I__4214\ : Span4Mux_h
    port map (
            O => \N__26978\,
            I => \N__26969\
        );

    \I__4213\ : InMux
    port map (
            O => \N__26975\,
            I => \N__26966\
        );

    \I__4212\ : LocalMux
    port map (
            O => \N__26972\,
            I => cmd_rdadctmp_10_adj_1462
        );

    \I__4211\ : Odrv4
    port map (
            O => \N__26969\,
            I => cmd_rdadctmp_10_adj_1462
        );

    \I__4210\ : LocalMux
    port map (
            O => \N__26966\,
            I => cmd_rdadctmp_10_adj_1462
        );

    \I__4209\ : CascadeMux
    port map (
            O => \N__26959\,
            I => \N__26954\
        );

    \I__4208\ : InMux
    port map (
            O => \N__26958\,
            I => \N__26949\
        );

    \I__4207\ : InMux
    port map (
            O => \N__26957\,
            I => \N__26949\
        );

    \I__4206\ : InMux
    port map (
            O => \N__26954\,
            I => \N__26946\
        );

    \I__4205\ : LocalMux
    port map (
            O => \N__26949\,
            I => cmd_rdadctmp_11_adj_1461
        );

    \I__4204\ : LocalMux
    port map (
            O => \N__26946\,
            I => cmd_rdadctmp_11_adj_1461
        );

    \I__4203\ : CascadeMux
    port map (
            O => \N__26941\,
            I => \ADC_VDC.n21673_cascade_\
        );

    \I__4202\ : IoInMux
    port map (
            O => \N__26938\,
            I => \N__26935\
        );

    \I__4201\ : LocalMux
    port map (
            O => \N__26935\,
            I => \N__26932\
        );

    \I__4200\ : Span12Mux_s11_h
    port map (
            O => \N__26932\,
            I => \N__26928\
        );

    \I__4199\ : InMux
    port map (
            O => \N__26931\,
            I => \N__26925\
        );

    \I__4198\ : Odrv12
    port map (
            O => \N__26928\,
            I => \VDC_SCLK\
        );

    \I__4197\ : LocalMux
    port map (
            O => \N__26925\,
            I => \VDC_SCLK\
        );

    \I__4196\ : InMux
    port map (
            O => \N__26920\,
            I => \N__26916\
        );

    \I__4195\ : CascadeMux
    port map (
            O => \N__26919\,
            I => \N__26912\
        );

    \I__4194\ : LocalMux
    port map (
            O => \N__26916\,
            I => \N__26909\
        );

    \I__4193\ : InMux
    port map (
            O => \N__26915\,
            I => \N__26906\
        );

    \I__4192\ : InMux
    port map (
            O => \N__26912\,
            I => \N__26903\
        );

    \I__4191\ : Odrv4
    port map (
            O => \N__26909\,
            I => cmd_rdadctmp_19_adj_1453
        );

    \I__4190\ : LocalMux
    port map (
            O => \N__26906\,
            I => cmd_rdadctmp_19_adj_1453
        );

    \I__4189\ : LocalMux
    port map (
            O => \N__26903\,
            I => cmd_rdadctmp_19_adj_1453
        );

    \I__4188\ : CascadeMux
    port map (
            O => \N__26896\,
            I => \N__26892\
        );

    \I__4187\ : CascadeMux
    port map (
            O => \N__26895\,
            I => \N__26885\
        );

    \I__4186\ : InMux
    port map (
            O => \N__26892\,
            I => \N__26875\
        );

    \I__4185\ : InMux
    port map (
            O => \N__26891\,
            I => \N__26864\
        );

    \I__4184\ : InMux
    port map (
            O => \N__26890\,
            I => \N__26864\
        );

    \I__4183\ : InMux
    port map (
            O => \N__26889\,
            I => \N__26864\
        );

    \I__4182\ : InMux
    port map (
            O => \N__26888\,
            I => \N__26864\
        );

    \I__4181\ : InMux
    port map (
            O => \N__26885\,
            I => \N__26864\
        );

    \I__4180\ : CascadeMux
    port map (
            O => \N__26884\,
            I => \N__26861\
        );

    \I__4179\ : CascadeMux
    port map (
            O => \N__26883\,
            I => \N__26858\
        );

    \I__4178\ : CascadeMux
    port map (
            O => \N__26882\,
            I => \N__26855\
        );

    \I__4177\ : CascadeMux
    port map (
            O => \N__26881\,
            I => \N__26852\
        );

    \I__4176\ : CascadeMux
    port map (
            O => \N__26880\,
            I => \N__26847\
        );

    \I__4175\ : CascadeMux
    port map (
            O => \N__26879\,
            I => \N__26843\
        );

    \I__4174\ : CascadeMux
    port map (
            O => \N__26878\,
            I => \N__26838\
        );

    \I__4173\ : LocalMux
    port map (
            O => \N__26875\,
            I => \N__26831\
        );

    \I__4172\ : LocalMux
    port map (
            O => \N__26864\,
            I => \N__26831\
        );

    \I__4171\ : InMux
    port map (
            O => \N__26861\,
            I => \N__26818\
        );

    \I__4170\ : InMux
    port map (
            O => \N__26858\,
            I => \N__26818\
        );

    \I__4169\ : InMux
    port map (
            O => \N__26855\,
            I => \N__26818\
        );

    \I__4168\ : InMux
    port map (
            O => \N__26852\,
            I => \N__26818\
        );

    \I__4167\ : InMux
    port map (
            O => \N__26851\,
            I => \N__26818\
        );

    \I__4166\ : InMux
    port map (
            O => \N__26850\,
            I => \N__26818\
        );

    \I__4165\ : InMux
    port map (
            O => \N__26847\,
            I => \N__26805\
        );

    \I__4164\ : InMux
    port map (
            O => \N__26846\,
            I => \N__26805\
        );

    \I__4163\ : InMux
    port map (
            O => \N__26843\,
            I => \N__26805\
        );

    \I__4162\ : InMux
    port map (
            O => \N__26842\,
            I => \N__26805\
        );

    \I__4161\ : InMux
    port map (
            O => \N__26841\,
            I => \N__26805\
        );

    \I__4160\ : InMux
    port map (
            O => \N__26838\,
            I => \N__26805\
        );

    \I__4159\ : CascadeMux
    port map (
            O => \N__26837\,
            I => \N__26802\
        );

    \I__4158\ : CascadeMux
    port map (
            O => \N__26836\,
            I => \N__26799\
        );

    \I__4157\ : Span4Mux_v
    port map (
            O => \N__26831\,
            I => \N__26792\
        );

    \I__4156\ : LocalMux
    port map (
            O => \N__26818\,
            I => \N__26792\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__26805\,
            I => \N__26789\
        );

    \I__4154\ : InMux
    port map (
            O => \N__26802\,
            I => \N__26780\
        );

    \I__4153\ : InMux
    port map (
            O => \N__26799\,
            I => \N__26780\
        );

    \I__4152\ : InMux
    port map (
            O => \N__26798\,
            I => \N__26780\
        );

    \I__4151\ : InMux
    port map (
            O => \N__26797\,
            I => \N__26780\
        );

    \I__4150\ : Odrv4
    port map (
            O => \N__26792\,
            I => n12853
        );

    \I__4149\ : Odrv4
    port map (
            O => \N__26789\,
            I => n12853
        );

    \I__4148\ : LocalMux
    port map (
            O => \N__26780\,
            I => n12853
        );

    \I__4147\ : CascadeMux
    port map (
            O => \N__26773\,
            I => \N__26770\
        );

    \I__4146\ : InMux
    port map (
            O => \N__26770\,
            I => \N__26765\
        );

    \I__4145\ : CascadeMux
    port map (
            O => \N__26769\,
            I => \N__26762\
        );

    \I__4144\ : InMux
    port map (
            O => \N__26768\,
            I => \N__26759\
        );

    \I__4143\ : LocalMux
    port map (
            O => \N__26765\,
            I => \N__26756\
        );

    \I__4142\ : InMux
    port map (
            O => \N__26762\,
            I => \N__26753\
        );

    \I__4141\ : LocalMux
    port map (
            O => \N__26759\,
            I => cmd_rdadctmp_20_adj_1452
        );

    \I__4140\ : Odrv12
    port map (
            O => \N__26756\,
            I => cmd_rdadctmp_20_adj_1452
        );

    \I__4139\ : LocalMux
    port map (
            O => \N__26753\,
            I => cmd_rdadctmp_20_adj_1452
        );

    \I__4138\ : InMux
    port map (
            O => \N__26746\,
            I => \N__26742\
        );

    \I__4137\ : InMux
    port map (
            O => \N__26745\,
            I => \N__26739\
        );

    \I__4136\ : LocalMux
    port map (
            O => \N__26742\,
            I => cmd_rdadcbuf_23
        );

    \I__4135\ : LocalMux
    port map (
            O => \N__26739\,
            I => cmd_rdadcbuf_23
        );

    \I__4134\ : InMux
    port map (
            O => \N__26734\,
            I => \N__26731\
        );

    \I__4133\ : LocalMux
    port map (
            O => \N__26731\,
            I => \N__26728\
        );

    \I__4132\ : Span4Mux_v
    port map (
            O => \N__26728\,
            I => \N__26724\
        );

    \I__4131\ : CascadeMux
    port map (
            O => \N__26727\,
            I => \N__26721\
        );

    \I__4130\ : Span4Mux_v
    port map (
            O => \N__26724\,
            I => \N__26718\
        );

    \I__4129\ : InMux
    port map (
            O => \N__26721\,
            I => \N__26715\
        );

    \I__4128\ : Odrv4
    port map (
            O => \N__26718\,
            I => buf_adcdata_vdc_12
        );

    \I__4127\ : LocalMux
    port map (
            O => \N__26715\,
            I => buf_adcdata_vdc_12
        );

    \I__4126\ : InMux
    port map (
            O => \N__26710\,
            I => \N__26706\
        );

    \I__4125\ : InMux
    port map (
            O => \N__26709\,
            I => \N__26703\
        );

    \I__4124\ : LocalMux
    port map (
            O => \N__26706\,
            I => cmd_rdadcbuf_22
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__26703\,
            I => cmd_rdadcbuf_22
        );

    \I__4122\ : InMux
    port map (
            O => \N__26698\,
            I => \N__26695\
        );

    \I__4121\ : LocalMux
    port map (
            O => \N__26695\,
            I => \N__26692\
        );

    \I__4120\ : Span4Mux_v
    port map (
            O => \N__26692\,
            I => \N__26688\
        );

    \I__4119\ : CascadeMux
    port map (
            O => \N__26691\,
            I => \N__26685\
        );

    \I__4118\ : Span4Mux_v
    port map (
            O => \N__26688\,
            I => \N__26682\
        );

    \I__4117\ : InMux
    port map (
            O => \N__26685\,
            I => \N__26679\
        );

    \I__4116\ : Odrv4
    port map (
            O => \N__26682\,
            I => buf_adcdata_vdc_11
        );

    \I__4115\ : LocalMux
    port map (
            O => \N__26679\,
            I => buf_adcdata_vdc_11
        );

    \I__4114\ : CascadeMux
    port map (
            O => \N__26674\,
            I => \N__26671\
        );

    \I__4113\ : InMux
    port map (
            O => \N__26671\,
            I => \N__26667\
        );

    \I__4112\ : InMux
    port map (
            O => \N__26670\,
            I => \N__26664\
        );

    \I__4111\ : LocalMux
    port map (
            O => \N__26667\,
            I => cmd_rdadcbuf_15
        );

    \I__4110\ : LocalMux
    port map (
            O => \N__26664\,
            I => cmd_rdadcbuf_15
        );

    \I__4109\ : InMux
    port map (
            O => \N__26659\,
            I => \N__26655\
        );

    \I__4108\ : InMux
    port map (
            O => \N__26658\,
            I => \N__26652\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__26655\,
            I => cmd_rdadcbuf_20
        );

    \I__4106\ : LocalMux
    port map (
            O => \N__26652\,
            I => cmd_rdadcbuf_20
        );

    \I__4105\ : InMux
    port map (
            O => \N__26647\,
            I => \N__26643\
        );

    \I__4104\ : InMux
    port map (
            O => \N__26646\,
            I => \N__26640\
        );

    \I__4103\ : LocalMux
    port map (
            O => \N__26643\,
            I => cmd_rdadcbuf_19
        );

    \I__4102\ : LocalMux
    port map (
            O => \N__26640\,
            I => cmd_rdadcbuf_19
        );

    \I__4101\ : InMux
    port map (
            O => \N__26635\,
            I => \N__26632\
        );

    \I__4100\ : LocalMux
    port map (
            O => \N__26632\,
            I => \N__26629\
        );

    \I__4099\ : Span4Mux_h
    port map (
            O => \N__26629\,
            I => \N__26625\
        );

    \I__4098\ : CascadeMux
    port map (
            O => \N__26628\,
            I => \N__26622\
        );

    \I__4097\ : Span4Mux_v
    port map (
            O => \N__26625\,
            I => \N__26619\
        );

    \I__4096\ : InMux
    port map (
            O => \N__26622\,
            I => \N__26616\
        );

    \I__4095\ : Odrv4
    port map (
            O => \N__26619\,
            I => buf_adcdata_vdc_8
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__26616\,
            I => buf_adcdata_vdc_8
        );

    \I__4093\ : CascadeMux
    port map (
            O => \N__26611\,
            I => \N__26606\
        );

    \I__4092\ : InMux
    port map (
            O => \N__26610\,
            I => \N__26603\
        );

    \I__4091\ : InMux
    port map (
            O => \N__26609\,
            I => \N__26600\
        );

    \I__4090\ : InMux
    port map (
            O => \N__26606\,
            I => \N__26597\
        );

    \I__4089\ : LocalMux
    port map (
            O => \N__26603\,
            I => cmd_rdadctmp_0_adj_1472
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__26600\,
            I => cmd_rdadctmp_0_adj_1472
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__26597\,
            I => cmd_rdadctmp_0_adj_1472
        );

    \I__4086\ : CascadeMux
    port map (
            O => \N__26590\,
            I => \N__26587\
        );

    \I__4085\ : InMux
    port map (
            O => \N__26587\,
            I => \N__26582\
        );

    \I__4084\ : InMux
    port map (
            O => \N__26586\,
            I => \N__26577\
        );

    \I__4083\ : InMux
    port map (
            O => \N__26585\,
            I => \N__26577\
        );

    \I__4082\ : LocalMux
    port map (
            O => \N__26582\,
            I => \N__26574\
        );

    \I__4081\ : LocalMux
    port map (
            O => \N__26577\,
            I => cmd_rdadctmp_3_adj_1469
        );

    \I__4080\ : Odrv4
    port map (
            O => \N__26574\,
            I => cmd_rdadctmp_3_adj_1469
        );

    \I__4079\ : InMux
    port map (
            O => \N__26569\,
            I => \N__26565\
        );

    \I__4078\ : CascadeMux
    port map (
            O => \N__26568\,
            I => \N__26561\
        );

    \I__4077\ : LocalMux
    port map (
            O => \N__26565\,
            I => \N__26558\
        );

    \I__4076\ : InMux
    port map (
            O => \N__26564\,
            I => \N__26555\
        );

    \I__4075\ : InMux
    port map (
            O => \N__26561\,
            I => \N__26552\
        );

    \I__4074\ : Odrv4
    port map (
            O => \N__26558\,
            I => cmd_rdadctmp_4_adj_1468
        );

    \I__4073\ : LocalMux
    port map (
            O => \N__26555\,
            I => cmd_rdadctmp_4_adj_1468
        );

    \I__4072\ : LocalMux
    port map (
            O => \N__26552\,
            I => cmd_rdadctmp_4_adj_1468
        );

    \I__4071\ : CEMux
    port map (
            O => \N__26545\,
            I => \N__26542\
        );

    \I__4070\ : LocalMux
    port map (
            O => \N__26542\,
            I => \N__26539\
        );

    \I__4069\ : Span4Mux_h
    port map (
            O => \N__26539\,
            I => \N__26536\
        );

    \I__4068\ : Odrv4
    port map (
            O => \N__26536\,
            I => \ADC_VDC.n12885\
        );

    \I__4067\ : CascadeMux
    port map (
            O => \N__26533\,
            I => \N__26529\
        );

    \I__4066\ : InMux
    port map (
            O => \N__26532\,
            I => \N__26525\
        );

    \I__4065\ : InMux
    port map (
            O => \N__26529\,
            I => \N__26522\
        );

    \I__4064\ : InMux
    port map (
            O => \N__26528\,
            I => \N__26519\
        );

    \I__4063\ : LocalMux
    port map (
            O => \N__26525\,
            I => \N__26514\
        );

    \I__4062\ : LocalMux
    port map (
            O => \N__26522\,
            I => \N__26514\
        );

    \I__4061\ : LocalMux
    port map (
            O => \N__26519\,
            I => cmd_rdadctmp_7_adj_1465
        );

    \I__4060\ : Odrv4
    port map (
            O => \N__26514\,
            I => cmd_rdadctmp_7_adj_1465
        );

    \I__4059\ : InMux
    port map (
            O => \N__26509\,
            I => \N__26505\
        );

    \I__4058\ : CascadeMux
    port map (
            O => \N__26508\,
            I => \N__26501\
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__26505\,
            I => \N__26498\
        );

    \I__4056\ : InMux
    port map (
            O => \N__26504\,
            I => \N__26495\
        );

    \I__4055\ : InMux
    port map (
            O => \N__26501\,
            I => \N__26492\
        );

    \I__4054\ : Odrv4
    port map (
            O => \N__26498\,
            I => cmd_rdadctmp_8_adj_1464
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__26495\,
            I => cmd_rdadctmp_8_adj_1464
        );

    \I__4052\ : LocalMux
    port map (
            O => \N__26492\,
            I => cmd_rdadctmp_8_adj_1464
        );

    \I__4051\ : CascadeMux
    port map (
            O => \N__26485\,
            I => \N__26482\
        );

    \I__4050\ : InMux
    port map (
            O => \N__26482\,
            I => \N__26477\
        );

    \I__4049\ : CascadeMux
    port map (
            O => \N__26481\,
            I => \N__26474\
        );

    \I__4048\ : InMux
    port map (
            O => \N__26480\,
            I => \N__26471\
        );

    \I__4047\ : LocalMux
    port map (
            O => \N__26477\,
            I => \N__26468\
        );

    \I__4046\ : InMux
    port map (
            O => \N__26474\,
            I => \N__26465\
        );

    \I__4045\ : LocalMux
    port map (
            O => \N__26471\,
            I => cmd_rdadctmp_17_adj_1455
        );

    \I__4044\ : Odrv12
    port map (
            O => \N__26468\,
            I => cmd_rdadctmp_17_adj_1455
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__26465\,
            I => cmd_rdadctmp_17_adj_1455
        );

    \I__4042\ : CascadeMux
    port map (
            O => \N__26458\,
            I => \N__26455\
        );

    \I__4041\ : InMux
    port map (
            O => \N__26455\,
            I => \N__26452\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__26452\,
            I => \N__26447\
        );

    \I__4039\ : CascadeMux
    port map (
            O => \N__26451\,
            I => \N__26444\
        );

    \I__4038\ : InMux
    port map (
            O => \N__26450\,
            I => \N__26441\
        );

    \I__4037\ : Span4Mux_h
    port map (
            O => \N__26447\,
            I => \N__26438\
        );

    \I__4036\ : InMux
    port map (
            O => \N__26444\,
            I => \N__26435\
        );

    \I__4035\ : LocalMux
    port map (
            O => \N__26441\,
            I => cmd_rdadctmp_15_adj_1457
        );

    \I__4034\ : Odrv4
    port map (
            O => \N__26438\,
            I => cmd_rdadctmp_15_adj_1457
        );

    \I__4033\ : LocalMux
    port map (
            O => \N__26435\,
            I => cmd_rdadctmp_15_adj_1457
        );

    \I__4032\ : CascadeMux
    port map (
            O => \N__26428\,
            I => \N__26423\
        );

    \I__4031\ : InMux
    port map (
            O => \N__26427\,
            I => \N__26418\
        );

    \I__4030\ : InMux
    port map (
            O => \N__26426\,
            I => \N__26418\
        );

    \I__4029\ : InMux
    port map (
            O => \N__26423\,
            I => \N__26415\
        );

    \I__4028\ : LocalMux
    port map (
            O => \N__26418\,
            I => cmd_rdadctmp_16_adj_1456
        );

    \I__4027\ : LocalMux
    port map (
            O => \N__26415\,
            I => cmd_rdadctmp_16_adj_1456
        );

    \I__4026\ : CascadeMux
    port map (
            O => \N__26410\,
            I => \N__26405\
        );

    \I__4025\ : InMux
    port map (
            O => \N__26409\,
            I => \N__26402\
        );

    \I__4024\ : InMux
    port map (
            O => \N__26408\,
            I => \N__26399\
        );

    \I__4023\ : InMux
    port map (
            O => \N__26405\,
            I => \N__26396\
        );

    \I__4022\ : LocalMux
    port map (
            O => \N__26402\,
            I => cmd_rdadctmp_1_adj_1471
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__26399\,
            I => cmd_rdadctmp_1_adj_1471
        );

    \I__4020\ : LocalMux
    port map (
            O => \N__26396\,
            I => cmd_rdadctmp_1_adj_1471
        );

    \I__4019\ : CascadeMux
    port map (
            O => \N__26389\,
            I => \N__26384\
        );

    \I__4018\ : InMux
    port map (
            O => \N__26388\,
            I => \N__26381\
        );

    \I__4017\ : InMux
    port map (
            O => \N__26387\,
            I => \N__26378\
        );

    \I__4016\ : InMux
    port map (
            O => \N__26384\,
            I => \N__26375\
        );

    \I__4015\ : LocalMux
    port map (
            O => \N__26381\,
            I => \N__26372\
        );

    \I__4014\ : LocalMux
    port map (
            O => \N__26378\,
            I => cmd_rdadctmp_2_adj_1470
        );

    \I__4013\ : LocalMux
    port map (
            O => \N__26375\,
            I => cmd_rdadctmp_2_adj_1470
        );

    \I__4012\ : Odrv4
    port map (
            O => \N__26372\,
            I => cmd_rdadctmp_2_adj_1470
        );

    \I__4011\ : CascadeMux
    port map (
            O => \N__26365\,
            I => \N__26360\
        );

    \I__4010\ : CascadeMux
    port map (
            O => \N__26364\,
            I => \N__26357\
        );

    \I__4009\ : InMux
    port map (
            O => \N__26363\,
            I => \N__26354\
        );

    \I__4008\ : InMux
    port map (
            O => \N__26360\,
            I => \N__26351\
        );

    \I__4007\ : InMux
    port map (
            O => \N__26357\,
            I => \N__26348\
        );

    \I__4006\ : LocalMux
    port map (
            O => \N__26354\,
            I => \N__26345\
        );

    \I__4005\ : LocalMux
    port map (
            O => \N__26351\,
            I => \N__26342\
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__26348\,
            I => cmd_rdadctmp_12_adj_1460
        );

    \I__4003\ : Odrv4
    port map (
            O => \N__26345\,
            I => cmd_rdadctmp_12_adj_1460
        );

    \I__4002\ : Odrv4
    port map (
            O => \N__26342\,
            I => cmd_rdadctmp_12_adj_1460
        );

    \I__4001\ : CascadeMux
    port map (
            O => \N__26335\,
            I => \ADC_VDC.n31_cascade_\
        );

    \I__4000\ : CascadeMux
    port map (
            O => \N__26332\,
            I => \ADC_VDC.n21925_cascade_\
        );

    \I__3999\ : InMux
    port map (
            O => \N__26329\,
            I => \N__26326\
        );

    \I__3998\ : LocalMux
    port map (
            O => \N__26326\,
            I => \ADC_VDC.n18397\
        );

    \I__3997\ : CascadeMux
    port map (
            O => \N__26323\,
            I => \ADC_VDC.n21928_cascade_\
        );

    \I__3996\ : CEMux
    port map (
            O => \N__26320\,
            I => \N__26317\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__26317\,
            I => \N__26314\
        );

    \I__3994\ : Odrv4
    port map (
            O => \N__26314\,
            I => \ADC_VDC.n20514\
        );

    \I__3993\ : CascadeMux
    port map (
            O => \N__26311\,
            I => \ADC_VDC.n6_cascade_\
        );

    \I__3992\ : InMux
    port map (
            O => \N__26308\,
            I => \N__26304\
        );

    \I__3991\ : InMux
    port map (
            O => \N__26307\,
            I => \N__26301\
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__26304\,
            I => \ADC_VDC.n10519\
        );

    \I__3989\ : LocalMux
    port map (
            O => \N__26301\,
            I => \ADC_VDC.n10519\
        );

    \I__3988\ : CascadeMux
    port map (
            O => \N__26296\,
            I => \n12853_cascade_\
        );

    \I__3987\ : CascadeMux
    port map (
            O => \N__26293\,
            I => \N__26289\
        );

    \I__3986\ : CascadeMux
    port map (
            O => \N__26292\,
            I => \N__26286\
        );

    \I__3985\ : InMux
    port map (
            O => \N__26289\,
            I => \N__26283\
        );

    \I__3984\ : InMux
    port map (
            O => \N__26286\,
            I => \N__26280\
        );

    \I__3983\ : LocalMux
    port map (
            O => \N__26283\,
            I => cmd_rdadctmp_31
        );

    \I__3982\ : LocalMux
    port map (
            O => \N__26280\,
            I => cmd_rdadctmp_31
        );

    \I__3981\ : InMux
    port map (
            O => \N__26275\,
            I => \N__26272\
        );

    \I__3980\ : LocalMux
    port map (
            O => \N__26272\,
            I => \N__26269\
        );

    \I__3979\ : Span4Mux_v
    port map (
            O => \N__26269\,
            I => \N__26266\
        );

    \I__3978\ : Span4Mux_v
    port map (
            O => \N__26266\,
            I => \N__26263\
        );

    \I__3977\ : Span4Mux_h
    port map (
            O => \N__26263\,
            I => \N__26259\
        );

    \I__3976\ : CascadeMux
    port map (
            O => \N__26262\,
            I => \N__26255\
        );

    \I__3975\ : Sp12to4
    port map (
            O => \N__26259\,
            I => \N__26252\
        );

    \I__3974\ : InMux
    port map (
            O => \N__26258\,
            I => \N__26247\
        );

    \I__3973\ : InMux
    port map (
            O => \N__26255\,
            I => \N__26247\
        );

    \I__3972\ : Odrv12
    port map (
            O => \N__26252\,
            I => buf_adcdata_iac_23
        );

    \I__3971\ : LocalMux
    port map (
            O => \N__26247\,
            I => buf_adcdata_iac_23
        );

    \I__3970\ : IoInMux
    port map (
            O => \N__26242\,
            I => \N__26239\
        );

    \I__3969\ : LocalMux
    port map (
            O => \N__26239\,
            I => \N__26236\
        );

    \I__3968\ : Span4Mux_s0_v
    port map (
            O => \N__26236\,
            I => \N__26233\
        );

    \I__3967\ : Span4Mux_v
    port map (
            O => \N__26233\,
            I => \N__26230\
        );

    \I__3966\ : Span4Mux_v
    port map (
            O => \N__26230\,
            I => \N__26227\
        );

    \I__3965\ : Sp12to4
    port map (
            O => \N__26227\,
            I => \N__26224\
        );

    \I__3964\ : Odrv12
    port map (
            O => \N__26224\,
            I => \AC_ADC_SYNC\
        );

    \I__3963\ : IoInMux
    port map (
            O => \N__26221\,
            I => \N__26218\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__26218\,
            I => \N__26215\
        );

    \I__3961\ : Span4Mux_s3_h
    port map (
            O => \N__26215\,
            I => \N__26212\
        );

    \I__3960\ : Span4Mux_v
    port map (
            O => \N__26212\,
            I => \N__26209\
        );

    \I__3959\ : Sp12to4
    port map (
            O => \N__26209\,
            I => \N__26204\
        );

    \I__3958\ : InMux
    port map (
            O => \N__26208\,
            I => \N__26199\
        );

    \I__3957\ : InMux
    port map (
            O => \N__26207\,
            I => \N__26199\
        );

    \I__3956\ : Odrv12
    port map (
            O => \N__26204\,
            I => \VAC_FLT1\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__26199\,
            I => \VAC_FLT1\
        );

    \I__3954\ : IoInMux
    port map (
            O => \N__26194\,
            I => \N__26191\
        );

    \I__3953\ : LocalMux
    port map (
            O => \N__26191\,
            I => \N__26188\
        );

    \I__3952\ : Span4Mux_s3_v
    port map (
            O => \N__26188\,
            I => \N__26185\
        );

    \I__3951\ : Span4Mux_h
    port map (
            O => \N__26185\,
            I => \N__26181\
        );

    \I__3950\ : CascadeMux
    port map (
            O => \N__26184\,
            I => \N__26178\
        );

    \I__3949\ : Span4Mux_v
    port map (
            O => \N__26181\,
            I => \N__26175\
        );

    \I__3948\ : InMux
    port map (
            O => \N__26178\,
            I => \N__26172\
        );

    \I__3947\ : Odrv4
    port map (
            O => \N__26175\,
            I => \IAC_SCLK\
        );

    \I__3946\ : LocalMux
    port map (
            O => \N__26172\,
            I => \IAC_SCLK\
        );

    \I__3945\ : CascadeMux
    port map (
            O => \N__26167\,
            I => \ADC_VDC.n18394_cascade_\
        );

    \I__3944\ : InMux
    port map (
            O => \N__26164\,
            I => \N__26161\
        );

    \I__3943\ : LocalMux
    port map (
            O => \N__26161\,
            I => \N__26158\
        );

    \I__3942\ : Sp12to4
    port map (
            O => \N__26158\,
            I => \N__26155\
        );

    \I__3941\ : Odrv12
    port map (
            O => \N__26155\,
            I => \EIS_SYNCCLK\
        );

    \I__3940\ : IoInMux
    port map (
            O => \N__26152\,
            I => \N__26149\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__26149\,
            I => \N__26145\
        );

    \I__3938\ : IoInMux
    port map (
            O => \N__26148\,
            I => \N__26142\
        );

    \I__3937\ : Span4Mux_s3_v
    port map (
            O => \N__26145\,
            I => \N__26139\
        );

    \I__3936\ : LocalMux
    port map (
            O => \N__26142\,
            I => \N__26136\
        );

    \I__3935\ : Span4Mux_h
    port map (
            O => \N__26139\,
            I => \N__26133\
        );

    \I__3934\ : Span4Mux_s3_h
    port map (
            O => \N__26136\,
            I => \N__26130\
        );

    \I__3933\ : Sp12to4
    port map (
            O => \N__26133\,
            I => \N__26127\
        );

    \I__3932\ : Span4Mux_v
    port map (
            O => \N__26130\,
            I => \N__26124\
        );

    \I__3931\ : Span12Mux_s11_v
    port map (
            O => \N__26127\,
            I => \N__26119\
        );

    \I__3930\ : Sp12to4
    port map (
            O => \N__26124\,
            I => \N__26119\
        );

    \I__3929\ : Span12Mux_v
    port map (
            O => \N__26119\,
            I => \N__26116\
        );

    \I__3928\ : Odrv12
    port map (
            O => \N__26116\,
            I => \IAC_CLK\
        );

    \I__3927\ : IoInMux
    port map (
            O => \N__26113\,
            I => \N__26110\
        );

    \I__3926\ : LocalMux
    port map (
            O => \N__26110\,
            I => \N__26107\
        );

    \I__3925\ : Span4Mux_s3_h
    port map (
            O => \N__26107\,
            I => \N__26104\
        );

    \I__3924\ : Span4Mux_v
    port map (
            O => \N__26104\,
            I => \N__26101\
        );

    \I__3923\ : Span4Mux_v
    port map (
            O => \N__26101\,
            I => \N__26097\
        );

    \I__3922\ : InMux
    port map (
            O => \N__26100\,
            I => \N__26093\
        );

    \I__3921\ : Sp12to4
    port map (
            O => \N__26097\,
            I => \N__26090\
        );

    \I__3920\ : InMux
    port map (
            O => \N__26096\,
            I => \N__26087\
        );

    \I__3919\ : LocalMux
    port map (
            O => \N__26093\,
            I => \N__26084\
        );

    \I__3918\ : Odrv12
    port map (
            O => \N__26090\,
            I => \VAC_OSR0\
        );

    \I__3917\ : LocalMux
    port map (
            O => \N__26087\,
            I => \VAC_OSR0\
        );

    \I__3916\ : Odrv4
    port map (
            O => \N__26084\,
            I => \VAC_OSR0\
        );

    \I__3915\ : InMux
    port map (
            O => \N__26077\,
            I => \N__26074\
        );

    \I__3914\ : LocalMux
    port map (
            O => \N__26074\,
            I => \N__26071\
        );

    \I__3913\ : Span4Mux_h
    port map (
            O => \N__26071\,
            I => \N__26066\
        );

    \I__3912\ : CascadeMux
    port map (
            O => \N__26070\,
            I => \N__26063\
        );

    \I__3911\ : InMux
    port map (
            O => \N__26069\,
            I => \N__26060\
        );

    \I__3910\ : Span4Mux_v
    port map (
            O => \N__26066\,
            I => \N__26057\
        );

    \I__3909\ : InMux
    port map (
            O => \N__26063\,
            I => \N__26054\
        );

    \I__3908\ : LocalMux
    port map (
            O => \N__26060\,
            I => buf_adcdata_iac_19
        );

    \I__3907\ : Odrv4
    port map (
            O => \N__26057\,
            I => buf_adcdata_iac_19
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__26054\,
            I => buf_adcdata_iac_19
        );

    \I__3905\ : InMux
    port map (
            O => \N__26047\,
            I => \N__26044\
        );

    \I__3904\ : LocalMux
    port map (
            O => \N__26044\,
            I => \N__26041\
        );

    \I__3903\ : Odrv12
    port map (
            O => \N__26041\,
            I => n11417
        );

    \I__3902\ : InMux
    port map (
            O => \N__26038\,
            I => \N__26035\
        );

    \I__3901\ : LocalMux
    port map (
            O => \N__26035\,
            I => \N__26032\
        );

    \I__3900\ : Span4Mux_v
    port map (
            O => \N__26032\,
            I => \N__26028\
        );

    \I__3899\ : CascadeMux
    port map (
            O => \N__26031\,
            I => \N__26024\
        );

    \I__3898\ : Span4Mux_h
    port map (
            O => \N__26028\,
            I => \N__26021\
        );

    \I__3897\ : InMux
    port map (
            O => \N__26027\,
            I => \N__26016\
        );

    \I__3896\ : InMux
    port map (
            O => \N__26024\,
            I => \N__26016\
        );

    \I__3895\ : Odrv4
    port map (
            O => \N__26021\,
            I => buf_adcdata_iac_17
        );

    \I__3894\ : LocalMux
    port map (
            O => \N__26016\,
            I => buf_adcdata_iac_17
        );

    \I__3893\ : CascadeMux
    port map (
            O => \N__26011\,
            I => \n22201_cascade_\
        );

    \I__3892\ : CascadeMux
    port map (
            O => \N__26008\,
            I => \N__26005\
        );

    \I__3891\ : InMux
    port map (
            O => \N__26005\,
            I => \N__26002\
        );

    \I__3890\ : LocalMux
    port map (
            O => \N__26002\,
            I => \N__25999\
        );

    \I__3889\ : Span4Mux_v
    port map (
            O => \N__25999\,
            I => \N__25996\
        );

    \I__3888\ : Odrv4
    port map (
            O => \N__25996\,
            I => n20805
        );

    \I__3887\ : CascadeMux
    port map (
            O => \N__25993\,
            I => \N__25989\
        );

    \I__3886\ : InMux
    port map (
            O => \N__25992\,
            I => \N__25986\
        );

    \I__3885\ : InMux
    port map (
            O => \N__25989\,
            I => \N__25983\
        );

    \I__3884\ : LocalMux
    port map (
            O => \N__25986\,
            I => \N__25977\
        );

    \I__3883\ : LocalMux
    port map (
            O => \N__25983\,
            I => \N__25977\
        );

    \I__3882\ : InMux
    port map (
            O => \N__25982\,
            I => \N__25974\
        );

    \I__3881\ : Odrv12
    port map (
            O => \N__25977\,
            I => cmd_rdadctmp_24
        );

    \I__3880\ : LocalMux
    port map (
            O => \N__25974\,
            I => cmd_rdadctmp_24
        );

    \I__3879\ : InMux
    port map (
            O => \N__25969\,
            I => \N__25965\
        );

    \I__3878\ : InMux
    port map (
            O => \N__25968\,
            I => \N__25962\
        );

    \I__3877\ : LocalMux
    port map (
            O => \N__25965\,
            I => \N__25958\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__25962\,
            I => \N__25955\
        );

    \I__3875\ : InMux
    port map (
            O => \N__25961\,
            I => \N__25952\
        );

    \I__3874\ : Span4Mux_v
    port map (
            O => \N__25958\,
            I => \N__25949\
        );

    \I__3873\ : Span4Mux_h
    port map (
            O => \N__25955\,
            I => \N__25946\
        );

    \I__3872\ : LocalMux
    port map (
            O => \N__25952\,
            I => buf_adcdata_iac_10
        );

    \I__3871\ : Odrv4
    port map (
            O => \N__25949\,
            I => buf_adcdata_iac_10
        );

    \I__3870\ : Odrv4
    port map (
            O => \N__25946\,
            I => buf_adcdata_iac_10
        );

    \I__3869\ : CascadeMux
    port map (
            O => \N__25939\,
            I => \N__25934\
        );

    \I__3868\ : CascadeMux
    port map (
            O => \N__25938\,
            I => \N__25931\
        );

    \I__3867\ : CascadeMux
    port map (
            O => \N__25937\,
            I => \N__25927\
        );

    \I__3866\ : InMux
    port map (
            O => \N__25934\,
            I => \N__25920\
        );

    \I__3865\ : InMux
    port map (
            O => \N__25931\,
            I => \N__25920\
        );

    \I__3864\ : InMux
    port map (
            O => \N__25930\,
            I => \N__25920\
        );

    \I__3863\ : InMux
    port map (
            O => \N__25927\,
            I => \N__25917\
        );

    \I__3862\ : LocalMux
    port map (
            O => \N__25920\,
            I => \SIG_DDS.bit_cnt_1\
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__25917\,
            I => \SIG_DDS.bit_cnt_1\
        );

    \I__3860\ : InMux
    port map (
            O => \N__25912\,
            I => \N__25905\
        );

    \I__3859\ : InMux
    port map (
            O => \N__25911\,
            I => \N__25905\
        );

    \I__3858\ : InMux
    port map (
            O => \N__25910\,
            I => \N__25902\
        );

    \I__3857\ : LocalMux
    port map (
            O => \N__25905\,
            I => \SIG_DDS.bit_cnt_2\
        );

    \I__3856\ : LocalMux
    port map (
            O => \N__25902\,
            I => \SIG_DDS.bit_cnt_2\
        );

    \I__3855\ : InMux
    port map (
            O => \N__25897\,
            I => \N__25894\
        );

    \I__3854\ : LocalMux
    port map (
            O => \N__25894\,
            I => \N__25890\
        );

    \I__3853\ : InMux
    port map (
            O => \N__25893\,
            I => \N__25886\
        );

    \I__3852\ : Span12Mux_v
    port map (
            O => \N__25890\,
            I => \N__25883\
        );

    \I__3851\ : InMux
    port map (
            O => \N__25889\,
            I => \N__25880\
        );

    \I__3850\ : LocalMux
    port map (
            O => \N__25886\,
            I => buf_adcdata_vac_11
        );

    \I__3849\ : Odrv12
    port map (
            O => \N__25883\,
            I => buf_adcdata_vac_11
        );

    \I__3848\ : LocalMux
    port map (
            O => \N__25880\,
            I => buf_adcdata_vac_11
        );

    \I__3847\ : CascadeMux
    port map (
            O => \N__25873\,
            I => \N__25869\
        );

    \I__3846\ : CascadeMux
    port map (
            O => \N__25872\,
            I => \N__25866\
        );

    \I__3845\ : InMux
    port map (
            O => \N__25869\,
            I => \N__25863\
        );

    \I__3844\ : InMux
    port map (
            O => \N__25866\,
            I => \N__25860\
        );

    \I__3843\ : LocalMux
    port map (
            O => \N__25863\,
            I => \N__25857\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__25860\,
            I => \N__25853\
        );

    \I__3841\ : Span4Mux_h
    port map (
            O => \N__25857\,
            I => \N__25850\
        );

    \I__3840\ : InMux
    port map (
            O => \N__25856\,
            I => \N__25847\
        );

    \I__3839\ : Odrv4
    port map (
            O => \N__25853\,
            I => cmd_rdadctmp_23
        );

    \I__3838\ : Odrv4
    port map (
            O => \N__25850\,
            I => cmd_rdadctmp_23
        );

    \I__3837\ : LocalMux
    port map (
            O => \N__25847\,
            I => cmd_rdadctmp_23
        );

    \I__3836\ : CascadeMux
    port map (
            O => \N__25840\,
            I => \N__25837\
        );

    \I__3835\ : InMux
    port map (
            O => \N__25837\,
            I => \N__25834\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__25834\,
            I => n8
        );

    \I__3833\ : InMux
    port map (
            O => \N__25831\,
            I => \N__25828\
        );

    \I__3832\ : LocalMux
    port map (
            O => \N__25828\,
            I => \N__25825\
        );

    \I__3831\ : Span4Mux_h
    port map (
            O => \N__25825\,
            I => \N__25822\
        );

    \I__3830\ : Odrv4
    port map (
            O => \N__25822\,
            I => n22117
        );

    \I__3829\ : CascadeMux
    port map (
            O => \N__25819\,
            I => \N__25816\
        );

    \I__3828\ : InMux
    port map (
            O => \N__25816\,
            I => \N__25813\
        );

    \I__3827\ : LocalMux
    port map (
            O => \N__25813\,
            I => \N__25809\
        );

    \I__3826\ : InMux
    port map (
            O => \N__25812\,
            I => \N__25805\
        );

    \I__3825\ : Span4Mux_h
    port map (
            O => \N__25809\,
            I => \N__25802\
        );

    \I__3824\ : InMux
    port map (
            O => \N__25808\,
            I => \N__25799\
        );

    \I__3823\ : LocalMux
    port map (
            O => \N__25805\,
            I => \N__25796\
        );

    \I__3822\ : Span4Mux_h
    port map (
            O => \N__25802\,
            I => \N__25793\
        );

    \I__3821\ : LocalMux
    port map (
            O => \N__25799\,
            I => buf_adcdata_iac_13
        );

    \I__3820\ : Odrv4
    port map (
            O => \N__25796\,
            I => buf_adcdata_iac_13
        );

    \I__3819\ : Odrv4
    port map (
            O => \N__25793\,
            I => buf_adcdata_iac_13
        );

    \I__3818\ : InMux
    port map (
            O => \N__25786\,
            I => \N__25782\
        );

    \I__3817\ : InMux
    port map (
            O => \N__25785\,
            I => \N__25779\
        );

    \I__3816\ : LocalMux
    port map (
            O => \N__25782\,
            I => \SIG_DDS.bit_cnt_3\
        );

    \I__3815\ : LocalMux
    port map (
            O => \N__25779\,
            I => \SIG_DDS.bit_cnt_3\
        );

    \I__3814\ : InMux
    port map (
            O => \N__25774\,
            I => \N__25771\
        );

    \I__3813\ : LocalMux
    port map (
            O => \N__25771\,
            I => \N__25768\
        );

    \I__3812\ : Odrv12
    port map (
            O => \N__25768\,
            I => \SIG_DDS.n21292\
        );

    \I__3811\ : CascadeMux
    port map (
            O => \N__25765\,
            I => \n20624_cascade_\
        );

    \I__3810\ : CascadeMux
    port map (
            O => \N__25762\,
            I => \SIG_DDS.n10_cascade_\
        );

    \I__3809\ : CascadeMux
    port map (
            O => \N__25759\,
            I => \N__25756\
        );

    \I__3808\ : InMux
    port map (
            O => \N__25756\,
            I => \N__25753\
        );

    \I__3807\ : LocalMux
    port map (
            O => \N__25753\,
            I => \N__25750\
        );

    \I__3806\ : Span4Mux_v
    port map (
            O => \N__25750\,
            I => \N__25747\
        );

    \I__3805\ : Span4Mux_h
    port map (
            O => \N__25747\,
            I => \N__25743\
        );

    \I__3804\ : CascadeMux
    port map (
            O => \N__25746\,
            I => \N__25740\
        );

    \I__3803\ : Span4Mux_v
    port map (
            O => \N__25743\,
            I => \N__25737\
        );

    \I__3802\ : InMux
    port map (
            O => \N__25740\,
            I => \N__25734\
        );

    \I__3801\ : Odrv4
    port map (
            O => \N__25737\,
            I => \buf_readRTD_12\
        );

    \I__3800\ : LocalMux
    port map (
            O => \N__25734\,
            I => \buf_readRTD_12\
        );

    \I__3799\ : InMux
    port map (
            O => \N__25729\,
            I => \N__25726\
        );

    \I__3798\ : LocalMux
    port map (
            O => \N__25726\,
            I => n22006
        );

    \I__3797\ : CascadeMux
    port map (
            O => \N__25723\,
            I => \n22027_cascade_\
        );

    \I__3796\ : InMux
    port map (
            O => \N__25720\,
            I => \N__25717\
        );

    \I__3795\ : LocalMux
    port map (
            O => \N__25717\,
            I => \N__25714\
        );

    \I__3794\ : Odrv4
    port map (
            O => \N__25714\,
            I => n22030
        );

    \I__3793\ : InMux
    port map (
            O => \N__25711\,
            I => \N__25707\
        );

    \I__3792\ : InMux
    port map (
            O => \N__25710\,
            I => \N__25703\
        );

    \I__3791\ : LocalMux
    port map (
            O => \N__25707\,
            I => \N__25700\
        );

    \I__3790\ : CascadeMux
    port map (
            O => \N__25706\,
            I => \N__25697\
        );

    \I__3789\ : LocalMux
    port map (
            O => \N__25703\,
            I => \N__25694\
        );

    \I__3788\ : Span4Mux_v
    port map (
            O => \N__25700\,
            I => \N__25691\
        );

    \I__3787\ : InMux
    port map (
            O => \N__25697\,
            I => \N__25688\
        );

    \I__3786\ : Span4Mux_h
    port map (
            O => \N__25694\,
            I => \N__25685\
        );

    \I__3785\ : Span4Mux_v
    port map (
            O => \N__25691\,
            I => \N__25682\
        );

    \I__3784\ : LocalMux
    port map (
            O => \N__25688\,
            I => buf_adcdata_vac_20
        );

    \I__3783\ : Odrv4
    port map (
            O => \N__25685\,
            I => buf_adcdata_vac_20
        );

    \I__3782\ : Odrv4
    port map (
            O => \N__25682\,
            I => buf_adcdata_vac_20
        );

    \I__3781\ : CascadeMux
    port map (
            O => \N__25675\,
            I => \N__25672\
        );

    \I__3780\ : InMux
    port map (
            O => \N__25672\,
            I => \N__25669\
        );

    \I__3779\ : LocalMux
    port map (
            O => \N__25669\,
            I => \N__25665\
        );

    \I__3778\ : CascadeMux
    port map (
            O => \N__25668\,
            I => \N__25662\
        );

    \I__3777\ : Span4Mux_v
    port map (
            O => \N__25665\,
            I => \N__25659\
        );

    \I__3776\ : InMux
    port map (
            O => \N__25662\,
            I => \N__25656\
        );

    \I__3775\ : Odrv4
    port map (
            O => \N__25659\,
            I => buf_adcdata_vdc_20
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__25656\,
            I => buf_adcdata_vdc_20
        );

    \I__3773\ : InMux
    port map (
            O => \N__25651\,
            I => \N__25648\
        );

    \I__3772\ : LocalMux
    port map (
            O => \N__25648\,
            I => n22207
        );

    \I__3771\ : InMux
    port map (
            O => \N__25645\,
            I => \N__25642\
        );

    \I__3770\ : LocalMux
    port map (
            O => \N__25642\,
            I => n20801
        );

    \I__3769\ : InMux
    port map (
            O => \N__25639\,
            I => \N__25636\
        );

    \I__3768\ : LocalMux
    port map (
            O => \N__25636\,
            I => \N__25633\
        );

    \I__3767\ : Span4Mux_h
    port map (
            O => \N__25633\,
            I => \N__25630\
        );

    \I__3766\ : Span4Mux_h
    port map (
            O => \N__25630\,
            I => \N__25627\
        );

    \I__3765\ : Odrv4
    port map (
            O => \N__25627\,
            I => buf_data_iac_17
        );

    \I__3764\ : CascadeMux
    port map (
            O => \N__25624\,
            I => \n20818_cascade_\
        );

    \I__3763\ : InMux
    port map (
            O => \N__25621\,
            I => \N__25618\
        );

    \I__3762\ : LocalMux
    port map (
            O => \N__25618\,
            I => n20871
        );

    \I__3761\ : CascadeMux
    port map (
            O => \N__25615\,
            I => \n20820_cascade_\
        );

    \I__3760\ : InMux
    port map (
            O => \N__25612\,
            I => \N__25609\
        );

    \I__3759\ : LocalMux
    port map (
            O => \N__25609\,
            I => n21967
        );

    \I__3758\ : InMux
    port map (
            O => \N__25606\,
            I => \N__25603\
        );

    \I__3757\ : LocalMux
    port map (
            O => \N__25603\,
            I => n21970
        );

    \I__3756\ : CascadeMux
    port map (
            O => \N__25600\,
            I => \n22003_cascade_\
        );

    \I__3755\ : InMux
    port map (
            O => \N__25597\,
            I => \N__25594\
        );

    \I__3754\ : LocalMux
    port map (
            O => \N__25594\,
            I => \N__25591\
        );

    \I__3753\ : Odrv4
    port map (
            O => \N__25591\,
            I => n22060
        );

    \I__3752\ : InMux
    port map (
            O => \N__25588\,
            I => \N__25585\
        );

    \I__3751\ : LocalMux
    port map (
            O => \N__25585\,
            I => n22054
        );

    \I__3750\ : CascadeMux
    port map (
            O => \N__25582\,
            I => \n22015_cascade_\
        );

    \I__3749\ : InMux
    port map (
            O => \N__25579\,
            I => \N__25575\
        );

    \I__3748\ : InMux
    port map (
            O => \N__25578\,
            I => \N__25572\
        );

    \I__3747\ : LocalMux
    port map (
            O => \N__25575\,
            I => cmd_rdadcbuf_28
        );

    \I__3746\ : LocalMux
    port map (
            O => \N__25572\,
            I => cmd_rdadcbuf_28
        );

    \I__3745\ : InMux
    port map (
            O => \N__25567\,
            I => \ADC_VDC.n19391\
        );

    \I__3744\ : InMux
    port map (
            O => \N__25564\,
            I => \N__25560\
        );

    \I__3743\ : InMux
    port map (
            O => \N__25563\,
            I => \N__25557\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__25560\,
            I => cmd_rdadcbuf_29
        );

    \I__3741\ : LocalMux
    port map (
            O => \N__25557\,
            I => cmd_rdadcbuf_29
        );

    \I__3740\ : InMux
    port map (
            O => \N__25552\,
            I => \ADC_VDC.n19392\
        );

    \I__3739\ : InMux
    port map (
            O => \N__25549\,
            I => \N__25545\
        );

    \I__3738\ : InMux
    port map (
            O => \N__25548\,
            I => \N__25542\
        );

    \I__3737\ : LocalMux
    port map (
            O => \N__25545\,
            I => cmd_rdadcbuf_30
        );

    \I__3736\ : LocalMux
    port map (
            O => \N__25542\,
            I => cmd_rdadcbuf_30
        );

    \I__3735\ : InMux
    port map (
            O => \N__25537\,
            I => \ADC_VDC.n19393\
        );

    \I__3734\ : InMux
    port map (
            O => \N__25534\,
            I => \N__25530\
        );

    \I__3733\ : InMux
    port map (
            O => \N__25533\,
            I => \N__25527\
        );

    \I__3732\ : LocalMux
    port map (
            O => \N__25530\,
            I => cmd_rdadcbuf_31
        );

    \I__3731\ : LocalMux
    port map (
            O => \N__25527\,
            I => cmd_rdadcbuf_31
        );

    \I__3730\ : InMux
    port map (
            O => \N__25522\,
            I => \ADC_VDC.n19394\
        );

    \I__3729\ : InMux
    port map (
            O => \N__25519\,
            I => \N__25515\
        );

    \I__3728\ : InMux
    port map (
            O => \N__25518\,
            I => \N__25512\
        );

    \I__3727\ : LocalMux
    port map (
            O => \N__25515\,
            I => cmd_rdadcbuf_32
        );

    \I__3726\ : LocalMux
    port map (
            O => \N__25512\,
            I => cmd_rdadcbuf_32
        );

    \I__3725\ : InMux
    port map (
            O => \N__25507\,
            I => \bfn_9_9_0_\
        );

    \I__3724\ : InMux
    port map (
            O => \N__25504\,
            I => \N__25500\
        );

    \I__3723\ : InMux
    port map (
            O => \N__25503\,
            I => \N__25497\
        );

    \I__3722\ : LocalMux
    port map (
            O => \N__25500\,
            I => cmd_rdadcbuf_33
        );

    \I__3721\ : LocalMux
    port map (
            O => \N__25497\,
            I => cmd_rdadcbuf_33
        );

    \I__3720\ : InMux
    port map (
            O => \N__25492\,
            I => \ADC_VDC.n19396\
        );

    \I__3719\ : InMux
    port map (
            O => \N__25489\,
            I => \ADC_VDC.n19397\
        );

    \I__3718\ : InMux
    port map (
            O => \N__25486\,
            I => \N__25483\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__25483\,
            I => \N__25480\
        );

    \I__3716\ : Odrv4
    port map (
            O => \N__25480\,
            I => n20772
        );

    \I__3715\ : InMux
    port map (
            O => \N__25477\,
            I => \N__25474\
        );

    \I__3714\ : LocalMux
    port map (
            O => \N__25474\,
            I => n21943
        );

    \I__3713\ : CascadeMux
    port map (
            O => \N__25471\,
            I => \n21946_cascade_\
        );

    \I__3712\ : InMux
    port map (
            O => \N__25468\,
            I => \ADC_VDC.n19383\
        );

    \I__3711\ : CascadeMux
    port map (
            O => \N__25465\,
            I => \N__25460\
        );

    \I__3710\ : InMux
    port map (
            O => \N__25464\,
            I => \N__25457\
        );

    \I__3709\ : InMux
    port map (
            O => \N__25463\,
            I => \N__25454\
        );

    \I__3708\ : InMux
    port map (
            O => \N__25460\,
            I => \N__25451\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__25457\,
            I => cmd_rdadctmp_21_adj_1451
        );

    \I__3706\ : LocalMux
    port map (
            O => \N__25454\,
            I => cmd_rdadctmp_21_adj_1451
        );

    \I__3705\ : LocalMux
    port map (
            O => \N__25451\,
            I => cmd_rdadctmp_21_adj_1451
        );

    \I__3704\ : InMux
    port map (
            O => \N__25444\,
            I => \N__25440\
        );

    \I__3703\ : InMux
    port map (
            O => \N__25443\,
            I => \N__25437\
        );

    \I__3702\ : LocalMux
    port map (
            O => \N__25440\,
            I => cmd_rdadcbuf_21
        );

    \I__3701\ : LocalMux
    port map (
            O => \N__25437\,
            I => cmd_rdadcbuf_21
        );

    \I__3700\ : InMux
    port map (
            O => \N__25432\,
            I => \ADC_VDC.n19384\
        );

    \I__3699\ : InMux
    port map (
            O => \N__25429\,
            I => \N__25425\
        );

    \I__3698\ : CascadeMux
    port map (
            O => \N__25428\,
            I => \N__25421\
        );

    \I__3697\ : LocalMux
    port map (
            O => \N__25425\,
            I => \N__25418\
        );

    \I__3696\ : InMux
    port map (
            O => \N__25424\,
            I => \N__25415\
        );

    \I__3695\ : InMux
    port map (
            O => \N__25421\,
            I => \N__25412\
        );

    \I__3694\ : Odrv4
    port map (
            O => \N__25418\,
            I => cmd_rdadctmp_22_adj_1450
        );

    \I__3693\ : LocalMux
    port map (
            O => \N__25415\,
            I => cmd_rdadctmp_22_adj_1450
        );

    \I__3692\ : LocalMux
    port map (
            O => \N__25412\,
            I => cmd_rdadctmp_22_adj_1450
        );

    \I__3691\ : InMux
    port map (
            O => \N__25405\,
            I => \ADC_VDC.n19385\
        );

    \I__3690\ : CascadeMux
    port map (
            O => \N__25402\,
            I => \N__25398\
        );

    \I__3689\ : CascadeMux
    port map (
            O => \N__25401\,
            I => \N__25395\
        );

    \I__3688\ : InMux
    port map (
            O => \N__25398\,
            I => \N__25392\
        );

    \I__3687\ : InMux
    port map (
            O => \N__25395\,
            I => \N__25389\
        );

    \I__3686\ : LocalMux
    port map (
            O => \N__25392\,
            I => \N__25386\
        );

    \I__3685\ : LocalMux
    port map (
            O => \N__25389\,
            I => \ADC_VDC.cmd_rdadctmp_23\
        );

    \I__3684\ : Odrv4
    port map (
            O => \N__25386\,
            I => \ADC_VDC.cmd_rdadctmp_23\
        );

    \I__3683\ : InMux
    port map (
            O => \N__25381\,
            I => \ADC_VDC.n19386\
        );

    \I__3682\ : InMux
    port map (
            O => \N__25378\,
            I => \N__25374\
        );

    \I__3681\ : InMux
    port map (
            O => \N__25377\,
            I => \N__25371\
        );

    \I__3680\ : LocalMux
    port map (
            O => \N__25374\,
            I => cmd_rdadcbuf_24
        );

    \I__3679\ : LocalMux
    port map (
            O => \N__25371\,
            I => cmd_rdadcbuf_24
        );

    \I__3678\ : InMux
    port map (
            O => \N__25366\,
            I => \bfn_9_8_0_\
        );

    \I__3677\ : InMux
    port map (
            O => \N__25363\,
            I => \N__25359\
        );

    \I__3676\ : InMux
    port map (
            O => \N__25362\,
            I => \N__25356\
        );

    \I__3675\ : LocalMux
    port map (
            O => \N__25359\,
            I => cmd_rdadcbuf_25
        );

    \I__3674\ : LocalMux
    port map (
            O => \N__25356\,
            I => cmd_rdadcbuf_25
        );

    \I__3673\ : InMux
    port map (
            O => \N__25351\,
            I => \ADC_VDC.n19388\
        );

    \I__3672\ : InMux
    port map (
            O => \N__25348\,
            I => \N__25344\
        );

    \I__3671\ : InMux
    port map (
            O => \N__25347\,
            I => \N__25341\
        );

    \I__3670\ : LocalMux
    port map (
            O => \N__25344\,
            I => cmd_rdadcbuf_26
        );

    \I__3669\ : LocalMux
    port map (
            O => \N__25341\,
            I => cmd_rdadcbuf_26
        );

    \I__3668\ : InMux
    port map (
            O => \N__25336\,
            I => \ADC_VDC.n19389\
        );

    \I__3667\ : InMux
    port map (
            O => \N__25333\,
            I => \N__25329\
        );

    \I__3666\ : InMux
    port map (
            O => \N__25332\,
            I => \N__25326\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__25329\,
            I => cmd_rdadcbuf_27
        );

    \I__3664\ : LocalMux
    port map (
            O => \N__25326\,
            I => cmd_rdadcbuf_27
        );

    \I__3663\ : InMux
    port map (
            O => \N__25321\,
            I => \ADC_VDC.n19390\
        );

    \I__3662\ : InMux
    port map (
            O => \N__25318\,
            I => \N__25314\
        );

    \I__3661\ : InMux
    port map (
            O => \N__25317\,
            I => \N__25311\
        );

    \I__3660\ : LocalMux
    port map (
            O => \N__25314\,
            I => cmd_rdadcbuf_11
        );

    \I__3659\ : LocalMux
    port map (
            O => \N__25311\,
            I => cmd_rdadcbuf_11
        );

    \I__3658\ : InMux
    port map (
            O => \N__25306\,
            I => \ADC_VDC.n19374\
        );

    \I__3657\ : InMux
    port map (
            O => \N__25303\,
            I => \N__25299\
        );

    \I__3656\ : InMux
    port map (
            O => \N__25302\,
            I => \N__25296\
        );

    \I__3655\ : LocalMux
    port map (
            O => \N__25299\,
            I => cmd_rdadcbuf_12
        );

    \I__3654\ : LocalMux
    port map (
            O => \N__25296\,
            I => cmd_rdadcbuf_12
        );

    \I__3653\ : InMux
    port map (
            O => \N__25291\,
            I => \ADC_VDC.n19375\
        );

    \I__3652\ : CascadeMux
    port map (
            O => \N__25288\,
            I => \N__25283\
        );

    \I__3651\ : InMux
    port map (
            O => \N__25287\,
            I => \N__25278\
        );

    \I__3650\ : InMux
    port map (
            O => \N__25286\,
            I => \N__25278\
        );

    \I__3649\ : InMux
    port map (
            O => \N__25283\,
            I => \N__25275\
        );

    \I__3648\ : LocalMux
    port map (
            O => \N__25278\,
            I => cmd_rdadctmp_13_adj_1459
        );

    \I__3647\ : LocalMux
    port map (
            O => \N__25275\,
            I => cmd_rdadctmp_13_adj_1459
        );

    \I__3646\ : InMux
    port map (
            O => \N__25270\,
            I => \N__25267\
        );

    \I__3645\ : LocalMux
    port map (
            O => \N__25267\,
            I => \N__25263\
        );

    \I__3644\ : InMux
    port map (
            O => \N__25266\,
            I => \N__25260\
        );

    \I__3643\ : Odrv4
    port map (
            O => \N__25263\,
            I => cmd_rdadcbuf_13
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__25260\,
            I => cmd_rdadcbuf_13
        );

    \I__3641\ : InMux
    port map (
            O => \N__25255\,
            I => \ADC_VDC.n19376\
        );

    \I__3640\ : CascadeMux
    port map (
            O => \N__25252\,
            I => \N__25249\
        );

    \I__3639\ : InMux
    port map (
            O => \N__25249\,
            I => \N__25244\
        );

    \I__3638\ : CascadeMux
    port map (
            O => \N__25248\,
            I => \N__25241\
        );

    \I__3637\ : CascadeMux
    port map (
            O => \N__25247\,
            I => \N__25238\
        );

    \I__3636\ : LocalMux
    port map (
            O => \N__25244\,
            I => \N__25235\
        );

    \I__3635\ : InMux
    port map (
            O => \N__25241\,
            I => \N__25232\
        );

    \I__3634\ : InMux
    port map (
            O => \N__25238\,
            I => \N__25229\
        );

    \I__3633\ : Odrv4
    port map (
            O => \N__25235\,
            I => cmd_rdadctmp_14_adj_1458
        );

    \I__3632\ : LocalMux
    port map (
            O => \N__25232\,
            I => cmd_rdadctmp_14_adj_1458
        );

    \I__3631\ : LocalMux
    port map (
            O => \N__25229\,
            I => cmd_rdadctmp_14_adj_1458
        );

    \I__3630\ : InMux
    port map (
            O => \N__25222\,
            I => \N__25218\
        );

    \I__3629\ : InMux
    port map (
            O => \N__25221\,
            I => \N__25215\
        );

    \I__3628\ : LocalMux
    port map (
            O => \N__25218\,
            I => cmd_rdadcbuf_14
        );

    \I__3627\ : LocalMux
    port map (
            O => \N__25215\,
            I => cmd_rdadcbuf_14
        );

    \I__3626\ : InMux
    port map (
            O => \N__25210\,
            I => \ADC_VDC.n19377\
        );

    \I__3625\ : InMux
    port map (
            O => \N__25207\,
            I => \ADC_VDC.n19378\
        );

    \I__3624\ : InMux
    port map (
            O => \N__25204\,
            I => \bfn_9_7_0_\
        );

    \I__3623\ : InMux
    port map (
            O => \N__25201\,
            I => \ADC_VDC.n19380\
        );

    \I__3622\ : CascadeMux
    port map (
            O => \N__25198\,
            I => \N__25194\
        );

    \I__3621\ : CascadeMux
    port map (
            O => \N__25197\,
            I => \N__25190\
        );

    \I__3620\ : InMux
    port map (
            O => \N__25194\,
            I => \N__25187\
        );

    \I__3619\ : InMux
    port map (
            O => \N__25193\,
            I => \N__25184\
        );

    \I__3618\ : InMux
    port map (
            O => \N__25190\,
            I => \N__25181\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__25187\,
            I => cmd_rdadctmp_18_adj_1454
        );

    \I__3616\ : LocalMux
    port map (
            O => \N__25184\,
            I => cmd_rdadctmp_18_adj_1454
        );

    \I__3615\ : LocalMux
    port map (
            O => \N__25181\,
            I => cmd_rdadctmp_18_adj_1454
        );

    \I__3614\ : InMux
    port map (
            O => \N__25174\,
            I => \ADC_VDC.n19381\
        );

    \I__3613\ : InMux
    port map (
            O => \N__25171\,
            I => \ADC_VDC.n19382\
        );

    \I__3612\ : InMux
    port map (
            O => \N__25168\,
            I => \N__25165\
        );

    \I__3611\ : LocalMux
    port map (
            O => \N__25165\,
            I => \ADC_VDC.cmd_rdadcbuf_3\
        );

    \I__3610\ : InMux
    port map (
            O => \N__25162\,
            I => \ADC_VDC.n19366\
        );

    \I__3609\ : InMux
    port map (
            O => \N__25159\,
            I => \N__25156\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__25156\,
            I => \ADC_VDC.cmd_rdadcbuf_4\
        );

    \I__3607\ : InMux
    port map (
            O => \N__25153\,
            I => \ADC_VDC.n19367\
        );

    \I__3606\ : CascadeMux
    port map (
            O => \N__25150\,
            I => \N__25145\
        );

    \I__3605\ : InMux
    port map (
            O => \N__25149\,
            I => \N__25140\
        );

    \I__3604\ : InMux
    port map (
            O => \N__25148\,
            I => \N__25140\
        );

    \I__3603\ : InMux
    port map (
            O => \N__25145\,
            I => \N__25137\
        );

    \I__3602\ : LocalMux
    port map (
            O => \N__25140\,
            I => cmd_rdadctmp_5_adj_1467
        );

    \I__3601\ : LocalMux
    port map (
            O => \N__25137\,
            I => cmd_rdadctmp_5_adj_1467
        );

    \I__3600\ : InMux
    port map (
            O => \N__25132\,
            I => \N__25129\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__25129\,
            I => \ADC_VDC.cmd_rdadcbuf_5\
        );

    \I__3598\ : InMux
    port map (
            O => \N__25126\,
            I => \ADC_VDC.n19368\
        );

    \I__3597\ : CascadeMux
    port map (
            O => \N__25123\,
            I => \N__25118\
        );

    \I__3596\ : InMux
    port map (
            O => \N__25122\,
            I => \N__25113\
        );

    \I__3595\ : InMux
    port map (
            O => \N__25121\,
            I => \N__25113\
        );

    \I__3594\ : InMux
    port map (
            O => \N__25118\,
            I => \N__25110\
        );

    \I__3593\ : LocalMux
    port map (
            O => \N__25113\,
            I => cmd_rdadctmp_6_adj_1466
        );

    \I__3592\ : LocalMux
    port map (
            O => \N__25110\,
            I => cmd_rdadctmp_6_adj_1466
        );

    \I__3591\ : InMux
    port map (
            O => \N__25105\,
            I => \N__25102\
        );

    \I__3590\ : LocalMux
    port map (
            O => \N__25102\,
            I => \ADC_VDC.cmd_rdadcbuf_6\
        );

    \I__3589\ : InMux
    port map (
            O => \N__25099\,
            I => \ADC_VDC.n19369\
        );

    \I__3588\ : InMux
    port map (
            O => \N__25096\,
            I => \N__25093\
        );

    \I__3587\ : LocalMux
    port map (
            O => \N__25093\,
            I => \ADC_VDC.cmd_rdadcbuf_7\
        );

    \I__3586\ : InMux
    port map (
            O => \N__25090\,
            I => \ADC_VDC.n19370\
        );

    \I__3585\ : InMux
    port map (
            O => \N__25087\,
            I => \N__25084\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__25084\,
            I => \ADC_VDC.cmd_rdadcbuf_8\
        );

    \I__3583\ : InMux
    port map (
            O => \N__25081\,
            I => \bfn_9_6_0_\
        );

    \I__3582\ : InMux
    port map (
            O => \N__25078\,
            I => \N__25071\
        );

    \I__3581\ : InMux
    port map (
            O => \N__25077\,
            I => \N__25071\
        );

    \I__3580\ : InMux
    port map (
            O => \N__25076\,
            I => \N__25068\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__25071\,
            I => cmd_rdadctmp_9_adj_1463
        );

    \I__3578\ : LocalMux
    port map (
            O => \N__25068\,
            I => cmd_rdadctmp_9_adj_1463
        );

    \I__3577\ : CascadeMux
    port map (
            O => \N__25063\,
            I => \N__25060\
        );

    \I__3576\ : InMux
    port map (
            O => \N__25060\,
            I => \N__25057\
        );

    \I__3575\ : LocalMux
    port map (
            O => \N__25057\,
            I => \ADC_VDC.cmd_rdadcbuf_9\
        );

    \I__3574\ : InMux
    port map (
            O => \N__25054\,
            I => \ADC_VDC.n19372\
        );

    \I__3573\ : InMux
    port map (
            O => \N__25051\,
            I => \N__25048\
        );

    \I__3572\ : LocalMux
    port map (
            O => \N__25048\,
            I => \ADC_VDC.cmd_rdadcbuf_10\
        );

    \I__3571\ : InMux
    port map (
            O => \N__25045\,
            I => \ADC_VDC.n19373\
        );

    \I__3570\ : InMux
    port map (
            O => \N__25042\,
            I => \N__25038\
        );

    \I__3569\ : InMux
    port map (
            O => \N__25041\,
            I => \N__25035\
        );

    \I__3568\ : LocalMux
    port map (
            O => \N__25038\,
            I => \N__25032\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__25035\,
            I => \ADC_IAC.bit_cnt_5\
        );

    \I__3566\ : Odrv4
    port map (
            O => \N__25032\,
            I => \ADC_IAC.bit_cnt_5\
        );

    \I__3565\ : CascadeMux
    port map (
            O => \N__25027\,
            I => \ADC_IAC.n20765_cascade_\
        );

    \I__3564\ : CascadeMux
    port map (
            O => \N__25024\,
            I => \ADC_IAC.n21007_cascade_\
        );

    \I__3563\ : CEMux
    port map (
            O => \N__25021\,
            I => \N__25018\
        );

    \I__3562\ : LocalMux
    port map (
            O => \N__25018\,
            I => \N__25015\
        );

    \I__3561\ : Odrv4
    port map (
            O => \N__25015\,
            I => \ADC_IAC.n20670\
        );

    \I__3560\ : CascadeMux
    port map (
            O => \N__25012\,
            I => \N__25009\
        );

    \I__3559\ : InMux
    port map (
            O => \N__25009\,
            I => \N__25004\
        );

    \I__3558\ : InMux
    port map (
            O => \N__25008\,
            I => \N__25001\
        );

    \I__3557\ : InMux
    port map (
            O => \N__25007\,
            I => \N__24998\
        );

    \I__3556\ : LocalMux
    port map (
            O => \N__25004\,
            I => \N__24990\
        );

    \I__3555\ : LocalMux
    port map (
            O => \N__25001\,
            I => \N__24990\
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__24998\,
            I => \N__24990\
        );

    \I__3553\ : CascadeMux
    port map (
            O => \N__24997\,
            I => \N__24986\
        );

    \I__3552\ : Span4Mux_h
    port map (
            O => \N__24990\,
            I => \N__24983\
        );

    \I__3551\ : InMux
    port map (
            O => \N__24989\,
            I => \N__24978\
        );

    \I__3550\ : InMux
    port map (
            O => \N__24986\,
            I => \N__24978\
        );

    \I__3549\ : Span4Mux_v
    port map (
            O => \N__24983\,
            I => \N__24975\
        );

    \I__3548\ : LocalMux
    port map (
            O => \N__24978\,
            I => \N__24972\
        );

    \I__3547\ : Span4Mux_v
    port map (
            O => \N__24975\,
            I => \N__24969\
        );

    \I__3546\ : Span12Mux_h
    port map (
            O => \N__24972\,
            I => \N__24966\
        );

    \I__3545\ : Span4Mux_h
    port map (
            O => \N__24969\,
            I => \N__24963\
        );

    \I__3544\ : Odrv12
    port map (
            O => \N__24966\,
            I => \IAC_DRDY\
        );

    \I__3543\ : Odrv4
    port map (
            O => \N__24963\,
            I => \IAC_DRDY\
        );

    \I__3542\ : CascadeMux
    port map (
            O => \N__24958\,
            I => \ADC_IAC.n17_cascade_\
        );

    \I__3541\ : CEMux
    port map (
            O => \N__24955\,
            I => \N__24952\
        );

    \I__3540\ : LocalMux
    port map (
            O => \N__24952\,
            I => \N__24949\
        );

    \I__3539\ : Odrv4
    port map (
            O => \N__24949\,
            I => \ADC_IAC.n12\
        );

    \I__3538\ : SRMux
    port map (
            O => \N__24946\,
            I => \N__24943\
        );

    \I__3537\ : LocalMux
    port map (
            O => \N__24943\,
            I => \N__24940\
        );

    \I__3536\ : Span4Mux_h
    port map (
            O => \N__24940\,
            I => \N__24937\
        );

    \I__3535\ : Span4Mux_h
    port map (
            O => \N__24937\,
            I => \N__24934\
        );

    \I__3534\ : Odrv4
    port map (
            O => \N__24934\,
            I => \ADC_VDC.n20345\
        );

    \I__3533\ : InMux
    port map (
            O => \N__24931\,
            I => \N__24928\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__24928\,
            I => \ADC_VDC.cmd_rdadcbuf_0\
        );

    \I__3531\ : InMux
    port map (
            O => \N__24925\,
            I => \N__24922\
        );

    \I__3530\ : LocalMux
    port map (
            O => \N__24922\,
            I => \ADC_VDC.cmd_rdadcbuf_1\
        );

    \I__3529\ : InMux
    port map (
            O => \N__24919\,
            I => \ADC_VDC.n19364\
        );

    \I__3528\ : CascadeMux
    port map (
            O => \N__24916\,
            I => \N__24913\
        );

    \I__3527\ : InMux
    port map (
            O => \N__24913\,
            I => \N__24910\
        );

    \I__3526\ : LocalMux
    port map (
            O => \N__24910\,
            I => \ADC_VDC.cmd_rdadcbuf_2\
        );

    \I__3525\ : InMux
    port map (
            O => \N__24907\,
            I => \ADC_VDC.n19365\
        );

    \I__3524\ : CascadeMux
    port map (
            O => \N__24904\,
            I => \N__24900\
        );

    \I__3523\ : InMux
    port map (
            O => \N__24903\,
            I => \N__24896\
        );

    \I__3522\ : InMux
    port map (
            O => \N__24900\,
            I => \N__24891\
        );

    \I__3521\ : InMux
    port map (
            O => \N__24899\,
            I => \N__24891\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__24896\,
            I => cmd_rdadctmp_30
        );

    \I__3519\ : LocalMux
    port map (
            O => \N__24891\,
            I => cmd_rdadctmp_30
        );

    \I__3518\ : InMux
    port map (
            O => \N__24886\,
            I => \N__24882\
        );

    \I__3517\ : InMux
    port map (
            O => \N__24885\,
            I => \N__24879\
        );

    \I__3516\ : LocalMux
    port map (
            O => \N__24882\,
            I => cmd_rdadctmp_4
        );

    \I__3515\ : LocalMux
    port map (
            O => \N__24879\,
            I => cmd_rdadctmp_4
        );

    \I__3514\ : CascadeMux
    port map (
            O => \N__24874\,
            I => \N__24871\
        );

    \I__3513\ : InMux
    port map (
            O => \N__24871\,
            I => \N__24867\
        );

    \I__3512\ : InMux
    port map (
            O => \N__24870\,
            I => \N__24864\
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__24867\,
            I => cmd_rdadctmp_2
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__24864\,
            I => cmd_rdadctmp_2
        );

    \I__3509\ : CascadeMux
    port map (
            O => \N__24859\,
            I => \N__24856\
        );

    \I__3508\ : InMux
    port map (
            O => \N__24856\,
            I => \N__24850\
        );

    \I__3507\ : InMux
    port map (
            O => \N__24855\,
            I => \N__24850\
        );

    \I__3506\ : LocalMux
    port map (
            O => \N__24850\,
            I => cmd_rdadctmp_3
        );

    \I__3505\ : IoInMux
    port map (
            O => \N__24847\,
            I => \N__24844\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__24844\,
            I => \N__24841\
        );

    \I__3503\ : Span4Mux_s0_v
    port map (
            O => \N__24841\,
            I => \N__24838\
        );

    \I__3502\ : Sp12to4
    port map (
            O => \N__24838\,
            I => \N__24834\
        );

    \I__3501\ : CascadeMux
    port map (
            O => \N__24837\,
            I => \N__24831\
        );

    \I__3500\ : Span12Mux_s11_h
    port map (
            O => \N__24834\,
            I => \N__24828\
        );

    \I__3499\ : InMux
    port map (
            O => \N__24831\,
            I => \N__24825\
        );

    \I__3498\ : Odrv12
    port map (
            O => \N__24828\,
            I => \IAC_CS\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__24825\,
            I => \IAC_CS\
        );

    \I__3496\ : InMux
    port map (
            O => \N__24820\,
            I => \N__24817\
        );

    \I__3495\ : LocalMux
    port map (
            O => \N__24817\,
            I => n14_adj_1581
        );

    \I__3494\ : InMux
    port map (
            O => \N__24814\,
            I => \N__24811\
        );

    \I__3493\ : LocalMux
    port map (
            O => \N__24811\,
            I => \ADC_IAC.n20669\
        );

    \I__3492\ : InMux
    port map (
            O => \N__24808\,
            I => \N__24804\
        );

    \I__3491\ : InMux
    port map (
            O => \N__24807\,
            I => \N__24801\
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__24804\,
            I => \ADC_IAC.bit_cnt_4\
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__24801\,
            I => \ADC_IAC.bit_cnt_4\
        );

    \I__3488\ : InMux
    port map (
            O => \N__24796\,
            I => \N__24792\
        );

    \I__3487\ : InMux
    port map (
            O => \N__24795\,
            I => \N__24789\
        );

    \I__3486\ : LocalMux
    port map (
            O => \N__24792\,
            I => \ADC_IAC.bit_cnt_3\
        );

    \I__3485\ : LocalMux
    port map (
            O => \N__24789\,
            I => \ADC_IAC.bit_cnt_3\
        );

    \I__3484\ : CascadeMux
    port map (
            O => \N__24784\,
            I => \N__24780\
        );

    \I__3483\ : InMux
    port map (
            O => \N__24783\,
            I => \N__24777\
        );

    \I__3482\ : InMux
    port map (
            O => \N__24780\,
            I => \N__24774\
        );

    \I__3481\ : LocalMux
    port map (
            O => \N__24777\,
            I => \ADC_IAC.bit_cnt_1\
        );

    \I__3480\ : LocalMux
    port map (
            O => \N__24774\,
            I => \ADC_IAC.bit_cnt_1\
        );

    \I__3479\ : InMux
    port map (
            O => \N__24769\,
            I => \N__24765\
        );

    \I__3478\ : InMux
    port map (
            O => \N__24768\,
            I => \N__24762\
        );

    \I__3477\ : LocalMux
    port map (
            O => \N__24765\,
            I => \ADC_IAC.bit_cnt_2\
        );

    \I__3476\ : LocalMux
    port map (
            O => \N__24762\,
            I => \ADC_IAC.bit_cnt_2\
        );

    \I__3475\ : InMux
    port map (
            O => \N__24757\,
            I => \N__24753\
        );

    \I__3474\ : InMux
    port map (
            O => \N__24756\,
            I => \N__24750\
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__24753\,
            I => \ADC_IAC.bit_cnt_6\
        );

    \I__3472\ : LocalMux
    port map (
            O => \N__24750\,
            I => \ADC_IAC.bit_cnt_6\
        );

    \I__3471\ : InMux
    port map (
            O => \N__24745\,
            I => \N__24741\
        );

    \I__3470\ : InMux
    port map (
            O => \N__24744\,
            I => \N__24738\
        );

    \I__3469\ : LocalMux
    port map (
            O => \N__24741\,
            I => \ADC_IAC.bit_cnt_0\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__24738\,
            I => \ADC_IAC.bit_cnt_0\
        );

    \I__3467\ : CascadeMux
    port map (
            O => \N__24733\,
            I => \ADC_IAC.n20753_cascade_\
        );

    \I__3466\ : InMux
    port map (
            O => \N__24730\,
            I => \N__24726\
        );

    \I__3465\ : InMux
    port map (
            O => \N__24729\,
            I => \N__24723\
        );

    \I__3464\ : LocalMux
    port map (
            O => \N__24726\,
            I => \ADC_IAC.bit_cnt_7\
        );

    \I__3463\ : LocalMux
    port map (
            O => \N__24723\,
            I => \ADC_IAC.bit_cnt_7\
        );

    \I__3462\ : CascadeMux
    port map (
            O => \N__24718\,
            I => \N__24715\
        );

    \I__3461\ : InMux
    port map (
            O => \N__24715\,
            I => \N__24712\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__24712\,
            I => \N__24708\
        );

    \I__3459\ : InMux
    port map (
            O => \N__24711\,
            I => \N__24705\
        );

    \I__3458\ : Odrv4
    port map (
            O => \N__24708\,
            I => cmd_rdadctmp_5
        );

    \I__3457\ : LocalMux
    port map (
            O => \N__24705\,
            I => cmd_rdadctmp_5
        );

    \I__3456\ : InMux
    port map (
            O => \N__24700\,
            I => \N__24697\
        );

    \I__3455\ : LocalMux
    port map (
            O => \N__24697\,
            I => \N__24694\
        );

    \I__3454\ : Span4Mux_v
    port map (
            O => \N__24694\,
            I => \N__24691\
        );

    \I__3453\ : Span4Mux_v
    port map (
            O => \N__24691\,
            I => \N__24687\
        );

    \I__3452\ : InMux
    port map (
            O => \N__24690\,
            I => \N__24684\
        );

    \I__3451\ : Span4Mux_v
    port map (
            O => \N__24687\,
            I => \N__24678\
        );

    \I__3450\ : LocalMux
    port map (
            O => \N__24684\,
            I => \N__24678\
        );

    \I__3449\ : InMux
    port map (
            O => \N__24683\,
            I => \N__24675\
        );

    \I__3448\ : Span4Mux_h
    port map (
            O => \N__24678\,
            I => \N__24672\
        );

    \I__3447\ : LocalMux
    port map (
            O => \N__24675\,
            I => buf_adcdata_iac_22
        );

    \I__3446\ : Odrv4
    port map (
            O => \N__24672\,
            I => buf_adcdata_iac_22
        );

    \I__3445\ : InMux
    port map (
            O => \N__24667\,
            I => \N__24661\
        );

    \I__3444\ : InMux
    port map (
            O => \N__24666\,
            I => \N__24661\
        );

    \I__3443\ : LocalMux
    port map (
            O => \N__24661\,
            I => cmd_rdadctmp_1
        );

    \I__3442\ : InMux
    port map (
            O => \N__24658\,
            I => \N__24654\
        );

    \I__3441\ : InMux
    port map (
            O => \N__24657\,
            I => \N__24651\
        );

    \I__3440\ : LocalMux
    port map (
            O => \N__24654\,
            I => n20553
        );

    \I__3439\ : LocalMux
    port map (
            O => \N__24651\,
            I => n20553
        );

    \I__3438\ : CascadeMux
    port map (
            O => \N__24646\,
            I => \N__24641\
        );

    \I__3437\ : CascadeMux
    port map (
            O => \N__24645\,
            I => \N__24638\
        );

    \I__3436\ : CascadeMux
    port map (
            O => \N__24644\,
            I => \N__24635\
        );

    \I__3435\ : InMux
    port map (
            O => \N__24641\,
            I => \N__24632\
        );

    \I__3434\ : InMux
    port map (
            O => \N__24638\,
            I => \N__24629\
        );

    \I__3433\ : InMux
    port map (
            O => \N__24635\,
            I => \N__24626\
        );

    \I__3432\ : LocalMux
    port map (
            O => \N__24632\,
            I => \N__24623\
        );

    \I__3431\ : LocalMux
    port map (
            O => \N__24629\,
            I => cmd_rdadctmp_29
        );

    \I__3430\ : LocalMux
    port map (
            O => \N__24626\,
            I => cmd_rdadctmp_29
        );

    \I__3429\ : Odrv4
    port map (
            O => \N__24623\,
            I => cmd_rdadctmp_29
        );

    \I__3428\ : CascadeMux
    port map (
            O => \N__24616\,
            I => \N__24613\
        );

    \I__3427\ : InMux
    port map (
            O => \N__24613\,
            I => \N__24608\
        );

    \I__3426\ : InMux
    port map (
            O => \N__24612\,
            I => \N__24605\
        );

    \I__3425\ : InMux
    port map (
            O => \N__24611\,
            I => \N__24602\
        );

    \I__3424\ : LocalMux
    port map (
            O => \N__24608\,
            I => cmd_rdadctmp_27
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__24605\,
            I => cmd_rdadctmp_27
        );

    \I__3422\ : LocalMux
    port map (
            O => \N__24602\,
            I => cmd_rdadctmp_27
        );

    \I__3421\ : CascadeMux
    port map (
            O => \N__24595\,
            I => \N__24592\
        );

    \I__3420\ : InMux
    port map (
            O => \N__24592\,
            I => \N__24589\
        );

    \I__3419\ : LocalMux
    port map (
            O => \N__24589\,
            I => \N__24586\
        );

    \I__3418\ : Span4Mux_v
    port map (
            O => \N__24586\,
            I => \N__24583\
        );

    \I__3417\ : Sp12to4
    port map (
            O => \N__24583\,
            I => \N__24580\
        );

    \I__3416\ : Span12Mux_h
    port map (
            O => \N__24580\,
            I => \N__24577\
        );

    \I__3415\ : Odrv12
    port map (
            O => \N__24577\,
            I => \IAC_MISO\
        );

    \I__3414\ : InMux
    port map (
            O => \N__24574\,
            I => \N__24570\
        );

    \I__3413\ : InMux
    port map (
            O => \N__24573\,
            I => \N__24567\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__24570\,
            I => cmd_rdadctmp_0
        );

    \I__3411\ : LocalMux
    port map (
            O => \N__24567\,
            I => cmd_rdadctmp_0
        );

    \I__3410\ : CascadeMux
    port map (
            O => \N__24562\,
            I => \N__24559\
        );

    \I__3409\ : InMux
    port map (
            O => \N__24559\,
            I => \N__24553\
        );

    \I__3408\ : InMux
    port map (
            O => \N__24558\,
            I => \N__24553\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__24553\,
            I => cmd_rdadctmp_6
        );

    \I__3406\ : CascadeMux
    port map (
            O => \N__24550\,
            I => \N__24547\
        );

    \I__3405\ : CascadeBuf
    port map (
            O => \N__24547\,
            I => \N__24544\
        );

    \I__3404\ : CascadeMux
    port map (
            O => \N__24544\,
            I => \N__24541\
        );

    \I__3403\ : CascadeBuf
    port map (
            O => \N__24541\,
            I => \N__24538\
        );

    \I__3402\ : CascadeMux
    port map (
            O => \N__24538\,
            I => \N__24535\
        );

    \I__3401\ : CascadeBuf
    port map (
            O => \N__24535\,
            I => \N__24532\
        );

    \I__3400\ : CascadeMux
    port map (
            O => \N__24532\,
            I => \N__24529\
        );

    \I__3399\ : CascadeBuf
    port map (
            O => \N__24529\,
            I => \N__24526\
        );

    \I__3398\ : CascadeMux
    port map (
            O => \N__24526\,
            I => \N__24523\
        );

    \I__3397\ : CascadeBuf
    port map (
            O => \N__24523\,
            I => \N__24520\
        );

    \I__3396\ : CascadeMux
    port map (
            O => \N__24520\,
            I => \N__24517\
        );

    \I__3395\ : CascadeBuf
    port map (
            O => \N__24517\,
            I => \N__24514\
        );

    \I__3394\ : CascadeMux
    port map (
            O => \N__24514\,
            I => \N__24510\
        );

    \I__3393\ : CascadeMux
    port map (
            O => \N__24513\,
            I => \N__24507\
        );

    \I__3392\ : CascadeBuf
    port map (
            O => \N__24510\,
            I => \N__24504\
        );

    \I__3391\ : CascadeBuf
    port map (
            O => \N__24507\,
            I => \N__24501\
        );

    \I__3390\ : CascadeMux
    port map (
            O => \N__24504\,
            I => \N__24498\
        );

    \I__3389\ : CascadeMux
    port map (
            O => \N__24501\,
            I => \N__24495\
        );

    \I__3388\ : CascadeBuf
    port map (
            O => \N__24498\,
            I => \N__24492\
        );

    \I__3387\ : InMux
    port map (
            O => \N__24495\,
            I => \N__24489\
        );

    \I__3386\ : CascadeMux
    port map (
            O => \N__24492\,
            I => \N__24486\
        );

    \I__3385\ : LocalMux
    port map (
            O => \N__24489\,
            I => \N__24483\
        );

    \I__3384\ : CascadeBuf
    port map (
            O => \N__24486\,
            I => \N__24480\
        );

    \I__3383\ : Span4Mux_v
    port map (
            O => \N__24483\,
            I => \N__24477\
        );

    \I__3382\ : CascadeMux
    port map (
            O => \N__24480\,
            I => \N__24474\
        );

    \I__3381\ : Span4Mux_h
    port map (
            O => \N__24477\,
            I => \N__24471\
        );

    \I__3380\ : InMux
    port map (
            O => \N__24474\,
            I => \N__24468\
        );

    \I__3379\ : Span4Mux_h
    port map (
            O => \N__24471\,
            I => \N__24465\
        );

    \I__3378\ : LocalMux
    port map (
            O => \N__24468\,
            I => \N__24462\
        );

    \I__3377\ : Span4Mux_h
    port map (
            O => \N__24465\,
            I => \N__24457\
        );

    \I__3376\ : Span4Mux_v
    port map (
            O => \N__24462\,
            I => \N__24457\
        );

    \I__3375\ : Odrv4
    port map (
            O => \N__24457\,
            I => \data_index_9_N_212_8\
        );

    \I__3374\ : InMux
    port map (
            O => \N__24454\,
            I => \N__24450\
        );

    \I__3373\ : CascadeMux
    port map (
            O => \N__24453\,
            I => \N__24447\
        );

    \I__3372\ : LocalMux
    port map (
            O => \N__24450\,
            I => \N__24443\
        );

    \I__3371\ : InMux
    port map (
            O => \N__24447\,
            I => \N__24438\
        );

    \I__3370\ : InMux
    port map (
            O => \N__24446\,
            I => \N__24438\
        );

    \I__3369\ : Odrv4
    port map (
            O => \N__24443\,
            I => cmd_rdadctmp_22
        );

    \I__3368\ : LocalMux
    port map (
            O => \N__24438\,
            I => cmd_rdadctmp_22
        );

    \I__3367\ : InMux
    port map (
            O => \N__24433\,
            I => \N__24427\
        );

    \I__3366\ : InMux
    port map (
            O => \N__24432\,
            I => \N__24427\
        );

    \I__3365\ : LocalMux
    port map (
            O => \N__24427\,
            I => n8_adj_1534
        );

    \I__3364\ : InMux
    port map (
            O => \N__24424\,
            I => \N__24421\
        );

    \I__3363\ : LocalMux
    port map (
            O => \N__24421\,
            I => \N__24417\
        );

    \I__3362\ : CascadeMux
    port map (
            O => \N__24420\,
            I => \N__24414\
        );

    \I__3361\ : Span4Mux_v
    port map (
            O => \N__24417\,
            I => \N__24410\
        );

    \I__3360\ : InMux
    port map (
            O => \N__24414\,
            I => \N__24407\
        );

    \I__3359\ : InMux
    port map (
            O => \N__24413\,
            I => \N__24404\
        );

    \I__3358\ : Span4Mux_h
    port map (
            O => \N__24410\,
            I => \N__24399\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__24407\,
            I => \N__24399\
        );

    \I__3356\ : LocalMux
    port map (
            O => \N__24404\,
            I => buf_adcdata_iac_8
        );

    \I__3355\ : Odrv4
    port map (
            O => \N__24399\,
            I => buf_adcdata_iac_8
        );

    \I__3354\ : InMux
    port map (
            O => \N__24394\,
            I => \N__24391\
        );

    \I__3353\ : LocalMux
    port map (
            O => \N__24391\,
            I => \N__24388\
        );

    \I__3352\ : Span4Mux_v
    port map (
            O => \N__24388\,
            I => \N__24385\
        );

    \I__3351\ : Span4Mux_h
    port map (
            O => \N__24385\,
            I => \N__24382\
        );

    \I__3350\ : Sp12to4
    port map (
            O => \N__24382\,
            I => \N__24379\
        );

    \I__3349\ : Odrv12
    port map (
            O => \N__24379\,
            I => buf_data_iac_23
        );

    \I__3348\ : CascadeMux
    port map (
            O => \N__24376\,
            I => \n26_adj_1511_cascade_\
        );

    \I__3347\ : CascadeMux
    port map (
            O => \N__24373\,
            I => \n20834_cascade_\
        );

    \I__3346\ : CascadeMux
    port map (
            O => \N__24370\,
            I => \n22057_cascade_\
        );

    \I__3345\ : InMux
    port map (
            O => \N__24367\,
            I => \N__24364\
        );

    \I__3344\ : LocalMux
    port map (
            O => \N__24364\,
            I => \N__24361\
        );

    \I__3343\ : Span4Mux_v
    port map (
            O => \N__24361\,
            I => \N__24358\
        );

    \I__3342\ : Odrv4
    port map (
            O => \N__24358\,
            I => buf_data_iac_12
        );

    \I__3341\ : InMux
    port map (
            O => \N__24355\,
            I => \N__24352\
        );

    \I__3340\ : LocalMux
    port map (
            O => \N__24352\,
            I => \N__24349\
        );

    \I__3339\ : Odrv4
    port map (
            O => \N__24349\,
            I => n22135
        );

    \I__3338\ : InMux
    port map (
            O => \N__24346\,
            I => \N__24343\
        );

    \I__3337\ : LocalMux
    port map (
            O => \N__24343\,
            I => \N__24339\
        );

    \I__3336\ : InMux
    port map (
            O => \N__24342\,
            I => \N__24335\
        );

    \I__3335\ : Span4Mux_v
    port map (
            O => \N__24339\,
            I => \N__24332\
        );

    \I__3334\ : CascadeMux
    port map (
            O => \N__24338\,
            I => \N__24329\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__24335\,
            I => \N__24326\
        );

    \I__3332\ : Span4Mux_v
    port map (
            O => \N__24332\,
            I => \N__24323\
        );

    \I__3331\ : InMux
    port map (
            O => \N__24329\,
            I => \N__24320\
        );

    \I__3330\ : Span4Mux_v
    port map (
            O => \N__24326\,
            I => \N__24315\
        );

    \I__3329\ : Span4Mux_v
    port map (
            O => \N__24323\,
            I => \N__24315\
        );

    \I__3328\ : LocalMux
    port map (
            O => \N__24320\,
            I => buf_adcdata_vac_23
        );

    \I__3327\ : Odrv4
    port map (
            O => \N__24315\,
            I => buf_adcdata_vac_23
        );

    \I__3326\ : InMux
    port map (
            O => \N__24310\,
            I => \N__24306\
        );

    \I__3325\ : CascadeMux
    port map (
            O => \N__24309\,
            I => \N__24303\
        );

    \I__3324\ : LocalMux
    port map (
            O => \N__24306\,
            I => \N__24300\
        );

    \I__3323\ : InMux
    port map (
            O => \N__24303\,
            I => \N__24297\
        );

    \I__3322\ : Odrv12
    port map (
            O => \N__24300\,
            I => buf_adcdata_vdc_23
        );

    \I__3321\ : LocalMux
    port map (
            O => \N__24297\,
            I => buf_adcdata_vdc_23
        );

    \I__3320\ : InMux
    port map (
            O => \N__24292\,
            I => \N__24289\
        );

    \I__3319\ : LocalMux
    port map (
            O => \N__24289\,
            I => n20831
        );

    \I__3318\ : InMux
    port map (
            O => \N__24286\,
            I => \N__24283\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__24283\,
            I => \N__24280\
        );

    \I__3316\ : Span4Mux_h
    port map (
            O => \N__24280\,
            I => \N__24276\
        );

    \I__3315\ : InMux
    port map (
            O => \N__24279\,
            I => \N__24273\
        );

    \I__3314\ : Odrv4
    port map (
            O => \N__24276\,
            I => cmd_rdadctmp_7
        );

    \I__3313\ : LocalMux
    port map (
            O => \N__24273\,
            I => cmd_rdadctmp_7
        );

    \I__3312\ : InMux
    port map (
            O => \N__24268\,
            I => \N__24265\
        );

    \I__3311\ : LocalMux
    port map (
            O => \N__24265\,
            I => \N__24262\
        );

    \I__3310\ : Span4Mux_v
    port map (
            O => \N__24262\,
            I => \N__24259\
        );

    \I__3309\ : Odrv4
    port map (
            O => \N__24259\,
            I => n16_adj_1507
        );

    \I__3308\ : InMux
    port map (
            O => \N__24256\,
            I => \N__24252\
        );

    \I__3307\ : InMux
    port map (
            O => \N__24255\,
            I => \N__24248\
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__24252\,
            I => \N__24245\
        );

    \I__3305\ : InMux
    port map (
            O => \N__24251\,
            I => \N__24242\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__24248\,
            I => cmd_rdadctmp_24_adj_1419
        );

    \I__3303\ : Odrv4
    port map (
            O => \N__24245\,
            I => cmd_rdadctmp_24_adj_1419
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__24242\,
            I => cmd_rdadctmp_24_adj_1419
        );

    \I__3301\ : InMux
    port map (
            O => \N__24235\,
            I => \N__24231\
        );

    \I__3300\ : InMux
    port map (
            O => \N__24234\,
            I => \N__24227\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__24231\,
            I => \N__24224\
        );

    \I__3298\ : InMux
    port map (
            O => \N__24230\,
            I => \N__24221\
        );

    \I__3297\ : LocalMux
    port map (
            O => \N__24227\,
            I => cmd_rdadctmp_25_adj_1418
        );

    \I__3296\ : Odrv4
    port map (
            O => \N__24224\,
            I => cmd_rdadctmp_25_adj_1418
        );

    \I__3295\ : LocalMux
    port map (
            O => \N__24221\,
            I => cmd_rdadctmp_25_adj_1418
        );

    \I__3294\ : InMux
    port map (
            O => \N__24214\,
            I => \N__24211\
        );

    \I__3293\ : LocalMux
    port map (
            O => \N__24211\,
            I => \N__24208\
        );

    \I__3292\ : Odrv4
    port map (
            O => \N__24208\,
            I => n22039
        );

    \I__3291\ : InMux
    port map (
            O => \N__24205\,
            I => \N__24202\
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__24202\,
            I => n22042
        );

    \I__3289\ : CascadeMux
    port map (
            O => \N__24199\,
            I => \N__24196\
        );

    \I__3288\ : InMux
    port map (
            O => \N__24196\,
            I => \N__24191\
        );

    \I__3287\ : CascadeMux
    port map (
            O => \N__24195\,
            I => \N__24188\
        );

    \I__3286\ : CascadeMux
    port map (
            O => \N__24194\,
            I => \N__24185\
        );

    \I__3285\ : LocalMux
    port map (
            O => \N__24191\,
            I => \N__24182\
        );

    \I__3284\ : InMux
    port map (
            O => \N__24188\,
            I => \N__24179\
        );

    \I__3283\ : InMux
    port map (
            O => \N__24185\,
            I => \N__24176\
        );

    \I__3282\ : Span4Mux_v
    port map (
            O => \N__24182\,
            I => \N__24172\
        );

    \I__3281\ : LocalMux
    port map (
            O => \N__24179\,
            I => \N__24167\
        );

    \I__3280\ : LocalMux
    port map (
            O => \N__24176\,
            I => \N__24167\
        );

    \I__3279\ : InMux
    port map (
            O => \N__24175\,
            I => \N__24163\
        );

    \I__3278\ : Span4Mux_v
    port map (
            O => \N__24172\,
            I => \N__24160\
        );

    \I__3277\ : Span4Mux_h
    port map (
            O => \N__24167\,
            I => \N__24157\
        );

    \I__3276\ : InMux
    port map (
            O => \N__24166\,
            I => \N__24154\
        );

    \I__3275\ : LocalMux
    port map (
            O => \N__24163\,
            I => \N__24151\
        );

    \I__3274\ : Odrv4
    port map (
            O => \N__24160\,
            I => \buf_cfgRTD_7\
        );

    \I__3273\ : Odrv4
    port map (
            O => \N__24157\,
            I => \buf_cfgRTD_7\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__24154\,
            I => \buf_cfgRTD_7\
        );

    \I__3271\ : Odrv4
    port map (
            O => \N__24151\,
            I => \buf_cfgRTD_7\
        );

    \I__3270\ : CascadeMux
    port map (
            O => \N__24142\,
            I => \N__24139\
        );

    \I__3269\ : InMux
    port map (
            O => \N__24139\,
            I => \N__24135\
        );

    \I__3268\ : CascadeMux
    port map (
            O => \N__24138\,
            I => \N__24132\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__24135\,
            I => \N__24129\
        );

    \I__3266\ : InMux
    port map (
            O => \N__24132\,
            I => \N__24125\
        );

    \I__3265\ : Span4Mux_h
    port map (
            O => \N__24129\,
            I => \N__24122\
        );

    \I__3264\ : InMux
    port map (
            O => \N__24128\,
            I => \N__24119\
        );

    \I__3263\ : LocalMux
    port map (
            O => \N__24125\,
            I => cmd_rdadctmp_20_adj_1423
        );

    \I__3262\ : Odrv4
    port map (
            O => \N__24122\,
            I => cmd_rdadctmp_20_adj_1423
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__24119\,
            I => cmd_rdadctmp_20_adj_1423
        );

    \I__3260\ : InMux
    port map (
            O => \N__24112\,
            I => \N__24107\
        );

    \I__3259\ : InMux
    port map (
            O => \N__24111\,
            I => \N__24102\
        );

    \I__3258\ : InMux
    port map (
            O => \N__24110\,
            I => \N__24102\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__24107\,
            I => cmd_rdadctmp_18_adj_1425
        );

    \I__3256\ : LocalMux
    port map (
            O => \N__24102\,
            I => cmd_rdadctmp_18_adj_1425
        );

    \I__3255\ : InMux
    port map (
            O => \N__24097\,
            I => \N__24094\
        );

    \I__3254\ : LocalMux
    port map (
            O => \N__24094\,
            I => \N__24091\
        );

    \I__3253\ : Span4Mux_h
    port map (
            O => \N__24091\,
            I => \N__24086\
        );

    \I__3252\ : InMux
    port map (
            O => \N__24090\,
            I => \N__24081\
        );

    \I__3251\ : InMux
    port map (
            O => \N__24089\,
            I => \N__24081\
        );

    \I__3250\ : Odrv4
    port map (
            O => \N__24086\,
            I => buf_adcdata_vac_12
        );

    \I__3249\ : LocalMux
    port map (
            O => \N__24081\,
            I => buf_adcdata_vac_12
        );

    \I__3248\ : InMux
    port map (
            O => \N__24076\,
            I => \N__24073\
        );

    \I__3247\ : LocalMux
    port map (
            O => \N__24073\,
            I => \N__24069\
        );

    \I__3246\ : CascadeMux
    port map (
            O => \N__24072\,
            I => \N__24066\
        );

    \I__3245\ : Span4Mux_v
    port map (
            O => \N__24069\,
            I => \N__24063\
        );

    \I__3244\ : InMux
    port map (
            O => \N__24066\,
            I => \N__24060\
        );

    \I__3243\ : Odrv4
    port map (
            O => \N__24063\,
            I => buf_adcdata_vdc_10
        );

    \I__3242\ : LocalMux
    port map (
            O => \N__24060\,
            I => buf_adcdata_vdc_10
        );

    \I__3241\ : InMux
    port map (
            O => \N__24055\,
            I => \N__24052\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__24052\,
            I => \N__24049\
        );

    \I__3239\ : Span4Mux_v
    port map (
            O => \N__24049\,
            I => \N__24046\
        );

    \I__3238\ : Span4Mux_h
    port map (
            O => \N__24046\,
            I => \N__24041\
        );

    \I__3237\ : InMux
    port map (
            O => \N__24045\,
            I => \N__24036\
        );

    \I__3236\ : InMux
    port map (
            O => \N__24044\,
            I => \N__24036\
        );

    \I__3235\ : Odrv4
    port map (
            O => \N__24041\,
            I => buf_adcdata_vac_10
        );

    \I__3234\ : LocalMux
    port map (
            O => \N__24036\,
            I => buf_adcdata_vac_10
        );

    \I__3233\ : CascadeMux
    port map (
            O => \N__24031\,
            I => \N__24027\
        );

    \I__3232\ : CascadeMux
    port map (
            O => \N__24030\,
            I => \N__24024\
        );

    \I__3231\ : InMux
    port map (
            O => \N__24027\,
            I => \N__24021\
        );

    \I__3230\ : InMux
    port map (
            O => \N__24024\,
            I => \N__24017\
        );

    \I__3229\ : LocalMux
    port map (
            O => \N__24021\,
            I => \N__24014\
        );

    \I__3228\ : InMux
    port map (
            O => \N__24020\,
            I => \N__24011\
        );

    \I__3227\ : LocalMux
    port map (
            O => \N__24017\,
            I => cmd_rdadctmp_19_adj_1424
        );

    \I__3226\ : Odrv4
    port map (
            O => \N__24014\,
            I => cmd_rdadctmp_19_adj_1424
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__24011\,
            I => cmd_rdadctmp_19_adj_1424
        );

    \I__3224\ : CascadeMux
    port map (
            O => \N__24004\,
            I => \N__24001\
        );

    \I__3223\ : InMux
    port map (
            O => \N__24001\,
            I => \N__23998\
        );

    \I__3222\ : LocalMux
    port map (
            O => \N__23998\,
            I => \N__23995\
        );

    \I__3221\ : Span4Mux_h
    port map (
            O => \N__23995\,
            I => \N__23992\
        );

    \I__3220\ : Odrv4
    port map (
            O => \N__23992\,
            I => buf_data_iac_16
        );

    \I__3219\ : CascadeMux
    port map (
            O => \N__23989\,
            I => \n20781_cascade_\
        );

    \I__3218\ : InMux
    port map (
            O => \N__23986\,
            I => \N__23982\
        );

    \I__3217\ : CascadeMux
    port map (
            O => \N__23985\,
            I => \N__23979\
        );

    \I__3216\ : LocalMux
    port map (
            O => \N__23982\,
            I => \N__23976\
        );

    \I__3215\ : InMux
    port map (
            O => \N__23979\,
            I => \N__23973\
        );

    \I__3214\ : Odrv12
    port map (
            O => \N__23976\,
            I => buf_adcdata_vdc_1
        );

    \I__3213\ : LocalMux
    port map (
            O => \N__23973\,
            I => buf_adcdata_vdc_1
        );

    \I__3212\ : InMux
    port map (
            O => \N__23968\,
            I => \N__23965\
        );

    \I__3211\ : LocalMux
    port map (
            O => \N__23965\,
            I => \N__23962\
        );

    \I__3210\ : Span4Mux_v
    port map (
            O => \N__23962\,
            I => \N__23957\
        );

    \I__3209\ : InMux
    port map (
            O => \N__23961\,
            I => \N__23954\
        );

    \I__3208\ : InMux
    port map (
            O => \N__23960\,
            I => \N__23951\
        );

    \I__3207\ : Span4Mux_h
    port map (
            O => \N__23957\,
            I => \N__23946\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__23954\,
            I => \N__23946\
        );

    \I__3205\ : LocalMux
    port map (
            O => \N__23951\,
            I => buf_adcdata_vac_1
        );

    \I__3204\ : Odrv4
    port map (
            O => \N__23946\,
            I => buf_adcdata_vac_1
        );

    \I__3203\ : InMux
    port map (
            O => \N__23941\,
            I => \N__23938\
        );

    \I__3202\ : LocalMux
    port map (
            O => \N__23938\,
            I => n19_adj_1617
        );

    \I__3201\ : CascadeMux
    port map (
            O => \N__23935\,
            I => \n22171_cascade_\
        );

    \I__3200\ : InMux
    port map (
            O => \N__23932\,
            I => \N__23929\
        );

    \I__3199\ : LocalMux
    port map (
            O => \N__23929\,
            I => \N__23926\
        );

    \I__3198\ : Odrv4
    port map (
            O => \N__23926\,
            I => n20775
        );

    \I__3197\ : InMux
    port map (
            O => \N__23923\,
            I => \N__23920\
        );

    \I__3196\ : LocalMux
    port map (
            O => \N__23920\,
            I => \N__23917\
        );

    \I__3195\ : Span4Mux_h
    port map (
            O => \N__23917\,
            I => \N__23914\
        );

    \I__3194\ : Odrv4
    port map (
            O => \N__23914\,
            I => n20842
        );

    \I__3193\ : CascadeMux
    port map (
            O => \N__23911\,
            I => \N__23908\
        );

    \I__3192\ : InMux
    port map (
            O => \N__23908\,
            I => \N__23905\
        );

    \I__3191\ : LocalMux
    port map (
            O => \N__23905\,
            I => \N__23902\
        );

    \I__3190\ : Odrv4
    port map (
            O => \N__23902\,
            I => n20843
        );

    \I__3189\ : CascadeMux
    port map (
            O => \N__23899\,
            I => \n22051_cascade_\
        );

    \I__3188\ : InMux
    port map (
            O => \N__23896\,
            I => \N__23893\
        );

    \I__3187\ : LocalMux
    port map (
            O => \N__23893\,
            I => \N__23890\
        );

    \I__3186\ : Odrv4
    port map (
            O => \N__23890\,
            I => n20828
        );

    \I__3185\ : InMux
    port map (
            O => \N__23887\,
            I => \N__23884\
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__23884\,
            I => \N__23881\
        );

    \I__3183\ : Odrv4
    port map (
            O => \N__23881\,
            I => n20814
        );

    \I__3182\ : InMux
    port map (
            O => \N__23878\,
            I => \N__23875\
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__23875\,
            I => \N__23871\
        );

    \I__3180\ : CascadeMux
    port map (
            O => \N__23874\,
            I => \N__23868\
        );

    \I__3179\ : Span4Mux_v
    port map (
            O => \N__23871\,
            I => \N__23865\
        );

    \I__3178\ : InMux
    port map (
            O => \N__23868\,
            I => \N__23862\
        );

    \I__3177\ : Odrv4
    port map (
            O => \N__23865\,
            I => buf_adcdata_vdc_18
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__23862\,
            I => buf_adcdata_vdc_18
        );

    \I__3175\ : InMux
    port map (
            O => \N__23857\,
            I => \N__23853\
        );

    \I__3174\ : InMux
    port map (
            O => \N__23856\,
            I => \N__23849\
        );

    \I__3173\ : LocalMux
    port map (
            O => \N__23853\,
            I => \N__23846\
        );

    \I__3172\ : InMux
    port map (
            O => \N__23852\,
            I => \N__23843\
        );

    \I__3171\ : LocalMux
    port map (
            O => \N__23849\,
            I => \N__23840\
        );

    \I__3170\ : Span4Mux_v
    port map (
            O => \N__23846\,
            I => \N__23837\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__23843\,
            I => buf_adcdata_vac_18
        );

    \I__3168\ : Odrv4
    port map (
            O => \N__23840\,
            I => buf_adcdata_vac_18
        );

    \I__3167\ : Odrv4
    port map (
            O => \N__23837\,
            I => buf_adcdata_vac_18
        );

    \I__3166\ : CascadeMux
    port map (
            O => \N__23830\,
            I => \n21931_cascade_\
        );

    \I__3165\ : InMux
    port map (
            O => \N__23827\,
            I => \N__23824\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__23824\,
            I => \N__23820\
        );

    \I__3163\ : CascadeMux
    port map (
            O => \N__23823\,
            I => \N__23816\
        );

    \I__3162\ : Span4Mux_v
    port map (
            O => \N__23820\,
            I => \N__23813\
        );

    \I__3161\ : InMux
    port map (
            O => \N__23819\,
            I => \N__23810\
        );

    \I__3160\ : InMux
    port map (
            O => \N__23816\,
            I => \N__23807\
        );

    \I__3159\ : Sp12to4
    port map (
            O => \N__23813\,
            I => \N__23800\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__23810\,
            I => \N__23800\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__23807\,
            I => \N__23797\
        );

    \I__3156\ : InMux
    port map (
            O => \N__23806\,
            I => \N__23792\
        );

    \I__3155\ : InMux
    port map (
            O => \N__23805\,
            I => \N__23792\
        );

    \I__3154\ : Odrv12
    port map (
            O => \N__23800\,
            I => \buf_cfgRTD_2\
        );

    \I__3153\ : Odrv4
    port map (
            O => \N__23797\,
            I => \buf_cfgRTD_2\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__23792\,
            I => \buf_cfgRTD_2\
        );

    \I__3151\ : CascadeMux
    port map (
            O => \N__23785\,
            I => \N__23782\
        );

    \I__3150\ : InMux
    port map (
            O => \N__23782\,
            I => \N__23779\
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__23779\,
            I => \N__23774\
        );

    \I__3148\ : CascadeMux
    port map (
            O => \N__23778\,
            I => \N__23771\
        );

    \I__3147\ : CascadeMux
    port map (
            O => \N__23777\,
            I => \N__23768\
        );

    \I__3146\ : Span4Mux_h
    port map (
            O => \N__23774\,
            I => \N__23764\
        );

    \I__3145\ : InMux
    port map (
            O => \N__23771\,
            I => \N__23760\
        );

    \I__3144\ : InMux
    port map (
            O => \N__23768\,
            I => \N__23755\
        );

    \I__3143\ : InMux
    port map (
            O => \N__23767\,
            I => \N__23755\
        );

    \I__3142\ : Sp12to4
    port map (
            O => \N__23764\,
            I => \N__23752\
        );

    \I__3141\ : InMux
    port map (
            O => \N__23763\,
            I => \N__23749\
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__23760\,
            I => \N__23744\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__23755\,
            I => \N__23744\
        );

    \I__3138\ : Odrv12
    port map (
            O => \N__23752\,
            I => \buf_cfgRTD_3\
        );

    \I__3137\ : LocalMux
    port map (
            O => \N__23749\,
            I => \buf_cfgRTD_3\
        );

    \I__3136\ : Odrv4
    port map (
            O => \N__23744\,
            I => \buf_cfgRTD_3\
        );

    \I__3135\ : CascadeMux
    port map (
            O => \N__23737\,
            I => \N__23734\
        );

    \I__3134\ : InMux
    port map (
            O => \N__23734\,
            I => \N__23729\
        );

    \I__3133\ : InMux
    port map (
            O => \N__23733\,
            I => \N__23724\
        );

    \I__3132\ : InMux
    port map (
            O => \N__23732\,
            I => \N__23724\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__23729\,
            I => \N__23719\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__23724\,
            I => \N__23719\
        );

    \I__3129\ : Span4Mux_v
    port map (
            O => \N__23719\,
            I => \N__23714\
        );

    \I__3128\ : InMux
    port map (
            O => \N__23718\,
            I => \N__23711\
        );

    \I__3127\ : InMux
    port map (
            O => \N__23717\,
            I => \N__23708\
        );

    \I__3126\ : Odrv4
    port map (
            O => \N__23714\,
            I => \buf_cfgRTD_0\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__23711\,
            I => \buf_cfgRTD_0\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__23708\,
            I => \buf_cfgRTD_0\
        );

    \I__3123\ : CascadeMux
    port map (
            O => \N__23701\,
            I => \n14490_cascade_\
        );

    \I__3122\ : CascadeMux
    port map (
            O => \N__23698\,
            I => \N__23694\
        );

    \I__3121\ : InMux
    port map (
            O => \N__23697\,
            I => \N__23691\
        );

    \I__3120\ : InMux
    port map (
            O => \N__23694\,
            I => \N__23688\
        );

    \I__3119\ : LocalMux
    port map (
            O => \N__23691\,
            I => \N__23683\
        );

    \I__3118\ : LocalMux
    port map (
            O => \N__23688\,
            I => \N__23683\
        );

    \I__3117\ : Span4Mux_v
    port map (
            O => \N__23683\,
            I => \N__23677\
        );

    \I__3116\ : InMux
    port map (
            O => \N__23682\,
            I => \N__23674\
        );

    \I__3115\ : InMux
    port map (
            O => \N__23681\,
            I => \N__23671\
        );

    \I__3114\ : InMux
    port map (
            O => \N__23680\,
            I => \N__23668\
        );

    \I__3113\ : Odrv4
    port map (
            O => \N__23677\,
            I => \buf_cfgRTD_1\
        );

    \I__3112\ : LocalMux
    port map (
            O => \N__23674\,
            I => \buf_cfgRTD_1\
        );

    \I__3111\ : LocalMux
    port map (
            O => \N__23671\,
            I => \buf_cfgRTD_1\
        );

    \I__3110\ : LocalMux
    port map (
            O => \N__23668\,
            I => \buf_cfgRTD_1\
        );

    \I__3109\ : CascadeMux
    port map (
            O => \N__23659\,
            I => \N__23656\
        );

    \I__3108\ : InMux
    port map (
            O => \N__23656\,
            I => \N__23653\
        );

    \I__3107\ : LocalMux
    port map (
            O => \N__23653\,
            I => \N__23650\
        );

    \I__3106\ : Span4Mux_v
    port map (
            O => \N__23650\,
            I => \N__23647\
        );

    \I__3105\ : Span4Mux_h
    port map (
            O => \N__23647\,
            I => \N__23643\
        );

    \I__3104\ : InMux
    port map (
            O => \N__23646\,
            I => \N__23640\
        );

    \I__3103\ : Odrv4
    port map (
            O => \N__23643\,
            I => \buf_readRTD_9\
        );

    \I__3102\ : LocalMux
    port map (
            O => \N__23640\,
            I => \buf_readRTD_9\
        );

    \I__3101\ : InMux
    port map (
            O => \N__23635\,
            I => \N__23632\
        );

    \I__3100\ : LocalMux
    port map (
            O => \N__23632\,
            I => n22165
        );

    \I__3099\ : InMux
    port map (
            O => \N__23629\,
            I => \N__23624\
        );

    \I__3098\ : InMux
    port map (
            O => \N__23628\,
            I => \N__23621\
        );

    \I__3097\ : CascadeMux
    port map (
            O => \N__23627\,
            I => \N__23618\
        );

    \I__3096\ : LocalMux
    port map (
            O => \N__23624\,
            I => \N__23615\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__23621\,
            I => \N__23612\
        );

    \I__3094\ : InMux
    port map (
            O => \N__23618\,
            I => \N__23609\
        );

    \I__3093\ : Span4Mux_v
    port map (
            O => \N__23615\,
            I => \N__23606\
        );

    \I__3092\ : Span12Mux_s9_h
    port map (
            O => \N__23612\,
            I => \N__23603\
        );

    \I__3091\ : LocalMux
    port map (
            O => \N__23609\,
            I => buf_adcdata_iac_1
        );

    \I__3090\ : Odrv4
    port map (
            O => \N__23606\,
            I => buf_adcdata_iac_1
        );

    \I__3089\ : Odrv12
    port map (
            O => \N__23603\,
            I => buf_adcdata_iac_1
        );

    \I__3088\ : InMux
    port map (
            O => \N__23596\,
            I => \N__23593\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__23593\,
            I => \N__23590\
        );

    \I__3086\ : Span4Mux_v
    port map (
            O => \N__23590\,
            I => \N__23587\
        );

    \I__3085\ : Odrv4
    port map (
            O => \N__23587\,
            I => buf_data_iac_1
        );

    \I__3084\ : CascadeMux
    port map (
            O => \N__23584\,
            I => \n22_adj_1618_cascade_\
        );

    \I__3083\ : InMux
    port map (
            O => \N__23581\,
            I => \N__23578\
        );

    \I__3082\ : LocalMux
    port map (
            O => \N__23578\,
            I => \N__23574\
        );

    \I__3081\ : CascadeMux
    port map (
            O => \N__23577\,
            I => \N__23571\
        );

    \I__3080\ : Span4Mux_v
    port map (
            O => \N__23574\,
            I => \N__23568\
        );

    \I__3079\ : InMux
    port map (
            O => \N__23571\,
            I => \N__23565\
        );

    \I__3078\ : Odrv4
    port map (
            O => \N__23568\,
            I => buf_adcdata_vdc_15
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__23565\,
            I => buf_adcdata_vdc_15
        );

    \I__3076\ : InMux
    port map (
            O => \N__23560\,
            I => \N__23557\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__23557\,
            I => \N__23554\
        );

    \I__3074\ : Span4Mux_v
    port map (
            O => \N__23554\,
            I => \N__23550\
        );

    \I__3073\ : InMux
    port map (
            O => \N__23553\,
            I => \N__23547\
        );

    \I__3072\ : Odrv4
    port map (
            O => \N__23550\,
            I => buf_adcdata_vdc_14
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__23547\,
            I => buf_adcdata_vdc_14
        );

    \I__3070\ : CascadeMux
    port map (
            O => \N__23542\,
            I => \N__23538\
        );

    \I__3069\ : CascadeMux
    port map (
            O => \N__23541\,
            I => \N__23535\
        );

    \I__3068\ : InMux
    port map (
            O => \N__23538\,
            I => \N__23532\
        );

    \I__3067\ : InMux
    port map (
            O => \N__23535\,
            I => \N__23529\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__23532\,
            I => buf_adcdata_vdc_22
        );

    \I__3065\ : LocalMux
    port map (
            O => \N__23529\,
            I => buf_adcdata_vdc_22
        );

    \I__3064\ : CascadeMux
    port map (
            O => \N__23524\,
            I => \N__23520\
        );

    \I__3063\ : CascadeMux
    port map (
            O => \N__23523\,
            I => \N__23517\
        );

    \I__3062\ : InMux
    port map (
            O => \N__23520\,
            I => \N__23514\
        );

    \I__3061\ : InMux
    port map (
            O => \N__23517\,
            I => \N__23511\
        );

    \I__3060\ : LocalMux
    port map (
            O => \N__23514\,
            I => \N__23508\
        );

    \I__3059\ : LocalMux
    port map (
            O => \N__23511\,
            I => \N__23505\
        );

    \I__3058\ : Odrv4
    port map (
            O => \N__23508\,
            I => buf_adcdata_vdc_17
        );

    \I__3057\ : Odrv4
    port map (
            O => \N__23505\,
            I => buf_adcdata_vdc_17
        );

    \I__3056\ : InMux
    port map (
            O => \N__23500\,
            I => \N__23496\
        );

    \I__3055\ : CascadeMux
    port map (
            O => \N__23499\,
            I => \N__23493\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__23496\,
            I => \N__23490\
        );

    \I__3053\ : InMux
    port map (
            O => \N__23493\,
            I => \N__23487\
        );

    \I__3052\ : Odrv12
    port map (
            O => \N__23490\,
            I => buf_adcdata_vdc_0
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__23487\,
            I => buf_adcdata_vdc_0
        );

    \I__3050\ : InMux
    port map (
            O => \N__23482\,
            I => \N__23479\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__23479\,
            I => \N__23474\
        );

    \I__3048\ : InMux
    port map (
            O => \N__23478\,
            I => \N__23471\
        );

    \I__3047\ : InMux
    port map (
            O => \N__23477\,
            I => \N__23468\
        );

    \I__3046\ : Span4Mux_h
    port map (
            O => \N__23474\,
            I => \N__23463\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__23471\,
            I => \N__23463\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__23468\,
            I => buf_adcdata_vac_0
        );

    \I__3043\ : Odrv4
    port map (
            O => \N__23463\,
            I => buf_adcdata_vac_0
        );

    \I__3042\ : InMux
    port map (
            O => \N__23458\,
            I => \N__23454\
        );

    \I__3041\ : InMux
    port map (
            O => \N__23457\,
            I => \N__23451\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__23454\,
            I => \N__23447\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__23451\,
            I => \N__23444\
        );

    \I__3038\ : InMux
    port map (
            O => \N__23450\,
            I => \N__23441\
        );

    \I__3037\ : Span4Mux_v
    port map (
            O => \N__23447\,
            I => \N__23436\
        );

    \I__3036\ : Span4Mux_v
    port map (
            O => \N__23444\,
            I => \N__23436\
        );

    \I__3035\ : LocalMux
    port map (
            O => \N__23441\,
            I => buf_adcdata_iac_0
        );

    \I__3034\ : Odrv4
    port map (
            O => \N__23436\,
            I => buf_adcdata_iac_0
        );

    \I__3033\ : CascadeMux
    port map (
            O => \N__23431\,
            I => \n19_adj_1477_cascade_\
        );

    \I__3032\ : CascadeMux
    port map (
            O => \N__23428\,
            I => \N__23425\
        );

    \I__3031\ : InMux
    port map (
            O => \N__23425\,
            I => \N__23422\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__23422\,
            I => \N__23419\
        );

    \I__3029\ : Span4Mux_h
    port map (
            O => \N__23419\,
            I => \N__23416\
        );

    \I__3028\ : Span4Mux_h
    port map (
            O => \N__23416\,
            I => \N__23412\
        );

    \I__3027\ : InMux
    port map (
            O => \N__23415\,
            I => \N__23409\
        );

    \I__3026\ : Odrv4
    port map (
            O => \N__23412\,
            I => \buf_readRTD_14\
        );

    \I__3025\ : LocalMux
    port map (
            O => \N__23409\,
            I => \buf_readRTD_14\
        );

    \I__3024\ : InMux
    port map (
            O => \N__23404\,
            I => \N__23401\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__23401\,
            I => n22141
        );

    \I__3022\ : InMux
    port map (
            O => \N__23398\,
            I => \N__23395\
        );

    \I__3021\ : LocalMux
    port map (
            O => \N__23395\,
            I => \N__23392\
        );

    \I__3020\ : Span4Mux_v
    port map (
            O => \N__23392\,
            I => \N__23388\
        );

    \I__3019\ : CascadeMux
    port map (
            O => \N__23391\,
            I => \N__23385\
        );

    \I__3018\ : Span4Mux_h
    port map (
            O => \N__23388\,
            I => \N__23382\
        );

    \I__3017\ : InMux
    port map (
            O => \N__23385\,
            I => \N__23379\
        );

    \I__3016\ : Odrv4
    port map (
            O => \N__23382\,
            I => \buf_readRTD_10\
        );

    \I__3015\ : LocalMux
    port map (
            O => \N__23379\,
            I => \buf_readRTD_10\
        );

    \I__3014\ : CascadeMux
    port map (
            O => \N__23374\,
            I => \N__23371\
        );

    \I__3013\ : InMux
    port map (
            O => \N__23371\,
            I => \N__23368\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__23368\,
            I => \N__23364\
        );

    \I__3011\ : CascadeMux
    port map (
            O => \N__23367\,
            I => \N__23361\
        );

    \I__3010\ : Span4Mux_v
    port map (
            O => \N__23364\,
            I => \N__23358\
        );

    \I__3009\ : InMux
    port map (
            O => \N__23361\,
            I => \N__23355\
        );

    \I__3008\ : Odrv4
    port map (
            O => \N__23358\,
            I => buf_adcdata_vdc_21
        );

    \I__3007\ : LocalMux
    port map (
            O => \N__23355\,
            I => buf_adcdata_vdc_21
        );

    \I__3006\ : InMux
    port map (
            O => \N__23350\,
            I => \N__23347\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__23347\,
            I => \N__23344\
        );

    \I__3004\ : Span4Mux_v
    port map (
            O => \N__23344\,
            I => \N__23340\
        );

    \I__3003\ : CascadeMux
    port map (
            O => \N__23343\,
            I => \N__23337\
        );

    \I__3002\ : Span4Mux_v
    port map (
            O => \N__23340\,
            I => \N__23334\
        );

    \I__3001\ : InMux
    port map (
            O => \N__23337\,
            I => \N__23331\
        );

    \I__3000\ : Odrv4
    port map (
            O => \N__23334\,
            I => buf_adcdata_vdc_13
        );

    \I__2999\ : LocalMux
    port map (
            O => \N__23331\,
            I => buf_adcdata_vdc_13
        );

    \I__2998\ : InMux
    port map (
            O => \N__23326\,
            I => \N__23322\
        );

    \I__2997\ : CascadeMux
    port map (
            O => \N__23325\,
            I => \N__23319\
        );

    \I__2996\ : LocalMux
    port map (
            O => \N__23322\,
            I => \N__23316\
        );

    \I__2995\ : InMux
    port map (
            O => \N__23319\,
            I => \N__23313\
        );

    \I__2994\ : Odrv4
    port map (
            O => \N__23316\,
            I => buf_adcdata_vdc_16
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__23313\,
            I => buf_adcdata_vdc_16
        );

    \I__2992\ : InMux
    port map (
            O => \N__23308\,
            I => \N__23304\
        );

    \I__2991\ : CascadeMux
    port map (
            O => \N__23307\,
            I => \N__23301\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__23304\,
            I => \N__23298\
        );

    \I__2989\ : InMux
    port map (
            O => \N__23301\,
            I => \N__23295\
        );

    \I__2988\ : Odrv4
    port map (
            O => \N__23298\,
            I => buf_adcdata_vdc_2
        );

    \I__2987\ : LocalMux
    port map (
            O => \N__23295\,
            I => buf_adcdata_vdc_2
        );

    \I__2986\ : InMux
    port map (
            O => \N__23290\,
            I => \N__23287\
        );

    \I__2985\ : LocalMux
    port map (
            O => \N__23287\,
            I => \N__23283\
        );

    \I__2984\ : CascadeMux
    port map (
            O => \N__23286\,
            I => \N__23280\
        );

    \I__2983\ : Span4Mux_v
    port map (
            O => \N__23283\,
            I => \N__23277\
        );

    \I__2982\ : InMux
    port map (
            O => \N__23280\,
            I => \N__23274\
        );

    \I__2981\ : Odrv4
    port map (
            O => \N__23277\,
            I => buf_adcdata_vdc_19
        );

    \I__2980\ : LocalMux
    port map (
            O => \N__23274\,
            I => buf_adcdata_vdc_19
        );

    \I__2979\ : CEMux
    port map (
            O => \N__23269\,
            I => \N__23266\
        );

    \I__2978\ : LocalMux
    port map (
            O => \N__23266\,
            I => \N__23263\
        );

    \I__2977\ : Odrv4
    port map (
            O => \N__23263\,
            I => \CLK_DDS.n9_adj_1386\
        );

    \I__2976\ : InMux
    port map (
            O => \N__23260\,
            I => \ADC_IAC.n19355\
        );

    \I__2975\ : InMux
    port map (
            O => \N__23257\,
            I => \ADC_IAC.n19356\
        );

    \I__2974\ : CEMux
    port map (
            O => \N__23254\,
            I => \N__23251\
        );

    \I__2973\ : LocalMux
    port map (
            O => \N__23251\,
            I => \N__23248\
        );

    \I__2972\ : Span4Mux_v
    port map (
            O => \N__23248\,
            I => \N__23245\
        );

    \I__2971\ : Span4Mux_h
    port map (
            O => \N__23245\,
            I => \N__23242\
        );

    \I__2970\ : Odrv4
    port map (
            O => \N__23242\,
            I => \ADC_IAC.n12459\
        );

    \I__2969\ : SRMux
    port map (
            O => \N__23239\,
            I => \N__23236\
        );

    \I__2968\ : LocalMux
    port map (
            O => \N__23236\,
            I => \ADC_IAC.n14791\
        );

    \I__2967\ : InMux
    port map (
            O => \N__23233\,
            I => \N__23226\
        );

    \I__2966\ : InMux
    port map (
            O => \N__23232\,
            I => \N__23219\
        );

    \I__2965\ : InMux
    port map (
            O => \N__23231\,
            I => \N__23219\
        );

    \I__2964\ : InMux
    port map (
            O => \N__23230\,
            I => \N__23219\
        );

    \I__2963\ : InMux
    port map (
            O => \N__23229\,
            I => \N__23216\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__23226\,
            I => bit_cnt_0_adj_1449
        );

    \I__2961\ : LocalMux
    port map (
            O => \N__23219\,
            I => bit_cnt_0_adj_1449
        );

    \I__2960\ : LocalMux
    port map (
            O => \N__23216\,
            I => bit_cnt_0_adj_1449
        );

    \I__2959\ : CascadeMux
    port map (
            O => \N__23209\,
            I => \N__23206\
        );

    \I__2958\ : InMux
    port map (
            O => \N__23206\,
            I => \N__23202\
        );

    \I__2957\ : InMux
    port map (
            O => \N__23205\,
            I => \N__23199\
        );

    \I__2956\ : LocalMux
    port map (
            O => \N__23202\,
            I => \N__23194\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__23199\,
            I => \N__23194\
        );

    \I__2954\ : Odrv4
    port map (
            O => \N__23194\,
            I => bit_cnt_3
        );

    \I__2953\ : InMux
    port map (
            O => \N__23191\,
            I => \N__23188\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__23188\,
            I => \N__23185\
        );

    \I__2951\ : Span4Mux_v
    port map (
            O => \N__23185\,
            I => \N__23182\
        );

    \I__2950\ : Odrv4
    port map (
            O => \N__23182\,
            I => n21206
        );

    \I__2949\ : InMux
    port map (
            O => \N__23179\,
            I => \N__23176\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__23176\,
            I => \N__23173\
        );

    \I__2947\ : Span4Mux_v
    port map (
            O => \N__23173\,
            I => \N__23169\
        );

    \I__2946\ : CascadeMux
    port map (
            O => \N__23172\,
            I => \N__23166\
        );

    \I__2945\ : Span4Mux_v
    port map (
            O => \N__23169\,
            I => \N__23163\
        );

    \I__2944\ : InMux
    port map (
            O => \N__23166\,
            I => \N__23160\
        );

    \I__2943\ : Odrv4
    port map (
            O => \N__23163\,
            I => buf_adcdata_vdc_3
        );

    \I__2942\ : LocalMux
    port map (
            O => \N__23160\,
            I => buf_adcdata_vdc_3
        );

    \I__2941\ : CascadeMux
    port map (
            O => \N__23155\,
            I => \ADC_IAC.n12459_cascade_\
        );

    \I__2940\ : InMux
    port map (
            O => \N__23152\,
            I => \bfn_7_19_0_\
        );

    \I__2939\ : InMux
    port map (
            O => \N__23149\,
            I => \ADC_IAC.n19350\
        );

    \I__2938\ : InMux
    port map (
            O => \N__23146\,
            I => \ADC_IAC.n19351\
        );

    \I__2937\ : InMux
    port map (
            O => \N__23143\,
            I => \ADC_IAC.n19352\
        );

    \I__2936\ : InMux
    port map (
            O => \N__23140\,
            I => \ADC_IAC.n19353\
        );

    \I__2935\ : InMux
    port map (
            O => \N__23137\,
            I => \ADC_IAC.n19354\
        );

    \I__2934\ : InMux
    port map (
            O => \N__23134\,
            I => \N__23130\
        );

    \I__2933\ : InMux
    port map (
            O => \N__23133\,
            I => \N__23127\
        );

    \I__2932\ : LocalMux
    port map (
            O => \N__23130\,
            I => \ADC_VAC.bit_cnt_2\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__23127\,
            I => \ADC_VAC.bit_cnt_2\
        );

    \I__2930\ : InMux
    port map (
            O => \N__23122\,
            I => \ADC_VAC.n19358\
        );

    \I__2929\ : InMux
    port map (
            O => \N__23119\,
            I => \N__23115\
        );

    \I__2928\ : InMux
    port map (
            O => \N__23118\,
            I => \N__23112\
        );

    \I__2927\ : LocalMux
    port map (
            O => \N__23115\,
            I => \ADC_VAC.bit_cnt_3\
        );

    \I__2926\ : LocalMux
    port map (
            O => \N__23112\,
            I => \ADC_VAC.bit_cnt_3\
        );

    \I__2925\ : InMux
    port map (
            O => \N__23107\,
            I => \ADC_VAC.n19359\
        );

    \I__2924\ : InMux
    port map (
            O => \N__23104\,
            I => \N__23100\
        );

    \I__2923\ : InMux
    port map (
            O => \N__23103\,
            I => \N__23097\
        );

    \I__2922\ : LocalMux
    port map (
            O => \N__23100\,
            I => \N__23094\
        );

    \I__2921\ : LocalMux
    port map (
            O => \N__23097\,
            I => \ADC_VAC.bit_cnt_4\
        );

    \I__2920\ : Odrv4
    port map (
            O => \N__23094\,
            I => \ADC_VAC.bit_cnt_4\
        );

    \I__2919\ : InMux
    port map (
            O => \N__23089\,
            I => \ADC_VAC.n19360\
        );

    \I__2918\ : InMux
    port map (
            O => \N__23086\,
            I => \N__23082\
        );

    \I__2917\ : InMux
    port map (
            O => \N__23085\,
            I => \N__23079\
        );

    \I__2916\ : LocalMux
    port map (
            O => \N__23082\,
            I => \ADC_VAC.bit_cnt_5\
        );

    \I__2915\ : LocalMux
    port map (
            O => \N__23079\,
            I => \ADC_VAC.bit_cnt_5\
        );

    \I__2914\ : InMux
    port map (
            O => \N__23074\,
            I => \ADC_VAC.n19361\
        );

    \I__2913\ : InMux
    port map (
            O => \N__23071\,
            I => \N__23067\
        );

    \I__2912\ : InMux
    port map (
            O => \N__23070\,
            I => \N__23064\
        );

    \I__2911\ : LocalMux
    port map (
            O => \N__23067\,
            I => \ADC_VAC.bit_cnt_6\
        );

    \I__2910\ : LocalMux
    port map (
            O => \N__23064\,
            I => \ADC_VAC.bit_cnt_6\
        );

    \I__2909\ : InMux
    port map (
            O => \N__23059\,
            I => \ADC_VAC.n19362\
        );

    \I__2908\ : InMux
    port map (
            O => \N__23056\,
            I => \ADC_VAC.n19363\
        );

    \I__2907\ : InMux
    port map (
            O => \N__23053\,
            I => \N__23049\
        );

    \I__2906\ : InMux
    port map (
            O => \N__23052\,
            I => \N__23046\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__23049\,
            I => \ADC_VAC.bit_cnt_7\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__23046\,
            I => \ADC_VAC.bit_cnt_7\
        );

    \I__2903\ : CEMux
    port map (
            O => \N__23041\,
            I => \N__23038\
        );

    \I__2902\ : LocalMux
    port map (
            O => \N__23038\,
            I => \N__23035\
        );

    \I__2901\ : Span4Mux_v
    port map (
            O => \N__23035\,
            I => \N__23032\
        );

    \I__2900\ : Odrv4
    port map (
            O => \N__23032\,
            I => \ADC_VAC.n12556\
        );

    \I__2899\ : SRMux
    port map (
            O => \N__23029\,
            I => \N__23026\
        );

    \I__2898\ : LocalMux
    port map (
            O => \N__23026\,
            I => \N__23023\
        );

    \I__2897\ : Span4Mux_v
    port map (
            O => \N__23023\,
            I => \N__23020\
        );

    \I__2896\ : Odrv4
    port map (
            O => \N__23020\,
            I => \ADC_VAC.n14829\
        );

    \I__2895\ : CascadeMux
    port map (
            O => \N__23017\,
            I => \ADC_VAC.n20747_cascade_\
        );

    \I__2894\ : CascadeMux
    port map (
            O => \N__23014\,
            I => \ADC_VAC.n20763_cascade_\
        );

    \I__2893\ : CascadeMux
    port map (
            O => \N__23011\,
            I => \ADC_VAC.n21031_cascade_\
        );

    \I__2892\ : CEMux
    port map (
            O => \N__23008\,
            I => \N__23005\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__23005\,
            I => \N__23002\
        );

    \I__2890\ : Odrv4
    port map (
            O => \N__23002\,
            I => \ADC_VAC.n20668\
        );

    \I__2889\ : CascadeMux
    port map (
            O => \N__22999\,
            I => \N__22995\
        );

    \I__2888\ : InMux
    port map (
            O => \N__22998\,
            I => \N__22988\
        );

    \I__2887\ : InMux
    port map (
            O => \N__22995\,
            I => \N__22988\
        );

    \I__2886\ : InMux
    port map (
            O => \N__22994\,
            I => \N__22983\
        );

    \I__2885\ : InMux
    port map (
            O => \N__22993\,
            I => \N__22983\
        );

    \I__2884\ : LocalMux
    port map (
            O => \N__22988\,
            I => \N__22977\
        );

    \I__2883\ : LocalMux
    port map (
            O => \N__22983\,
            I => \N__22977\
        );

    \I__2882\ : InMux
    port map (
            O => \N__22982\,
            I => \N__22974\
        );

    \I__2881\ : Span4Mux_v
    port map (
            O => \N__22977\,
            I => \N__22971\
        );

    \I__2880\ : LocalMux
    port map (
            O => \N__22974\,
            I => \N__22968\
        );

    \I__2879\ : Span4Mux_h
    port map (
            O => \N__22971\,
            I => \N__22965\
        );

    \I__2878\ : Span4Mux_v
    port map (
            O => \N__22968\,
            I => \N__22962\
        );

    \I__2877\ : Sp12to4
    port map (
            O => \N__22965\,
            I => \N__22957\
        );

    \I__2876\ : Sp12to4
    port map (
            O => \N__22962\,
            I => \N__22957\
        );

    \I__2875\ : Odrv12
    port map (
            O => \N__22957\,
            I => \VAC_DRDY\
        );

    \I__2874\ : CascadeMux
    port map (
            O => \N__22954\,
            I => \ADC_VAC.n17_cascade_\
        );

    \I__2873\ : CEMux
    port map (
            O => \N__22951\,
            I => \N__22948\
        );

    \I__2872\ : LocalMux
    port map (
            O => \N__22948\,
            I => \N__22945\
        );

    \I__2871\ : Odrv4
    port map (
            O => \N__22945\,
            I => \ADC_VAC.n12\
        );

    \I__2870\ : InMux
    port map (
            O => \N__22942\,
            I => \N__22938\
        );

    \I__2869\ : InMux
    port map (
            O => \N__22941\,
            I => \N__22935\
        );

    \I__2868\ : LocalMux
    port map (
            O => \N__22938\,
            I => \ADC_VAC.bit_cnt_0\
        );

    \I__2867\ : LocalMux
    port map (
            O => \N__22935\,
            I => \ADC_VAC.bit_cnt_0\
        );

    \I__2866\ : InMux
    port map (
            O => \N__22930\,
            I => \bfn_7_17_0_\
        );

    \I__2865\ : CascadeMux
    port map (
            O => \N__22927\,
            I => \N__22923\
        );

    \I__2864\ : InMux
    port map (
            O => \N__22926\,
            I => \N__22920\
        );

    \I__2863\ : InMux
    port map (
            O => \N__22923\,
            I => \N__22917\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__22920\,
            I => \ADC_VAC.bit_cnt_1\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__22917\,
            I => \ADC_VAC.bit_cnt_1\
        );

    \I__2860\ : InMux
    port map (
            O => \N__22912\,
            I => \ADC_VAC.n19357\
        );

    \I__2859\ : CascadeMux
    port map (
            O => \N__22909\,
            I => \N__22906\
        );

    \I__2858\ : InMux
    port map (
            O => \N__22906\,
            I => \N__22900\
        );

    \I__2857\ : InMux
    port map (
            O => \N__22905\,
            I => \N__22900\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__22900\,
            I => cmd_rdadctmp_0_adj_1443
        );

    \I__2855\ : InMux
    port map (
            O => \N__22897\,
            I => \N__22891\
        );

    \I__2854\ : InMux
    port map (
            O => \N__22896\,
            I => \N__22891\
        );

    \I__2853\ : LocalMux
    port map (
            O => \N__22891\,
            I => cmd_rdadctmp_1_adj_1442
        );

    \I__2852\ : InMux
    port map (
            O => \N__22888\,
            I => \N__22882\
        );

    \I__2851\ : InMux
    port map (
            O => \N__22887\,
            I => \N__22882\
        );

    \I__2850\ : LocalMux
    port map (
            O => \N__22882\,
            I => cmd_rdadctmp_2_adj_1441
        );

    \I__2849\ : CascadeMux
    port map (
            O => \N__22879\,
            I => \N__22876\
        );

    \I__2848\ : InMux
    port map (
            O => \N__22876\,
            I => \N__22872\
        );

    \I__2847\ : InMux
    port map (
            O => \N__22875\,
            I => \N__22869\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__22872\,
            I => cmd_rdadctmp_3_adj_1440
        );

    \I__2845\ : LocalMux
    port map (
            O => \N__22869\,
            I => cmd_rdadctmp_3_adj_1440
        );

    \I__2844\ : InMux
    port map (
            O => \N__22864\,
            I => \N__22861\
        );

    \I__2843\ : LocalMux
    port map (
            O => \N__22861\,
            I => \N__22858\
        );

    \I__2842\ : Odrv12
    port map (
            O => \N__22858\,
            I => n20573
        );

    \I__2841\ : CascadeMux
    port map (
            O => \N__22855\,
            I => \ADC_VAC.n12556_cascade_\
        );

    \I__2840\ : InMux
    port map (
            O => \N__22852\,
            I => \N__22849\
        );

    \I__2839\ : LocalMux
    port map (
            O => \N__22849\,
            I => \ADC_VAC.n20667\
        );

    \I__2838\ : CascadeMux
    port map (
            O => \N__22846\,
            I => \N__22842\
        );

    \I__2837\ : CascadeMux
    port map (
            O => \N__22845\,
            I => \N__22839\
        );

    \I__2836\ : InMux
    port map (
            O => \N__22842\,
            I => \N__22835\
        );

    \I__2835\ : InMux
    port map (
            O => \N__22839\,
            I => \N__22830\
        );

    \I__2834\ : InMux
    port map (
            O => \N__22838\,
            I => \N__22830\
        );

    \I__2833\ : LocalMux
    port map (
            O => \N__22835\,
            I => cmd_rdadctmp_11_adj_1432
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__22830\,
            I => cmd_rdadctmp_11_adj_1432
        );

    \I__2831\ : InMux
    port map (
            O => \N__22825\,
            I => \N__22822\
        );

    \I__2830\ : LocalMux
    port map (
            O => \N__22822\,
            I => \N__22819\
        );

    \I__2829\ : Span4Mux_v
    port map (
            O => \N__22819\,
            I => \N__22815\
        );

    \I__2828\ : InMux
    port map (
            O => \N__22818\,
            I => \N__22812\
        );

    \I__2827\ : Odrv4
    port map (
            O => \N__22815\,
            I => cmd_rdadctmp_7_adj_1436
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__22812\,
            I => cmd_rdadctmp_7_adj_1436
        );

    \I__2825\ : CascadeMux
    port map (
            O => \N__22807\,
            I => \N__22804\
        );

    \I__2824\ : InMux
    port map (
            O => \N__22804\,
            I => \N__22800\
        );

    \I__2823\ : CascadeMux
    port map (
            O => \N__22803\,
            I => \N__22797\
        );

    \I__2822\ : LocalMux
    port map (
            O => \N__22800\,
            I => \N__22793\
        );

    \I__2821\ : InMux
    port map (
            O => \N__22797\,
            I => \N__22788\
        );

    \I__2820\ : InMux
    port map (
            O => \N__22796\,
            I => \N__22788\
        );

    \I__2819\ : Odrv4
    port map (
            O => \N__22793\,
            I => cmd_rdadctmp_8_adj_1435
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__22788\,
            I => cmd_rdadctmp_8_adj_1435
        );

    \I__2817\ : CascadeMux
    port map (
            O => \N__22783\,
            I => \N__22779\
        );

    \I__2816\ : CascadeMux
    port map (
            O => \N__22782\,
            I => \N__22776\
        );

    \I__2815\ : InMux
    port map (
            O => \N__22779\,
            I => \N__22768\
        );

    \I__2814\ : InMux
    port map (
            O => \N__22776\,
            I => \N__22768\
        );

    \I__2813\ : InMux
    port map (
            O => \N__22775\,
            I => \N__22768\
        );

    \I__2812\ : LocalMux
    port map (
            O => \N__22768\,
            I => cmd_rdadctmp_9_adj_1434
        );

    \I__2811\ : CascadeMux
    port map (
            O => \N__22765\,
            I => \N__22762\
        );

    \I__2810\ : InMux
    port map (
            O => \N__22762\,
            I => \N__22759\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__22759\,
            I => \N__22756\
        );

    \I__2808\ : Span4Mux_h
    port map (
            O => \N__22756\,
            I => \N__22753\
        );

    \I__2807\ : Sp12to4
    port map (
            O => \N__22753\,
            I => \N__22750\
        );

    \I__2806\ : Odrv12
    port map (
            O => \N__22750\,
            I => \VAC_MISO\
        );

    \I__2805\ : InMux
    port map (
            O => \N__22747\,
            I => \N__22744\
        );

    \I__2804\ : LocalMux
    port map (
            O => \N__22744\,
            I => n21973
        );

    \I__2803\ : InMux
    port map (
            O => \N__22741\,
            I => \N__22734\
        );

    \I__2802\ : InMux
    port map (
            O => \N__22740\,
            I => \N__22734\
        );

    \I__2801\ : InMux
    port map (
            O => \N__22739\,
            I => \N__22731\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__22734\,
            I => cmd_rdadctmp_17_adj_1426
        );

    \I__2799\ : LocalMux
    port map (
            O => \N__22731\,
            I => cmd_rdadctmp_17_adj_1426
        );

    \I__2798\ : InMux
    port map (
            O => \N__22726\,
            I => \N__22721\
        );

    \I__2797\ : InMux
    port map (
            O => \N__22725\,
            I => \N__22716\
        );

    \I__2796\ : InMux
    port map (
            O => \N__22724\,
            I => \N__22716\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__22721\,
            I => cmd_rdadctmp_16_adj_1427
        );

    \I__2794\ : LocalMux
    port map (
            O => \N__22716\,
            I => cmd_rdadctmp_16_adj_1427
        );

    \I__2793\ : InMux
    port map (
            O => \N__22711\,
            I => \N__22708\
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__22708\,
            I => \N__22705\
        );

    \I__2791\ : Span4Mux_h
    port map (
            O => \N__22705\,
            I => \N__22700\
        );

    \I__2790\ : InMux
    port map (
            O => \N__22704\,
            I => \N__22697\
        );

    \I__2789\ : InMux
    port map (
            O => \N__22703\,
            I => \N__22694\
        );

    \I__2788\ : Sp12to4
    port map (
            O => \N__22700\,
            I => \N__22691\
        );

    \I__2787\ : LocalMux
    port map (
            O => \N__22697\,
            I => \N__22688\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__22694\,
            I => buf_adcdata_vac_22
        );

    \I__2785\ : Odrv12
    port map (
            O => \N__22691\,
            I => buf_adcdata_vac_22
        );

    \I__2784\ : Odrv4
    port map (
            O => \N__22688\,
            I => buf_adcdata_vac_22
        );

    \I__2783\ : InMux
    port map (
            O => \N__22681\,
            I => \N__22678\
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__22678\,
            I => \N__22674\
        );

    \I__2781\ : InMux
    port map (
            O => \N__22677\,
            I => \N__22670\
        );

    \I__2780\ : Span4Mux_v
    port map (
            O => \N__22674\,
            I => \N__22667\
        );

    \I__2779\ : InMux
    port map (
            O => \N__22673\,
            I => \N__22664\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__22670\,
            I => buf_adcdata_vac_14
        );

    \I__2777\ : Odrv4
    port map (
            O => \N__22667\,
            I => buf_adcdata_vac_14
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__22664\,
            I => buf_adcdata_vac_14
        );

    \I__2775\ : InMux
    port map (
            O => \N__22657\,
            I => \N__22653\
        );

    \I__2774\ : CascadeMux
    port map (
            O => \N__22656\,
            I => \N__22649\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__22653\,
            I => \N__22646\
        );

    \I__2772\ : InMux
    port map (
            O => \N__22652\,
            I => \N__22643\
        );

    \I__2771\ : InMux
    port map (
            O => \N__22649\,
            I => \N__22640\
        );

    \I__2770\ : Span4Mux_h
    port map (
            O => \N__22646\,
            I => \N__22637\
        );

    \I__2769\ : LocalMux
    port map (
            O => \N__22643\,
            I => \N__22634\
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__22640\,
            I => buf_adcdata_vac_17
        );

    \I__2767\ : Odrv4
    port map (
            O => \N__22637\,
            I => buf_adcdata_vac_17
        );

    \I__2766\ : Odrv12
    port map (
            O => \N__22634\,
            I => buf_adcdata_vac_17
        );

    \I__2765\ : CascadeMux
    port map (
            O => \N__22627\,
            I => \N__22623\
        );

    \I__2764\ : CascadeMux
    port map (
            O => \N__22626\,
            I => \N__22620\
        );

    \I__2763\ : InMux
    port map (
            O => \N__22623\,
            I => \N__22614\
        );

    \I__2762\ : InMux
    port map (
            O => \N__22620\,
            I => \N__22614\
        );

    \I__2761\ : InMux
    port map (
            O => \N__22619\,
            I => \N__22611\
        );

    \I__2760\ : LocalMux
    port map (
            O => \N__22614\,
            I => cmd_rdadctmp_30_adj_1413
        );

    \I__2759\ : LocalMux
    port map (
            O => \N__22611\,
            I => cmd_rdadctmp_30_adj_1413
        );

    \I__2758\ : InMux
    port map (
            O => \N__22606\,
            I => \N__22600\
        );

    \I__2757\ : InMux
    port map (
            O => \N__22605\,
            I => \N__22600\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__22600\,
            I => cmd_rdadctmp_31_adj_1412
        );

    \I__2755\ : CascadeMux
    port map (
            O => \N__22597\,
            I => \N__22592\
        );

    \I__2754\ : InMux
    port map (
            O => \N__22596\,
            I => \N__22589\
        );

    \I__2753\ : InMux
    port map (
            O => \N__22595\,
            I => \N__22586\
        );

    \I__2752\ : InMux
    port map (
            O => \N__22592\,
            I => \N__22583\
        );

    \I__2751\ : LocalMux
    port map (
            O => \N__22589\,
            I => \N__22580\
        );

    \I__2750\ : LocalMux
    port map (
            O => \N__22586\,
            I => \N__22577\
        );

    \I__2749\ : LocalMux
    port map (
            O => \N__22583\,
            I => buf_adcdata_vac_16
        );

    \I__2748\ : Odrv4
    port map (
            O => \N__22580\,
            I => buf_adcdata_vac_16
        );

    \I__2747\ : Odrv12
    port map (
            O => \N__22577\,
            I => buf_adcdata_vac_16
        );

    \I__2746\ : CascadeMux
    port map (
            O => \N__22570\,
            I => \N__22567\
        );

    \I__2745\ : InMux
    port map (
            O => \N__22567\,
            I => \N__22563\
        );

    \I__2744\ : CascadeMux
    port map (
            O => \N__22566\,
            I => \N__22560\
        );

    \I__2743\ : LocalMux
    port map (
            O => \N__22563\,
            I => \N__22556\
        );

    \I__2742\ : InMux
    port map (
            O => \N__22560\,
            I => \N__22553\
        );

    \I__2741\ : InMux
    port map (
            O => \N__22559\,
            I => \N__22550\
        );

    \I__2740\ : Odrv12
    port map (
            O => \N__22556\,
            I => cmd_rdadctmp_10_adj_1433
        );

    \I__2739\ : LocalMux
    port map (
            O => \N__22553\,
            I => cmd_rdadctmp_10_adj_1433
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__22550\,
            I => cmd_rdadctmp_10_adj_1433
        );

    \I__2737\ : CascadeMux
    port map (
            O => \N__22543\,
            I => \n22183_cascade_\
        );

    \I__2736\ : CascadeMux
    port map (
            O => \N__22540\,
            I => \N__22537\
        );

    \I__2735\ : InMux
    port map (
            O => \N__22537\,
            I => \N__22534\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__22534\,
            I => \N__22531\
        );

    \I__2733\ : Span4Mux_v
    port map (
            O => \N__22531\,
            I => \N__22528\
        );

    \I__2732\ : Odrv4
    port map (
            O => \N__22528\,
            I => buf_data_iac_2
        );

    \I__2731\ : CascadeMux
    port map (
            O => \N__22525\,
            I => \N__22522\
        );

    \I__2730\ : InMux
    port map (
            O => \N__22522\,
            I => \N__22519\
        );

    \I__2729\ : LocalMux
    port map (
            O => \N__22519\,
            I => \N__22515\
        );

    \I__2728\ : CascadeMux
    port map (
            O => \N__22518\,
            I => \N__22512\
        );

    \I__2727\ : Span4Mux_v
    port map (
            O => \N__22515\,
            I => \N__22509\
        );

    \I__2726\ : InMux
    port map (
            O => \N__22512\,
            I => \N__22506\
        );

    \I__2725\ : Odrv4
    port map (
            O => \N__22509\,
            I => \buf_readRTD_13\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__22506\,
            I => \buf_readRTD_13\
        );

    \I__2723\ : InMux
    port map (
            O => \N__22501\,
            I => \N__22498\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__22498\,
            I => n22153
        );

    \I__2721\ : InMux
    port map (
            O => \N__22495\,
            I => \N__22492\
        );

    \I__2720\ : LocalMux
    port map (
            O => \N__22492\,
            I => \N__22487\
        );

    \I__2719\ : InMux
    port map (
            O => \N__22491\,
            I => \N__22484\
        );

    \I__2718\ : InMux
    port map (
            O => \N__22490\,
            I => \N__22481\
        );

    \I__2717\ : Span4Mux_v
    port map (
            O => \N__22487\,
            I => \N__22478\
        );

    \I__2716\ : LocalMux
    port map (
            O => \N__22484\,
            I => \N__22475\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__22481\,
            I => buf_adcdata_iac_2
        );

    \I__2714\ : Odrv4
    port map (
            O => \N__22478\,
            I => buf_adcdata_iac_2
        );

    \I__2713\ : Odrv12
    port map (
            O => \N__22475\,
            I => buf_adcdata_iac_2
        );

    \I__2712\ : CascadeMux
    port map (
            O => \N__22468\,
            I => \n19_adj_1613_cascade_\
        );

    \I__2711\ : InMux
    port map (
            O => \N__22465\,
            I => \N__22462\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__22462\,
            I => n22_adj_1614
        );

    \I__2709\ : CascadeMux
    port map (
            O => \N__22459\,
            I => \N__22456\
        );

    \I__2708\ : InMux
    port map (
            O => \N__22456\,
            I => \N__22453\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__22453\,
            I => \N__22449\
        );

    \I__2706\ : CascadeMux
    port map (
            O => \N__22452\,
            I => \N__22446\
        );

    \I__2705\ : Span4Mux_v
    port map (
            O => \N__22449\,
            I => \N__22443\
        );

    \I__2704\ : InMux
    port map (
            O => \N__22446\,
            I => \N__22440\
        );

    \I__2703\ : Odrv4
    port map (
            O => \N__22443\,
            I => \buf_readRTD_15\
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__22440\,
            I => \buf_readRTD_15\
        );

    \I__2701\ : InMux
    port map (
            O => \N__22435\,
            I => \N__22432\
        );

    \I__2700\ : LocalMux
    port map (
            O => \N__22432\,
            I => \N__22429\
        );

    \I__2699\ : Span4Mux_h
    port map (
            O => \N__22429\,
            I => \N__22426\
        );

    \I__2698\ : Span4Mux_v
    port map (
            O => \N__22426\,
            I => \N__22421\
        );

    \I__2697\ : InMux
    port map (
            O => \N__22425\,
            I => \N__22416\
        );

    \I__2696\ : InMux
    port map (
            O => \N__22424\,
            I => \N__22416\
        );

    \I__2695\ : Odrv4
    port map (
            O => \N__22421\,
            I => buf_adcdata_vac_2
        );

    \I__2694\ : LocalMux
    port map (
            O => \N__22416\,
            I => buf_adcdata_vac_2
        );

    \I__2693\ : CascadeMux
    port map (
            O => \N__22411\,
            I => \N__22405\
        );

    \I__2692\ : CascadeMux
    port map (
            O => \N__22410\,
            I => \N__22399\
        );

    \I__2691\ : CascadeMux
    port map (
            O => \N__22409\,
            I => \N__22396\
        );

    \I__2690\ : CascadeMux
    port map (
            O => \N__22408\,
            I => \N__22390\
        );

    \I__2689\ : InMux
    port map (
            O => \N__22405\,
            I => \N__22384\
        );

    \I__2688\ : InMux
    port map (
            O => \N__22404\,
            I => \N__22381\
        );

    \I__2687\ : InMux
    port map (
            O => \N__22403\,
            I => \N__22378\
        );

    \I__2686\ : CascadeMux
    port map (
            O => \N__22402\,
            I => \N__22375\
        );

    \I__2685\ : InMux
    port map (
            O => \N__22399\,
            I => \N__22362\
        );

    \I__2684\ : InMux
    port map (
            O => \N__22396\,
            I => \N__22362\
        );

    \I__2683\ : InMux
    port map (
            O => \N__22395\,
            I => \N__22362\
        );

    \I__2682\ : InMux
    port map (
            O => \N__22394\,
            I => \N__22362\
        );

    \I__2681\ : InMux
    port map (
            O => \N__22393\,
            I => \N__22362\
        );

    \I__2680\ : InMux
    port map (
            O => \N__22390\,
            I => \N__22362\
        );

    \I__2679\ : CascadeMux
    port map (
            O => \N__22389\,
            I => \N__22356\
        );

    \I__2678\ : InMux
    port map (
            O => \N__22388\,
            I => \N__22345\
        );

    \I__2677\ : InMux
    port map (
            O => \N__22387\,
            I => \N__22345\
        );

    \I__2676\ : LocalMux
    port map (
            O => \N__22384\,
            I => \N__22342\
        );

    \I__2675\ : LocalMux
    port map (
            O => \N__22381\,
            I => \N__22337\
        );

    \I__2674\ : LocalMux
    port map (
            O => \N__22378\,
            I => \N__22337\
        );

    \I__2673\ : InMux
    port map (
            O => \N__22375\,
            I => \N__22334\
        );

    \I__2672\ : LocalMux
    port map (
            O => \N__22362\,
            I => \N__22330\
        );

    \I__2671\ : InMux
    port map (
            O => \N__22361\,
            I => \N__22325\
        );

    \I__2670\ : InMux
    port map (
            O => \N__22360\,
            I => \N__22325\
        );

    \I__2669\ : InMux
    port map (
            O => \N__22359\,
            I => \N__22316\
        );

    \I__2668\ : InMux
    port map (
            O => \N__22356\,
            I => \N__22316\
        );

    \I__2667\ : InMux
    port map (
            O => \N__22355\,
            I => \N__22316\
        );

    \I__2666\ : InMux
    port map (
            O => \N__22354\,
            I => \N__22313\
        );

    \I__2665\ : InMux
    port map (
            O => \N__22353\,
            I => \N__22310\
        );

    \I__2664\ : InMux
    port map (
            O => \N__22352\,
            I => \N__22303\
        );

    \I__2663\ : InMux
    port map (
            O => \N__22351\,
            I => \N__22303\
        );

    \I__2662\ : InMux
    port map (
            O => \N__22350\,
            I => \N__22303\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__22345\,
            I => \N__22294\
        );

    \I__2660\ : Span4Mux_h
    port map (
            O => \N__22342\,
            I => \N__22294\
        );

    \I__2659\ : Span4Mux_v
    port map (
            O => \N__22337\,
            I => \N__22294\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__22334\,
            I => \N__22294\
        );

    \I__2657\ : InMux
    port map (
            O => \N__22333\,
            I => \N__22291\
        );

    \I__2656\ : Span4Mux_h
    port map (
            O => \N__22330\,
            I => \N__22286\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__22325\,
            I => \N__22286\
        );

    \I__2654\ : InMux
    port map (
            O => \N__22324\,
            I => \N__22281\
        );

    \I__2653\ : InMux
    port map (
            O => \N__22323\,
            I => \N__22281\
        );

    \I__2652\ : LocalMux
    port map (
            O => \N__22316\,
            I => \N__22278\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__22313\,
            I => \RTD.adc_state_3\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__22310\,
            I => \RTD.adc_state_3\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__22303\,
            I => \RTD.adc_state_3\
        );

    \I__2648\ : Odrv4
    port map (
            O => \N__22294\,
            I => \RTD.adc_state_3\
        );

    \I__2647\ : LocalMux
    port map (
            O => \N__22291\,
            I => \RTD.adc_state_3\
        );

    \I__2646\ : Odrv4
    port map (
            O => \N__22286\,
            I => \RTD.adc_state_3\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__22281\,
            I => \RTD.adc_state_3\
        );

    \I__2644\ : Odrv4
    port map (
            O => \N__22278\,
            I => \RTD.adc_state_3\
        );

    \I__2643\ : CascadeMux
    port map (
            O => \N__22261\,
            I => \N__22249\
        );

    \I__2642\ : InMux
    port map (
            O => \N__22260\,
            I => \N__22243\
        );

    \I__2641\ : InMux
    port map (
            O => \N__22259\,
            I => \N__22240\
        );

    \I__2640\ : InMux
    port map (
            O => \N__22258\,
            I => \N__22237\
        );

    \I__2639\ : InMux
    port map (
            O => \N__22257\,
            I => \N__22224\
        );

    \I__2638\ : InMux
    port map (
            O => \N__22256\,
            I => \N__22224\
        );

    \I__2637\ : InMux
    port map (
            O => \N__22255\,
            I => \N__22224\
        );

    \I__2636\ : InMux
    port map (
            O => \N__22254\,
            I => \N__22224\
        );

    \I__2635\ : InMux
    port map (
            O => \N__22253\,
            I => \N__22224\
        );

    \I__2634\ : InMux
    port map (
            O => \N__22252\,
            I => \N__22224\
        );

    \I__2633\ : InMux
    port map (
            O => \N__22249\,
            I => \N__22212\
        );

    \I__2632\ : InMux
    port map (
            O => \N__22248\,
            I => \N__22212\
        );

    \I__2631\ : InMux
    port map (
            O => \N__22247\,
            I => \N__22212\
        );

    \I__2630\ : InMux
    port map (
            O => \N__22246\,
            I => \N__22209\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__22243\,
            I => \N__22204\
        );

    \I__2628\ : LocalMux
    port map (
            O => \N__22240\,
            I => \N__22204\
        );

    \I__2627\ : LocalMux
    port map (
            O => \N__22237\,
            I => \N__22199\
        );

    \I__2626\ : LocalMux
    port map (
            O => \N__22224\,
            I => \N__22199\
        );

    \I__2625\ : InMux
    port map (
            O => \N__22223\,
            I => \N__22196\
        );

    \I__2624\ : InMux
    port map (
            O => \N__22222\,
            I => \N__22187\
        );

    \I__2623\ : InMux
    port map (
            O => \N__22221\,
            I => \N__22182\
        );

    \I__2622\ : InMux
    port map (
            O => \N__22220\,
            I => \N__22182\
        );

    \I__2621\ : InMux
    port map (
            O => \N__22219\,
            I => \N__22179\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__22212\,
            I => \N__22176\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__22209\,
            I => \N__22169\
        );

    \I__2618\ : Span4Mux_v
    port map (
            O => \N__22204\,
            I => \N__22169\
        );

    \I__2617\ : Span4Mux_v
    port map (
            O => \N__22199\,
            I => \N__22169\
        );

    \I__2616\ : LocalMux
    port map (
            O => \N__22196\,
            I => \N__22166\
        );

    \I__2615\ : InMux
    port map (
            O => \N__22195\,
            I => \N__22163\
        );

    \I__2614\ : InMux
    port map (
            O => \N__22194\,
            I => \N__22158\
        );

    \I__2613\ : InMux
    port map (
            O => \N__22193\,
            I => \N__22158\
        );

    \I__2612\ : InMux
    port map (
            O => \N__22192\,
            I => \N__22151\
        );

    \I__2611\ : InMux
    port map (
            O => \N__22191\,
            I => \N__22151\
        );

    \I__2610\ : InMux
    port map (
            O => \N__22190\,
            I => \N__22151\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__22187\,
            I => \RTD.adc_state_1\
        );

    \I__2608\ : LocalMux
    port map (
            O => \N__22182\,
            I => \RTD.adc_state_1\
        );

    \I__2607\ : LocalMux
    port map (
            O => \N__22179\,
            I => \RTD.adc_state_1\
        );

    \I__2606\ : Odrv4
    port map (
            O => \N__22176\,
            I => \RTD.adc_state_1\
        );

    \I__2605\ : Odrv4
    port map (
            O => \N__22169\,
            I => \RTD.adc_state_1\
        );

    \I__2604\ : Odrv4
    port map (
            O => \N__22166\,
            I => \RTD.adc_state_1\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__22163\,
            I => \RTD.adc_state_1\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__22158\,
            I => \RTD.adc_state_1\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__22151\,
            I => \RTD.adc_state_1\
        );

    \I__2600\ : CascadeMux
    port map (
            O => \N__22132\,
            I => \N__22110\
        );

    \I__2599\ : CascadeMux
    port map (
            O => \N__22131\,
            I => \N__22106\
        );

    \I__2598\ : CascadeMux
    port map (
            O => \N__22130\,
            I => \N__22096\
        );

    \I__2597\ : InMux
    port map (
            O => \N__22129\,
            I => \N__22088\
        );

    \I__2596\ : InMux
    port map (
            O => \N__22128\,
            I => \N__22088\
        );

    \I__2595\ : InMux
    port map (
            O => \N__22127\,
            I => \N__22085\
        );

    \I__2594\ : InMux
    port map (
            O => \N__22126\,
            I => \N__22076\
        );

    \I__2593\ : InMux
    port map (
            O => \N__22125\,
            I => \N__22076\
        );

    \I__2592\ : InMux
    port map (
            O => \N__22124\,
            I => \N__22076\
        );

    \I__2591\ : InMux
    port map (
            O => \N__22123\,
            I => \N__22076\
        );

    \I__2590\ : InMux
    port map (
            O => \N__22122\,
            I => \N__22069\
        );

    \I__2589\ : InMux
    port map (
            O => \N__22121\,
            I => \N__22069\
        );

    \I__2588\ : InMux
    port map (
            O => \N__22120\,
            I => \N__22069\
        );

    \I__2587\ : InMux
    port map (
            O => \N__22119\,
            I => \N__22064\
        );

    \I__2586\ : InMux
    port map (
            O => \N__22118\,
            I => \N__22064\
        );

    \I__2585\ : InMux
    port map (
            O => \N__22117\,
            I => \N__22057\
        );

    \I__2584\ : InMux
    port map (
            O => \N__22116\,
            I => \N__22057\
        );

    \I__2583\ : InMux
    port map (
            O => \N__22115\,
            I => \N__22057\
        );

    \I__2582\ : InMux
    port map (
            O => \N__22114\,
            I => \N__22044\
        );

    \I__2581\ : InMux
    port map (
            O => \N__22113\,
            I => \N__22044\
        );

    \I__2580\ : InMux
    port map (
            O => \N__22110\,
            I => \N__22044\
        );

    \I__2579\ : InMux
    port map (
            O => \N__22109\,
            I => \N__22044\
        );

    \I__2578\ : InMux
    port map (
            O => \N__22106\,
            I => \N__22044\
        );

    \I__2577\ : InMux
    port map (
            O => \N__22105\,
            I => \N__22044\
        );

    \I__2576\ : InMux
    port map (
            O => \N__22104\,
            I => \N__22041\
        );

    \I__2575\ : InMux
    port map (
            O => \N__22103\,
            I => \N__22038\
        );

    \I__2574\ : InMux
    port map (
            O => \N__22102\,
            I => \N__22027\
        );

    \I__2573\ : InMux
    port map (
            O => \N__22101\,
            I => \N__22018\
        );

    \I__2572\ : InMux
    port map (
            O => \N__22100\,
            I => \N__22018\
        );

    \I__2571\ : InMux
    port map (
            O => \N__22099\,
            I => \N__22018\
        );

    \I__2570\ : InMux
    port map (
            O => \N__22096\,
            I => \N__22015\
        );

    \I__2569\ : InMux
    port map (
            O => \N__22095\,
            I => \N__22008\
        );

    \I__2568\ : InMux
    port map (
            O => \N__22094\,
            I => \N__22008\
        );

    \I__2567\ : InMux
    port map (
            O => \N__22093\,
            I => \N__22008\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__22088\,
            I => \N__21999\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__22085\,
            I => \N__21999\
        );

    \I__2564\ : LocalMux
    port map (
            O => \N__22076\,
            I => \N__21999\
        );

    \I__2563\ : LocalMux
    port map (
            O => \N__22069\,
            I => \N__21999\
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__22064\,
            I => \N__21992\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__22057\,
            I => \N__21992\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__22044\,
            I => \N__21992\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__22041\,
            I => \N__21984\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__22038\,
            I => \N__21984\
        );

    \I__2557\ : InMux
    port map (
            O => \N__22037\,
            I => \N__21968\
        );

    \I__2556\ : InMux
    port map (
            O => \N__22036\,
            I => \N__21968\
        );

    \I__2555\ : InMux
    port map (
            O => \N__22035\,
            I => \N__21968\
        );

    \I__2554\ : InMux
    port map (
            O => \N__22034\,
            I => \N__21968\
        );

    \I__2553\ : InMux
    port map (
            O => \N__22033\,
            I => \N__21968\
        );

    \I__2552\ : InMux
    port map (
            O => \N__22032\,
            I => \N__21968\
        );

    \I__2551\ : InMux
    port map (
            O => \N__22031\,
            I => \N__21968\
        );

    \I__2550\ : InMux
    port map (
            O => \N__22030\,
            I => \N__21965\
        );

    \I__2549\ : LocalMux
    port map (
            O => \N__22027\,
            I => \N__21962\
        );

    \I__2548\ : InMux
    port map (
            O => \N__22026\,
            I => \N__21959\
        );

    \I__2547\ : InMux
    port map (
            O => \N__22025\,
            I => \N__21956\
        );

    \I__2546\ : LocalMux
    port map (
            O => \N__22018\,
            I => \N__21953\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__22015\,
            I => \N__21944\
        );

    \I__2544\ : LocalMux
    port map (
            O => \N__22008\,
            I => \N__21944\
        );

    \I__2543\ : Span4Mux_v
    port map (
            O => \N__21999\,
            I => \N__21944\
        );

    \I__2542\ : Span4Mux_v
    port map (
            O => \N__21992\,
            I => \N__21944\
        );

    \I__2541\ : InMux
    port map (
            O => \N__21991\,
            I => \N__21937\
        );

    \I__2540\ : InMux
    port map (
            O => \N__21990\,
            I => \N__21937\
        );

    \I__2539\ : InMux
    port map (
            O => \N__21989\,
            I => \N__21937\
        );

    \I__2538\ : Span4Mux_h
    port map (
            O => \N__21984\,
            I => \N__21934\
        );

    \I__2537\ : InMux
    port map (
            O => \N__21983\,
            I => \N__21931\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__21968\,
            I => adc_state_2_adj_1474
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__21965\,
            I => adc_state_2_adj_1474
        );

    \I__2534\ : Odrv4
    port map (
            O => \N__21962\,
            I => adc_state_2_adj_1474
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__21959\,
            I => adc_state_2_adj_1474
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__21956\,
            I => adc_state_2_adj_1474
        );

    \I__2531\ : Odrv4
    port map (
            O => \N__21953\,
            I => adc_state_2_adj_1474
        );

    \I__2530\ : Odrv4
    port map (
            O => \N__21944\,
            I => adc_state_2_adj_1474
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__21937\,
            I => adc_state_2_adj_1474
        );

    \I__2528\ : Odrv4
    port map (
            O => \N__21934\,
            I => adc_state_2_adj_1474
        );

    \I__2527\ : LocalMux
    port map (
            O => \N__21931\,
            I => adc_state_2_adj_1474
        );

    \I__2526\ : CascadeMux
    port map (
            O => \N__21910\,
            I => \N__21907\
        );

    \I__2525\ : InMux
    port map (
            O => \N__21907\,
            I => \N__21904\
        );

    \I__2524\ : LocalMux
    port map (
            O => \N__21904\,
            I => \N__21900\
        );

    \I__2523\ : InMux
    port map (
            O => \N__21903\,
            I => \N__21897\
        );

    \I__2522\ : Span12Mux_v
    port map (
            O => \N__21900\,
            I => \N__21892\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__21897\,
            I => \N__21892\
        );

    \I__2520\ : Odrv12
    port map (
            O => \N__21892\,
            I => \RTD.n20487\
        );

    \I__2519\ : InMux
    port map (
            O => \N__21889\,
            I => \N__21886\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__21886\,
            I => \N__21883\
        );

    \I__2517\ : Span4Mux_h
    port map (
            O => \N__21883\,
            I => \N__21880\
        );

    \I__2516\ : Span4Mux_v
    port map (
            O => \N__21880\,
            I => \N__21877\
        );

    \I__2515\ : Odrv4
    port map (
            O => \N__21877\,
            I => buf_data_iac_22
        );

    \I__2514\ : IoInMux
    port map (
            O => \N__21874\,
            I => \N__21871\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__21871\,
            I => \N__21868\
        );

    \I__2512\ : Span12Mux_s6_v
    port map (
            O => \N__21868\,
            I => \N__21864\
        );

    \I__2511\ : InMux
    port map (
            O => \N__21867\,
            I => \N__21861\
        );

    \I__2510\ : Odrv12
    port map (
            O => \N__21864\,
            I => \DDS_MOSI1\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__21861\,
            I => \DDS_MOSI1\
        );

    \I__2508\ : InMux
    port map (
            O => \N__21856\,
            I => \N__21853\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__21853\,
            I => \N__21849\
        );

    \I__2506\ : InMux
    port map (
            O => \N__21852\,
            I => \N__21846\
        );

    \I__2505\ : Span4Mux_v
    port map (
            O => \N__21849\,
            I => \N__21843\
        );

    \I__2504\ : LocalMux
    port map (
            O => \N__21846\,
            I => \N__21840\
        );

    \I__2503\ : Span4Mux_v
    port map (
            O => \N__21843\,
            I => \N__21834\
        );

    \I__2502\ : Span4Mux_h
    port map (
            O => \N__21840\,
            I => \N__21834\
        );

    \I__2501\ : InMux
    port map (
            O => \N__21839\,
            I => \N__21831\
        );

    \I__2500\ : Sp12to4
    port map (
            O => \N__21834\,
            I => \N__21828\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__21831\,
            I => buf_adcdata_vac_21
        );

    \I__2498\ : Odrv12
    port map (
            O => \N__21828\,
            I => buf_adcdata_vac_21
        );

    \I__2497\ : CascadeMux
    port map (
            O => \N__21823\,
            I => \N__21820\
        );

    \I__2496\ : InMux
    port map (
            O => \N__21820\,
            I => \N__21817\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__21817\,
            I => \N__21814\
        );

    \I__2494\ : Span4Mux_h
    port map (
            O => \N__21814\,
            I => \N__21810\
        );

    \I__2493\ : InMux
    port map (
            O => \N__21813\,
            I => \N__21807\
        );

    \I__2492\ : Odrv4
    port map (
            O => \N__21810\,
            I => \buf_readRTD_8\
        );

    \I__2491\ : LocalMux
    port map (
            O => \N__21807\,
            I => \buf_readRTD_8\
        );

    \I__2490\ : CascadeMux
    port map (
            O => \N__21802\,
            I => \N__21798\
        );

    \I__2489\ : CascadeMux
    port map (
            O => \N__21801\,
            I => \N__21795\
        );

    \I__2488\ : InMux
    port map (
            O => \N__21798\,
            I => \N__21791\
        );

    \I__2487\ : InMux
    port map (
            O => \N__21795\,
            I => \N__21786\
        );

    \I__2486\ : InMux
    port map (
            O => \N__21794\,
            I => \N__21786\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__21791\,
            I => cmd_rdadctmp_20
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__21786\,
            I => cmd_rdadctmp_20
        );

    \I__2483\ : CascadeMux
    port map (
            O => \N__21781\,
            I => \N__21778\
        );

    \I__2482\ : InMux
    port map (
            O => \N__21778\,
            I => \N__21773\
        );

    \I__2481\ : InMux
    port map (
            O => \N__21777\,
            I => \N__21770\
        );

    \I__2480\ : InMux
    port map (
            O => \N__21776\,
            I => \N__21767\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__21773\,
            I => cmd_rdadctmp_21
        );

    \I__2478\ : LocalMux
    port map (
            O => \N__21770\,
            I => cmd_rdadctmp_21
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__21767\,
            I => cmd_rdadctmp_21
        );

    \I__2476\ : CascadeMux
    port map (
            O => \N__21760\,
            I => \N__21756\
        );

    \I__2475\ : CascadeMux
    port map (
            O => \N__21759\,
            I => \N__21753\
        );

    \I__2474\ : InMux
    port map (
            O => \N__21756\,
            I => \N__21749\
        );

    \I__2473\ : InMux
    port map (
            O => \N__21753\,
            I => \N__21746\
        );

    \I__2472\ : InMux
    port map (
            O => \N__21752\,
            I => \N__21743\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__21749\,
            I => cmd_rdadctmp_19
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__21746\,
            I => cmd_rdadctmp_19
        );

    \I__2469\ : LocalMux
    port map (
            O => \N__21743\,
            I => cmd_rdadctmp_19
        );

    \I__2468\ : CascadeMux
    port map (
            O => \N__21736\,
            I => \N__21733\
        );

    \I__2467\ : InMux
    port map (
            O => \N__21733\,
            I => \N__21729\
        );

    \I__2466\ : CascadeMux
    port map (
            O => \N__21732\,
            I => \N__21726\
        );

    \I__2465\ : LocalMux
    port map (
            O => \N__21729\,
            I => \N__21722\
        );

    \I__2464\ : InMux
    port map (
            O => \N__21726\,
            I => \N__21719\
        );

    \I__2463\ : InMux
    port map (
            O => \N__21725\,
            I => \N__21716\
        );

    \I__2462\ : Odrv4
    port map (
            O => \N__21722\,
            I => cmd_rdadctmp_18
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__21719\,
            I => cmd_rdadctmp_18
        );

    \I__2460\ : LocalMux
    port map (
            O => \N__21716\,
            I => cmd_rdadctmp_18
        );

    \I__2459\ : InMux
    port map (
            O => \N__21709\,
            I => \N__21706\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__21706\,
            I => \N__21703\
        );

    \I__2457\ : Odrv4
    port map (
            O => \N__21703\,
            I => buf_data_iac_11
        );

    \I__2456\ : CascadeMux
    port map (
            O => \N__21700\,
            I => \N__21697\
        );

    \I__2455\ : InMux
    port map (
            O => \N__21697\,
            I => \N__21692\
        );

    \I__2454\ : InMux
    port map (
            O => \N__21696\,
            I => \N__21687\
        );

    \I__2453\ : InMux
    port map (
            O => \N__21695\,
            I => \N__21687\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__21692\,
            I => \N__21684\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__21687\,
            I => \N__21681\
        );

    \I__2450\ : Odrv4
    port map (
            O => \N__21684\,
            I => cmd_rdadctmp_17
        );

    \I__2449\ : Odrv4
    port map (
            O => \N__21681\,
            I => cmd_rdadctmp_17
        );

    \I__2448\ : InMux
    port map (
            O => \N__21676\,
            I => \N__21673\
        );

    \I__2447\ : LocalMux
    port map (
            O => \N__21673\,
            I => \N__21668\
        );

    \I__2446\ : InMux
    port map (
            O => \N__21672\,
            I => \N__21665\
        );

    \I__2445\ : InMux
    port map (
            O => \N__21671\,
            I => \N__21662\
        );

    \I__2444\ : Span4Mux_h
    port map (
            O => \N__21668\,
            I => \N__21659\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__21665\,
            I => \N__21656\
        );

    \I__2442\ : LocalMux
    port map (
            O => \N__21662\,
            I => buf_adcdata_iac_9
        );

    \I__2441\ : Odrv4
    port map (
            O => \N__21659\,
            I => buf_adcdata_iac_9
        );

    \I__2440\ : Odrv12
    port map (
            O => \N__21656\,
            I => buf_adcdata_iac_9
        );

    \I__2439\ : IoInMux
    port map (
            O => \N__21649\,
            I => \N__21646\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__21646\,
            I => \N__21643\
        );

    \I__2437\ : Span4Mux_s2_v
    port map (
            O => \N__21643\,
            I => \N__21640\
        );

    \I__2436\ : Span4Mux_v
    port map (
            O => \N__21640\,
            I => \N__21637\
        );

    \I__2435\ : Span4Mux_h
    port map (
            O => \N__21637\,
            I => \N__21634\
        );

    \I__2434\ : Odrv4
    port map (
            O => \N__21634\,
            I => \DDS_MCLK1\
        );

    \I__2433\ : IoInMux
    port map (
            O => \N__21631\,
            I => \N__21628\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__21628\,
            I => \N__21625\
        );

    \I__2431\ : Span4Mux_s3_v
    port map (
            O => \N__21625\,
            I => \N__21622\
        );

    \I__2430\ : Span4Mux_v
    port map (
            O => \N__21622\,
            I => \N__21619\
        );

    \I__2429\ : Span4Mux_h
    port map (
            O => \N__21619\,
            I => \N__21616\
        );

    \I__2428\ : Odrv4
    port map (
            O => \N__21616\,
            I => \DDS_CS1\
        );

    \I__2427\ : IoInMux
    port map (
            O => \N__21613\,
            I => \N__21610\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__21610\,
            I => \N__21607\
        );

    \I__2425\ : IoSpan4Mux
    port map (
            O => \N__21607\,
            I => \N__21604\
        );

    \I__2424\ : Span4Mux_s2_v
    port map (
            O => \N__21604\,
            I => \N__21600\
        );

    \I__2423\ : CascadeMux
    port map (
            O => \N__21603\,
            I => \N__21597\
        );

    \I__2422\ : Sp12to4
    port map (
            O => \N__21600\,
            I => \N__21594\
        );

    \I__2421\ : InMux
    port map (
            O => \N__21597\,
            I => \N__21591\
        );

    \I__2420\ : Odrv12
    port map (
            O => \N__21594\,
            I => \DDS_SCK1\
        );

    \I__2419\ : LocalMux
    port map (
            O => \N__21591\,
            I => \DDS_SCK1\
        );

    \I__2418\ : CascadeMux
    port map (
            O => \N__21586\,
            I => \n23_adj_1512_cascade_\
        );

    \I__2417\ : CascadeMux
    port map (
            O => \N__21583\,
            I => \N__21580\
        );

    \I__2416\ : InMux
    port map (
            O => \N__21580\,
            I => \N__21576\
        );

    \I__2415\ : InMux
    port map (
            O => \N__21579\,
            I => \N__21573\
        );

    \I__2414\ : LocalMux
    port map (
            O => \N__21576\,
            I => cmd_rdadctmp_6_adj_1437
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__21573\,
            I => cmd_rdadctmp_6_adj_1437
        );

    \I__2412\ : CascadeMux
    port map (
            O => \N__21568\,
            I => \N__21564\
        );

    \I__2411\ : InMux
    port map (
            O => \N__21567\,
            I => \N__21561\
        );

    \I__2410\ : InMux
    port map (
            O => \N__21564\,
            I => \N__21558\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__21561\,
            I => \N__21554\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__21558\,
            I => \N__21551\
        );

    \I__2407\ : InMux
    port map (
            O => \N__21557\,
            I => \N__21548\
        );

    \I__2406\ : Odrv12
    port map (
            O => \N__21554\,
            I => cmd_rdadctmp_21_adj_1422
        );

    \I__2405\ : Odrv4
    port map (
            O => \N__21551\,
            I => cmd_rdadctmp_21_adj_1422
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__21548\,
            I => cmd_rdadctmp_21_adj_1422
        );

    \I__2403\ : CascadeMux
    port map (
            O => \N__21541\,
            I => \N__21537\
        );

    \I__2402\ : InMux
    port map (
            O => \N__21540\,
            I => \N__21534\
        );

    \I__2401\ : InMux
    port map (
            O => \N__21537\,
            I => \N__21530\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__21534\,
            I => \N__21527\
        );

    \I__2399\ : InMux
    port map (
            O => \N__21533\,
            I => \N__21524\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__21530\,
            I => buf_adcdata_vac_13
        );

    \I__2397\ : Odrv4
    port map (
            O => \N__21527\,
            I => buf_adcdata_vac_13
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__21524\,
            I => buf_adcdata_vac_13
        );

    \I__2395\ : CascadeMux
    port map (
            O => \N__21517\,
            I => \N__21514\
        );

    \I__2394\ : InMux
    port map (
            O => \N__21514\,
            I => \N__21510\
        );

    \I__2393\ : InMux
    port map (
            O => \N__21513\,
            I => \N__21507\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__21510\,
            I => cmd_rdadctmp_4_adj_1439
        );

    \I__2391\ : LocalMux
    port map (
            O => \N__21507\,
            I => cmd_rdadctmp_4_adj_1439
        );

    \I__2390\ : InMux
    port map (
            O => \N__21502\,
            I => \N__21496\
        );

    \I__2389\ : InMux
    port map (
            O => \N__21501\,
            I => \N__21496\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__21496\,
            I => cmd_rdadctmp_5_adj_1438
        );

    \I__2387\ : InMux
    port map (
            O => \N__21493\,
            I => \N__21490\
        );

    \I__2386\ : LocalMux
    port map (
            O => \N__21490\,
            I => \N__21487\
        );

    \I__2385\ : Span4Mux_h
    port map (
            O => \N__21487\,
            I => \N__21484\
        );

    \I__2384\ : Odrv4
    port map (
            O => \N__21484\,
            I => buf_data_iac_14
        );

    \I__2383\ : InMux
    port map (
            O => \N__21481\,
            I => \N__21478\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__21478\,
            I => \N__21475\
        );

    \I__2381\ : Span4Mux_h
    port map (
            O => \N__21475\,
            I => \N__21470\
        );

    \I__2380\ : InMux
    port map (
            O => \N__21474\,
            I => \N__21467\
        );

    \I__2379\ : InMux
    port map (
            O => \N__21473\,
            I => \N__21464\
        );

    \I__2378\ : Span4Mux_v
    port map (
            O => \N__21470\,
            I => \N__21461\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__21467\,
            I => \N__21458\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__21464\,
            I => buf_adcdata_vac_3
        );

    \I__2375\ : Odrv4
    port map (
            O => \N__21461\,
            I => buf_adcdata_vac_3
        );

    \I__2374\ : Odrv4
    port map (
            O => \N__21458\,
            I => buf_adcdata_vac_3
        );

    \I__2373\ : CascadeMux
    port map (
            O => \N__21451\,
            I => \N__21448\
        );

    \I__2372\ : InMux
    port map (
            O => \N__21448\,
            I => \N__21443\
        );

    \I__2371\ : CascadeMux
    port map (
            O => \N__21447\,
            I => \N__21440\
        );

    \I__2370\ : CascadeMux
    port map (
            O => \N__21446\,
            I => \N__21437\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__21443\,
            I => \N__21434\
        );

    \I__2368\ : InMux
    port map (
            O => \N__21440\,
            I => \N__21431\
        );

    \I__2367\ : InMux
    port map (
            O => \N__21437\,
            I => \N__21428\
        );

    \I__2366\ : Odrv4
    port map (
            O => \N__21434\,
            I => cmd_rdadctmp_8
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__21431\,
            I => cmd_rdadctmp_8
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__21428\,
            I => cmd_rdadctmp_8
        );

    \I__2363\ : CascadeMux
    port map (
            O => \N__21421\,
            I => \N__21417\
        );

    \I__2362\ : CascadeMux
    port map (
            O => \N__21420\,
            I => \N__21414\
        );

    \I__2361\ : InMux
    port map (
            O => \N__21417\,
            I => \N__21406\
        );

    \I__2360\ : InMux
    port map (
            O => \N__21414\,
            I => \N__21406\
        );

    \I__2359\ : InMux
    port map (
            O => \N__21413\,
            I => \N__21406\
        );

    \I__2358\ : LocalMux
    port map (
            O => \N__21406\,
            I => cmd_rdadctmp_22_adj_1421
        );

    \I__2357\ : InMux
    port map (
            O => \N__21403\,
            I => \N__21400\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__21400\,
            I => n19_adj_1487
        );

    \I__2355\ : InMux
    port map (
            O => \N__21397\,
            I => \N__21394\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__21394\,
            I => \N__21391\
        );

    \I__2353\ : Span4Mux_h
    port map (
            O => \N__21391\,
            I => \N__21388\
        );

    \I__2352\ : Span4Mux_v
    port map (
            O => \N__21388\,
            I => \N__21383\
        );

    \I__2351\ : InMux
    port map (
            O => \N__21387\,
            I => \N__21378\
        );

    \I__2350\ : InMux
    port map (
            O => \N__21386\,
            I => \N__21378\
        );

    \I__2349\ : Odrv4
    port map (
            O => \N__21383\,
            I => buf_adcdata_vac_8
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__21378\,
            I => buf_adcdata_vac_8
        );

    \I__2347\ : InMux
    port map (
            O => \N__21373\,
            I => \N__21370\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__21370\,
            I => \N__21367\
        );

    \I__2345\ : Span4Mux_v
    port map (
            O => \N__21367\,
            I => \N__21363\
        );

    \I__2344\ : CascadeMux
    port map (
            O => \N__21366\,
            I => \N__21360\
        );

    \I__2343\ : Span4Mux_h
    port map (
            O => \N__21363\,
            I => \N__21357\
        );

    \I__2342\ : InMux
    port map (
            O => \N__21360\,
            I => \N__21354\
        );

    \I__2341\ : Odrv4
    port map (
            O => \N__21357\,
            I => \buf_readRTD_0\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__21354\,
            I => \buf_readRTD_0\
        );

    \I__2339\ : CascadeMux
    port map (
            O => \N__21349\,
            I => \n19_adj_1479_cascade_\
        );

    \I__2338\ : CascadeMux
    port map (
            O => \N__21346\,
            I => \N__21342\
        );

    \I__2337\ : CascadeMux
    port map (
            O => \N__21345\,
            I => \N__21339\
        );

    \I__2336\ : InMux
    port map (
            O => \N__21342\,
            I => \N__21335\
        );

    \I__2335\ : InMux
    port map (
            O => \N__21339\,
            I => \N__21332\
        );

    \I__2334\ : InMux
    port map (
            O => \N__21338\,
            I => \N__21329\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__21335\,
            I => cmd_rdadctmp_29_adj_1414
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__21332\,
            I => cmd_rdadctmp_29_adj_1414
        );

    \I__2331\ : LocalMux
    port map (
            O => \N__21329\,
            I => cmd_rdadctmp_29_adj_1414
        );

    \I__2330\ : CascadeMux
    port map (
            O => \N__21322\,
            I => \N__21318\
        );

    \I__2329\ : CascadeMux
    port map (
            O => \N__21321\,
            I => \N__21315\
        );

    \I__2328\ : InMux
    port map (
            O => \N__21318\,
            I => \N__21311\
        );

    \I__2327\ : InMux
    port map (
            O => \N__21315\,
            I => \N__21308\
        );

    \I__2326\ : InMux
    port map (
            O => \N__21314\,
            I => \N__21305\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__21311\,
            I => cmd_rdadctmp_10
        );

    \I__2324\ : LocalMux
    port map (
            O => \N__21308\,
            I => cmd_rdadctmp_10
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__21305\,
            I => cmd_rdadctmp_10
        );

    \I__2322\ : CascadeMux
    port map (
            O => \N__21298\,
            I => \N__21294\
        );

    \I__2321\ : CascadeMux
    port map (
            O => \N__21297\,
            I => \N__21291\
        );

    \I__2320\ : InMux
    port map (
            O => \N__21294\,
            I => \N__21287\
        );

    \I__2319\ : InMux
    port map (
            O => \N__21291\,
            I => \N__21282\
        );

    \I__2318\ : InMux
    port map (
            O => \N__21290\,
            I => \N__21282\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__21287\,
            I => cmd_rdadctmp_26_adj_1417
        );

    \I__2316\ : LocalMux
    port map (
            O => \N__21282\,
            I => cmd_rdadctmp_26_adj_1417
        );

    \I__2315\ : CascadeMux
    port map (
            O => \N__21277\,
            I => \N__21273\
        );

    \I__2314\ : CascadeMux
    port map (
            O => \N__21276\,
            I => \N__21270\
        );

    \I__2313\ : InMux
    port map (
            O => \N__21273\,
            I => \N__21266\
        );

    \I__2312\ : InMux
    port map (
            O => \N__21270\,
            I => \N__21263\
        );

    \I__2311\ : InMux
    port map (
            O => \N__21269\,
            I => \N__21260\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__21266\,
            I => cmd_rdadctmp_27_adj_1416
        );

    \I__2309\ : LocalMux
    port map (
            O => \N__21263\,
            I => cmd_rdadctmp_27_adj_1416
        );

    \I__2308\ : LocalMux
    port map (
            O => \N__21260\,
            I => cmd_rdadctmp_27_adj_1416
        );

    \I__2307\ : InMux
    port map (
            O => \N__21253\,
            I => \N__21246\
        );

    \I__2306\ : InMux
    port map (
            O => \N__21252\,
            I => \N__21246\
        );

    \I__2305\ : InMux
    port map (
            O => \N__21251\,
            I => \N__21243\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__21246\,
            I => cmd_rdadctmp_9
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__21243\,
            I => cmd_rdadctmp_9
        );

    \I__2302\ : InMux
    port map (
            O => \N__21238\,
            I => \N__21234\
        );

    \I__2301\ : CascadeMux
    port map (
            O => \N__21237\,
            I => \N__21231\
        );

    \I__2300\ : LocalMux
    port map (
            O => \N__21234\,
            I => \N__21227\
        );

    \I__2299\ : InMux
    port map (
            O => \N__21231\,
            I => \N__21224\
        );

    \I__2298\ : InMux
    port map (
            O => \N__21230\,
            I => \N__21221\
        );

    \I__2297\ : Odrv4
    port map (
            O => \N__21227\,
            I => cmd_rdadctmp_23_adj_1420
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__21224\,
            I => cmd_rdadctmp_23_adj_1420
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__21221\,
            I => cmd_rdadctmp_23_adj_1420
        );

    \I__2294\ : InMux
    port map (
            O => \N__21214\,
            I => \N__21210\
        );

    \I__2293\ : InMux
    port map (
            O => \N__21213\,
            I => \N__21207\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__21210\,
            I => \RTD.cfg_buf_5\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__21207\,
            I => \RTD.cfg_buf_5\
        );

    \I__2290\ : InMux
    port map (
            O => \N__21202\,
            I => \N__21199\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__21199\,
            I => \RTD.n11_adj_1396\
        );

    \I__2288\ : InMux
    port map (
            O => \N__21196\,
            I => \N__21190\
        );

    \I__2287\ : InMux
    port map (
            O => \N__21195\,
            I => \N__21190\
        );

    \I__2286\ : LocalMux
    port map (
            O => \N__21190\,
            I => \RTD.cfg_buf_3\
        );

    \I__2285\ : InMux
    port map (
            O => \N__21187\,
            I => \N__21170\
        );

    \I__2284\ : InMux
    port map (
            O => \N__21186\,
            I => \N__21170\
        );

    \I__2283\ : InMux
    port map (
            O => \N__21185\,
            I => \N__21170\
        );

    \I__2282\ : InMux
    port map (
            O => \N__21184\,
            I => \N__21170\
        );

    \I__2281\ : InMux
    port map (
            O => \N__21183\,
            I => \N__21170\
        );

    \I__2280\ : InMux
    port map (
            O => \N__21182\,
            I => \N__21165\
        );

    \I__2279\ : InMux
    port map (
            O => \N__21181\,
            I => \N__21165\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__21170\,
            I => n18586
        );

    \I__2277\ : LocalMux
    port map (
            O => \N__21165\,
            I => n18586
        );

    \I__2276\ : InMux
    port map (
            O => \N__21160\,
            I => \N__21149\
        );

    \I__2275\ : InMux
    port map (
            O => \N__21159\,
            I => \N__21146\
        );

    \I__2274\ : InMux
    port map (
            O => \N__21158\,
            I => \N__21141\
        );

    \I__2273\ : InMux
    port map (
            O => \N__21157\,
            I => \N__21141\
        );

    \I__2272\ : InMux
    port map (
            O => \N__21156\,
            I => \N__21134\
        );

    \I__2271\ : InMux
    port map (
            O => \N__21155\,
            I => \N__21134\
        );

    \I__2270\ : InMux
    port map (
            O => \N__21154\,
            I => \N__21134\
        );

    \I__2269\ : InMux
    port map (
            O => \N__21153\,
            I => \N__21131\
        );

    \I__2268\ : InMux
    port map (
            O => \N__21152\,
            I => \N__21128\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__21149\,
            I => n13162
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__21146\,
            I => n13162
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__21141\,
            I => n13162
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__21134\,
            I => n13162
        );

    \I__2263\ : LocalMux
    port map (
            O => \N__21131\,
            I => n13162
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__21128\,
            I => n13162
        );

    \I__2261\ : InMux
    port map (
            O => \N__21115\,
            I => \N__21111\
        );

    \I__2260\ : InMux
    port map (
            O => \N__21114\,
            I => \N__21108\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__21111\,
            I => \RTD.cfg_buf_6\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__21108\,
            I => \RTD.cfg_buf_6\
        );

    \I__2257\ : CascadeMux
    port map (
            O => \N__21103\,
            I => \N__21100\
        );

    \I__2256\ : InMux
    port map (
            O => \N__21100\,
            I => \N__21097\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__21097\,
            I => \N__21093\
        );

    \I__2254\ : CascadeMux
    port map (
            O => \N__21096\,
            I => \N__21090\
        );

    \I__2253\ : Span4Mux_h
    port map (
            O => \N__21093\,
            I => \N__21087\
        );

    \I__2252\ : InMux
    port map (
            O => \N__21090\,
            I => \N__21084\
        );

    \I__2251\ : Odrv4
    port map (
            O => \N__21087\,
            I => \buf_readRTD_11\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__21084\,
            I => \buf_readRTD_11\
        );

    \I__2249\ : CascadeMux
    port map (
            O => \N__21079\,
            I => \n22099_cascade_\
        );

    \I__2248\ : CascadeMux
    port map (
            O => \N__21076\,
            I => \n22102_cascade_\
        );

    \I__2247\ : InMux
    port map (
            O => \N__21073\,
            I => \N__21070\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__21070\,
            I => \N__21066\
        );

    \I__2245\ : InMux
    port map (
            O => \N__21069\,
            I => \N__21062\
        );

    \I__2244\ : Span4Mux_h
    port map (
            O => \N__21066\,
            I => \N__21059\
        );

    \I__2243\ : InMux
    port map (
            O => \N__21065\,
            I => \N__21056\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__21062\,
            I => buf_adcdata_vac_19
        );

    \I__2241\ : Odrv4
    port map (
            O => \N__21059\,
            I => buf_adcdata_vac_19
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__21056\,
            I => buf_adcdata_vac_19
        );

    \I__2239\ : CascadeMux
    port map (
            O => \N__21049\,
            I => \n19_adj_1610_cascade_\
        );

    \I__2238\ : InMux
    port map (
            O => \N__21046\,
            I => \N__21043\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__21043\,
            I => \N__21039\
        );

    \I__2236\ : InMux
    port map (
            O => \N__21042\,
            I => \N__21035\
        );

    \I__2235\ : Span4Mux_v
    port map (
            O => \N__21039\,
            I => \N__21032\
        );

    \I__2234\ : InMux
    port map (
            O => \N__21038\,
            I => \N__21029\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__21035\,
            I => buf_adcdata_iac_3
        );

    \I__2232\ : Odrv4
    port map (
            O => \N__21032\,
            I => buf_adcdata_iac_3
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__21029\,
            I => buf_adcdata_iac_3
        );

    \I__2230\ : InMux
    port map (
            O => \N__21022\,
            I => \N__21019\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__21019\,
            I => n22_adj_1611
        );

    \I__2228\ : InMux
    port map (
            O => \N__21016\,
            I => \N__21013\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__21013\,
            I => \RTD.cfg_tmp_5\
        );

    \I__2226\ : InMux
    port map (
            O => \N__21010\,
            I => \N__21007\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__21007\,
            I => \RTD.cfg_tmp_6\
        );

    \I__2224\ : CascadeMux
    port map (
            O => \N__21004\,
            I => \N__21001\
        );

    \I__2223\ : InMux
    port map (
            O => \N__21001\,
            I => \N__20998\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__20998\,
            I => \N__20995\
        );

    \I__2221\ : Span4Mux_h
    port map (
            O => \N__20995\,
            I => \N__20991\
        );

    \I__2220\ : InMux
    port map (
            O => \N__20994\,
            I => \N__20988\
        );

    \I__2219\ : Odrv4
    port map (
            O => \N__20991\,
            I => \RTD.cfg_tmp_7\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__20988\,
            I => \RTD.cfg_tmp_7\
        );

    \I__2217\ : InMux
    port map (
            O => \N__20983\,
            I => \N__20980\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__20980\,
            I => \RTD.cfg_tmp_0\
        );

    \I__2215\ : CascadeMux
    port map (
            O => \N__20977\,
            I => \N__20974\
        );

    \I__2214\ : InMux
    port map (
            O => \N__20974\,
            I => \N__20971\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__20971\,
            I => \N__20960\
        );

    \I__2212\ : InMux
    port map (
            O => \N__20970\,
            I => \N__20949\
        );

    \I__2211\ : InMux
    port map (
            O => \N__20969\,
            I => \N__20949\
        );

    \I__2210\ : InMux
    port map (
            O => \N__20968\,
            I => \N__20949\
        );

    \I__2209\ : InMux
    port map (
            O => \N__20967\,
            I => \N__20949\
        );

    \I__2208\ : InMux
    port map (
            O => \N__20966\,
            I => \N__20949\
        );

    \I__2207\ : InMux
    port map (
            O => \N__20965\,
            I => \N__20946\
        );

    \I__2206\ : InMux
    port map (
            O => \N__20964\,
            I => \N__20929\
        );

    \I__2205\ : InMux
    port map (
            O => \N__20963\,
            I => \N__20920\
        );

    \I__2204\ : Span4Mux_v
    port map (
            O => \N__20960\,
            I => \N__20915\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__20949\,
            I => \N__20915\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__20946\,
            I => \N__20910\
        );

    \I__2201\ : InMux
    port map (
            O => \N__20945\,
            I => \N__20907\
        );

    \I__2200\ : InMux
    port map (
            O => \N__20944\,
            I => \N__20898\
        );

    \I__2199\ : InMux
    port map (
            O => \N__20943\,
            I => \N__20898\
        );

    \I__2198\ : InMux
    port map (
            O => \N__20942\,
            I => \N__20898\
        );

    \I__2197\ : InMux
    port map (
            O => \N__20941\,
            I => \N__20898\
        );

    \I__2196\ : InMux
    port map (
            O => \N__20940\,
            I => \N__20890\
        );

    \I__2195\ : InMux
    port map (
            O => \N__20939\,
            I => \N__20873\
        );

    \I__2194\ : InMux
    port map (
            O => \N__20938\,
            I => \N__20873\
        );

    \I__2193\ : InMux
    port map (
            O => \N__20937\,
            I => \N__20873\
        );

    \I__2192\ : InMux
    port map (
            O => \N__20936\,
            I => \N__20873\
        );

    \I__2191\ : InMux
    port map (
            O => \N__20935\,
            I => \N__20873\
        );

    \I__2190\ : InMux
    port map (
            O => \N__20934\,
            I => \N__20873\
        );

    \I__2189\ : InMux
    port map (
            O => \N__20933\,
            I => \N__20873\
        );

    \I__2188\ : InMux
    port map (
            O => \N__20932\,
            I => \N__20873\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__20929\,
            I => \N__20870\
        );

    \I__2186\ : InMux
    port map (
            O => \N__20928\,
            I => \N__20867\
        );

    \I__2185\ : InMux
    port map (
            O => \N__20927\,
            I => \N__20856\
        );

    \I__2184\ : InMux
    port map (
            O => \N__20926\,
            I => \N__20856\
        );

    \I__2183\ : InMux
    port map (
            O => \N__20925\,
            I => \N__20856\
        );

    \I__2182\ : InMux
    port map (
            O => \N__20924\,
            I => \N__20856\
        );

    \I__2181\ : InMux
    port map (
            O => \N__20923\,
            I => \N__20856\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__20920\,
            I => \N__20851\
        );

    \I__2179\ : Span4Mux_v
    port map (
            O => \N__20915\,
            I => \N__20851\
        );

    \I__2178\ : InMux
    port map (
            O => \N__20914\,
            I => \N__20846\
        );

    \I__2177\ : InMux
    port map (
            O => \N__20913\,
            I => \N__20846\
        );

    \I__2176\ : Span4Mux_h
    port map (
            O => \N__20910\,
            I => \N__20839\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__20907\,
            I => \N__20839\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__20898\,
            I => \N__20839\
        );

    \I__2173\ : InMux
    port map (
            O => \N__20897\,
            I => \N__20828\
        );

    \I__2172\ : InMux
    port map (
            O => \N__20896\,
            I => \N__20828\
        );

    \I__2171\ : InMux
    port map (
            O => \N__20895\,
            I => \N__20828\
        );

    \I__2170\ : InMux
    port map (
            O => \N__20894\,
            I => \N__20828\
        );

    \I__2169\ : InMux
    port map (
            O => \N__20893\,
            I => \N__20828\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__20890\,
            I => \RTD.adc_state_0\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__20873\,
            I => \RTD.adc_state_0\
        );

    \I__2166\ : Odrv12
    port map (
            O => \N__20870\,
            I => \RTD.adc_state_0\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__20867\,
            I => \RTD.adc_state_0\
        );

    \I__2164\ : LocalMux
    port map (
            O => \N__20856\,
            I => \RTD.adc_state_0\
        );

    \I__2163\ : Odrv4
    port map (
            O => \N__20851\,
            I => \RTD.adc_state_0\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__20846\,
            I => \RTD.adc_state_0\
        );

    \I__2161\ : Odrv4
    port map (
            O => \N__20839\,
            I => \RTD.adc_state_0\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__20828\,
            I => \RTD.adc_state_0\
        );

    \I__2159\ : CascadeMux
    port map (
            O => \N__20809\,
            I => \n18586_cascade_\
        );

    \I__2158\ : InMux
    port map (
            O => \N__20806\,
            I => \N__20800\
        );

    \I__2157\ : InMux
    port map (
            O => \N__20805\,
            I => \N__20800\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__20800\,
            I => cfg_buf_0
        );

    \I__2155\ : InMux
    port map (
            O => \N__20797\,
            I => \N__20794\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__20794\,
            I => \RTD.n9\
        );

    \I__2153\ : InMux
    port map (
            O => \N__20791\,
            I => \N__20787\
        );

    \I__2152\ : InMux
    port map (
            O => \N__20790\,
            I => \N__20784\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__20787\,
            I => \RTD.n11\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__20784\,
            I => \RTD.n11\
        );

    \I__2149\ : InMux
    port map (
            O => \N__20779\,
            I => \N__20776\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__20776\,
            I => \N__20773\
        );

    \I__2147\ : Odrv4
    port map (
            O => \N__20773\,
            I => \RTD.n14\
        );

    \I__2146\ : CascadeMux
    port map (
            O => \N__20770\,
            I => \RTD.n20722_cascade_\
        );

    \I__2145\ : CEMux
    port map (
            O => \N__20767\,
            I => \N__20764\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__20764\,
            I => \N__20761\
        );

    \I__2143\ : Span4Mux_h
    port map (
            O => \N__20761\,
            I => \N__20758\
        );

    \I__2142\ : Odrv4
    port map (
            O => \N__20758\,
            I => \RTD.n13198\
        );

    \I__2141\ : CascadeMux
    port map (
            O => \N__20755\,
            I => \RTD.n13198_cascade_\
        );

    \I__2140\ : SRMux
    port map (
            O => \N__20752\,
            I => \N__20749\
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__20749\,
            I => \N__20746\
        );

    \I__2138\ : Span4Mux_h
    port map (
            O => \N__20746\,
            I => \N__20743\
        );

    \I__2137\ : Odrv4
    port map (
            O => \N__20743\,
            I => \RTD.n14984\
        );

    \I__2136\ : SRMux
    port map (
            O => \N__20740\,
            I => \N__20737\
        );

    \I__2135\ : LocalMux
    port map (
            O => \N__20737\,
            I => \N__20734\
        );

    \I__2134\ : Odrv4
    port map (
            O => \N__20734\,
            I => \CLK_DDS.n16711\
        );

    \I__2133\ : InMux
    port map (
            O => \N__20731\,
            I => \N__20727\
        );

    \I__2132\ : InMux
    port map (
            O => \N__20730\,
            I => \N__20724\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__20727\,
            I => \RTD.n7285\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__20724\,
            I => \RTD.n7285\
        );

    \I__2129\ : CascadeMux
    port map (
            O => \N__20719\,
            I => \N__20716\
        );

    \I__2128\ : InMux
    port map (
            O => \N__20716\,
            I => \N__20713\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__20713\,
            I => \RTD.n11_adj_1394\
        );

    \I__2126\ : InMux
    port map (
            O => \N__20710\,
            I => \N__20707\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__20707\,
            I => \RTD.n21091\
        );

    \I__2124\ : CascadeMux
    port map (
            O => \N__20704\,
            I => \N__20701\
        );

    \I__2123\ : InMux
    port map (
            O => \N__20701\,
            I => \N__20698\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__20698\,
            I => \RTD.n33\
        );

    \I__2121\ : InMux
    port map (
            O => \N__20695\,
            I => \N__20692\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__20692\,
            I => \RTD.n17676\
        );

    \I__2119\ : InMux
    port map (
            O => \N__20689\,
            I => \N__20686\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__20686\,
            I => \RTD.n7_adj_1395\
        );

    \I__2117\ : CEMux
    port map (
            O => \N__20683\,
            I => \N__20680\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__20680\,
            I => \N__20676\
        );

    \I__2115\ : CEMux
    port map (
            O => \N__20679\,
            I => \N__20673\
        );

    \I__2114\ : Odrv12
    port map (
            O => \N__20676\,
            I => \RTD.n11712\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__20673\,
            I => \RTD.n11712\
        );

    \I__2112\ : CascadeMux
    port map (
            O => \N__20668\,
            I => \N__20665\
        );

    \I__2111\ : InMux
    port map (
            O => \N__20665\,
            I => \N__20662\
        );

    \I__2110\ : LocalMux
    port map (
            O => \N__20662\,
            I => \RTD.cfg_tmp_1\
        );

    \I__2109\ : InMux
    port map (
            O => \N__20659\,
            I => \N__20656\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__20656\,
            I => \RTD.cfg_tmp_2\
        );

    \I__2107\ : InMux
    port map (
            O => \N__20653\,
            I => \N__20650\
        );

    \I__2106\ : LocalMux
    port map (
            O => \N__20650\,
            I => \RTD.cfg_tmp_3\
        );

    \I__2105\ : InMux
    port map (
            O => \N__20647\,
            I => \N__20644\
        );

    \I__2104\ : LocalMux
    port map (
            O => \N__20644\,
            I => \RTD.cfg_tmp_4\
        );

    \I__2103\ : CEMux
    port map (
            O => \N__20641\,
            I => \N__20637\
        );

    \I__2102\ : CEMux
    port map (
            O => \N__20640\,
            I => \N__20634\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__20637\,
            I => \N__20631\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__20634\,
            I => \N__20628\
        );

    \I__2099\ : Span4Mux_h
    port map (
            O => \N__20631\,
            I => \N__20625\
        );

    \I__2098\ : Odrv12
    port map (
            O => \N__20628\,
            I => \CLK_DDS.n9\
        );

    \I__2097\ : Odrv4
    port map (
            O => \N__20625\,
            I => \CLK_DDS.n9\
        );

    \I__2096\ : InMux
    port map (
            O => \N__20620\,
            I => \N__20617\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__20617\,
            I => \N__20611\
        );

    \I__2094\ : InMux
    port map (
            O => \N__20616\,
            I => \N__20606\
        );

    \I__2093\ : InMux
    port map (
            O => \N__20615\,
            I => \N__20606\
        );

    \I__2092\ : InMux
    port map (
            O => \N__20614\,
            I => \N__20603\
        );

    \I__2091\ : Odrv4
    port map (
            O => \N__20611\,
            I => \RTD.bit_cnt_1\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__20606\,
            I => \RTD.bit_cnt_1\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__20603\,
            I => \RTD.bit_cnt_1\
        );

    \I__2088\ : InMux
    port map (
            O => \N__20596\,
            I => \N__20592\
        );

    \I__2087\ : CascadeMux
    port map (
            O => \N__20595\,
            I => \N__20589\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__20592\,
            I => \N__20583\
        );

    \I__2085\ : InMux
    port map (
            O => \N__20589\,
            I => \N__20576\
        );

    \I__2084\ : InMux
    port map (
            O => \N__20588\,
            I => \N__20576\
        );

    \I__2083\ : InMux
    port map (
            O => \N__20587\,
            I => \N__20576\
        );

    \I__2082\ : InMux
    port map (
            O => \N__20586\,
            I => \N__20573\
        );

    \I__2081\ : Odrv4
    port map (
            O => \N__20583\,
            I => \RTD.bit_cnt_0\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__20576\,
            I => \RTD.bit_cnt_0\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__20573\,
            I => \RTD.bit_cnt_0\
        );

    \I__2078\ : InMux
    port map (
            O => \N__20566\,
            I => \N__20563\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__20563\,
            I => \N__20558\
        );

    \I__2076\ : InMux
    port map (
            O => \N__20562\,
            I => \N__20555\
        );

    \I__2075\ : InMux
    port map (
            O => \N__20561\,
            I => \N__20552\
        );

    \I__2074\ : Odrv4
    port map (
            O => \N__20558\,
            I => \RTD.bit_cnt_2\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__20555\,
            I => \RTD.bit_cnt_2\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__20552\,
            I => \RTD.bit_cnt_2\
        );

    \I__2071\ : InMux
    port map (
            O => \N__20545\,
            I => \N__20541\
        );

    \I__2070\ : InMux
    port map (
            O => \N__20544\,
            I => \N__20537\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__20541\,
            I => \N__20534\
        );

    \I__2068\ : InMux
    port map (
            O => \N__20540\,
            I => \N__20531\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__20537\,
            I => \RTD.n17638\
        );

    \I__2066\ : Odrv4
    port map (
            O => \N__20534\,
            I => \RTD.n17638\
        );

    \I__2065\ : LocalMux
    port map (
            O => \N__20531\,
            I => \RTD.n17638\
        );

    \I__2064\ : CascadeMux
    port map (
            O => \N__20524\,
            I => \N__20521\
        );

    \I__2063\ : InMux
    port map (
            O => \N__20521\,
            I => \N__20514\
        );

    \I__2062\ : InMux
    port map (
            O => \N__20520\,
            I => \N__20511\
        );

    \I__2061\ : InMux
    port map (
            O => \N__20519\,
            I => \N__20508\
        );

    \I__2060\ : InMux
    port map (
            O => \N__20518\,
            I => \N__20505\
        );

    \I__2059\ : CascadeMux
    port map (
            O => \N__20517\,
            I => \N__20502\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__20514\,
            I => \N__20493\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__20511\,
            I => \N__20493\
        );

    \I__2056\ : LocalMux
    port map (
            O => \N__20508\,
            I => \N__20493\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__20505\,
            I => \N__20493\
        );

    \I__2054\ : InMux
    port map (
            O => \N__20502\,
            I => \N__20490\
        );

    \I__2053\ : Span4Mux_v
    port map (
            O => \N__20493\,
            I => \N__20487\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__20490\,
            I => \RTD.bit_cnt_3\
        );

    \I__2051\ : Odrv4
    port map (
            O => \N__20487\,
            I => \RTD.bit_cnt_3\
        );

    \I__2050\ : CascadeMux
    port map (
            O => \N__20482\,
            I => \RTD.n17638_cascade_\
        );

    \I__2049\ : InMux
    port map (
            O => \N__20479\,
            I => \N__20476\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__20476\,
            I => \N__20472\
        );

    \I__2047\ : InMux
    port map (
            O => \N__20475\,
            I => \N__20469\
        );

    \I__2046\ : Span4Mux_h
    port map (
            O => \N__20472\,
            I => \N__20466\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__20469\,
            I => \RTD.n1_adj_1392\
        );

    \I__2044\ : Odrv4
    port map (
            O => \N__20466\,
            I => \RTD.n1_adj_1392\
        );

    \I__2043\ : CascadeMux
    port map (
            O => \N__20461\,
            I => \RTD.n21063_cascade_\
        );

    \I__2042\ : CascadeMux
    port map (
            O => \N__20458\,
            I => \N__20454\
        );

    \I__2041\ : CascadeMux
    port map (
            O => \N__20457\,
            I => \N__20450\
        );

    \I__2040\ : InMux
    port map (
            O => \N__20454\,
            I => \N__20446\
        );

    \I__2039\ : InMux
    port map (
            O => \N__20453\,
            I => \N__20439\
        );

    \I__2038\ : InMux
    port map (
            O => \N__20450\,
            I => \N__20439\
        );

    \I__2037\ : InMux
    port map (
            O => \N__20449\,
            I => \N__20439\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__20446\,
            I => \N__20436\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__20439\,
            I => bit_cnt_1
        );

    \I__2034\ : Odrv4
    port map (
            O => \N__20436\,
            I => bit_cnt_1
        );

    \I__2033\ : InMux
    port map (
            O => \N__20431\,
            I => \N__20426\
        );

    \I__2032\ : InMux
    port map (
            O => \N__20430\,
            I => \N__20421\
        );

    \I__2031\ : InMux
    port map (
            O => \N__20429\,
            I => \N__20421\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__20426\,
            I => \N__20418\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__20421\,
            I => bit_cnt_2
        );

    \I__2028\ : Odrv4
    port map (
            O => \N__20418\,
            I => bit_cnt_2
        );

    \I__2027\ : InMux
    port map (
            O => \N__20413\,
            I => \N__20410\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__20410\,
            I => n8_adj_1409
        );

    \I__2025\ : InMux
    port map (
            O => \N__20407\,
            I => \N__20404\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__20404\,
            I => \N__20401\
        );

    \I__2023\ : Odrv4
    port map (
            O => \N__20401\,
            I => buf_data_iac_8
        );

    \I__2022\ : CascadeMux
    port map (
            O => \N__20398\,
            I => \N__20395\
        );

    \I__2021\ : CascadeBuf
    port map (
            O => \N__20395\,
            I => \N__20392\
        );

    \I__2020\ : CascadeMux
    port map (
            O => \N__20392\,
            I => \N__20389\
        );

    \I__2019\ : CascadeBuf
    port map (
            O => \N__20389\,
            I => \N__20386\
        );

    \I__2018\ : CascadeMux
    port map (
            O => \N__20386\,
            I => \N__20383\
        );

    \I__2017\ : CascadeBuf
    port map (
            O => \N__20383\,
            I => \N__20380\
        );

    \I__2016\ : CascadeMux
    port map (
            O => \N__20380\,
            I => \N__20377\
        );

    \I__2015\ : CascadeBuf
    port map (
            O => \N__20377\,
            I => \N__20374\
        );

    \I__2014\ : CascadeMux
    port map (
            O => \N__20374\,
            I => \N__20371\
        );

    \I__2013\ : CascadeBuf
    port map (
            O => \N__20371\,
            I => \N__20368\
        );

    \I__2012\ : CascadeMux
    port map (
            O => \N__20368\,
            I => \N__20364\
        );

    \I__2011\ : CascadeMux
    port map (
            O => \N__20367\,
            I => \N__20361\
        );

    \I__2010\ : CascadeBuf
    port map (
            O => \N__20364\,
            I => \N__20358\
        );

    \I__2009\ : CascadeBuf
    port map (
            O => \N__20361\,
            I => \N__20355\
        );

    \I__2008\ : CascadeMux
    port map (
            O => \N__20358\,
            I => \N__20352\
        );

    \I__2007\ : CascadeMux
    port map (
            O => \N__20355\,
            I => \N__20349\
        );

    \I__2006\ : CascadeBuf
    port map (
            O => \N__20352\,
            I => \N__20346\
        );

    \I__2005\ : InMux
    port map (
            O => \N__20349\,
            I => \N__20343\
        );

    \I__2004\ : CascadeMux
    port map (
            O => \N__20346\,
            I => \N__20340\
        );

    \I__2003\ : LocalMux
    port map (
            O => \N__20343\,
            I => \N__20337\
        );

    \I__2002\ : CascadeBuf
    port map (
            O => \N__20340\,
            I => \N__20334\
        );

    \I__2001\ : Span4Mux_v
    port map (
            O => \N__20337\,
            I => \N__20331\
        );

    \I__2000\ : CascadeMux
    port map (
            O => \N__20334\,
            I => \N__20328\
        );

    \I__1999\ : Span4Mux_v
    port map (
            O => \N__20331\,
            I => \N__20325\
        );

    \I__1998\ : CascadeBuf
    port map (
            O => \N__20328\,
            I => \N__20322\
        );

    \I__1997\ : Span4Mux_h
    port map (
            O => \N__20325\,
            I => \N__20319\
        );

    \I__1996\ : CascadeMux
    port map (
            O => \N__20322\,
            I => \N__20316\
        );

    \I__1995\ : Sp12to4
    port map (
            O => \N__20319\,
            I => \N__20313\
        );

    \I__1994\ : InMux
    port map (
            O => \N__20316\,
            I => \N__20310\
        );

    \I__1993\ : Odrv12
    port map (
            O => \N__20313\,
            I => \data_index_9_N_212_7\
        );

    \I__1992\ : LocalMux
    port map (
            O => \N__20310\,
            I => \data_index_9_N_212_7\
        );

    \I__1991\ : CascadeMux
    port map (
            O => \N__20305\,
            I => \N__20301\
        );

    \I__1990\ : InMux
    port map (
            O => \N__20304\,
            I => \N__20293\
        );

    \I__1989\ : InMux
    port map (
            O => \N__20301\,
            I => \N__20293\
        );

    \I__1988\ : InMux
    port map (
            O => \N__20300\,
            I => \N__20293\
        );

    \I__1987\ : LocalMux
    port map (
            O => \N__20293\,
            I => cmd_rdadctmp_28_adj_1415
        );

    \I__1986\ : CascadeMux
    port map (
            O => \N__20290\,
            I => \N__20287\
        );

    \I__1985\ : InMux
    port map (
            O => \N__20287\,
            I => \N__20284\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__20284\,
            I => \N__20281\
        );

    \I__1983\ : Span4Mux_v
    port map (
            O => \N__20281\,
            I => \N__20277\
        );

    \I__1982\ : CascadeMux
    port map (
            O => \N__20280\,
            I => \N__20274\
        );

    \I__1981\ : Span4Mux_v
    port map (
            O => \N__20277\,
            I => \N__20271\
        );

    \I__1980\ : InMux
    port map (
            O => \N__20274\,
            I => \N__20268\
        );

    \I__1979\ : Odrv4
    port map (
            O => \N__20271\,
            I => \buf_readRTD_5\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__20268\,
            I => \buf_readRTD_5\
        );

    \I__1977\ : InMux
    port map (
            O => \N__20263\,
            I => \N__20260\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__20260\,
            I => n14_adj_1577
        );

    \I__1975\ : CascadeMux
    port map (
            O => \N__20257\,
            I => \n20573_cascade_\
        );

    \I__1974\ : IoInMux
    port map (
            O => \N__20254\,
            I => \N__20251\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__20251\,
            I => \N__20248\
        );

    \I__1972\ : Span4Mux_s2_h
    port map (
            O => \N__20248\,
            I => \N__20245\
        );

    \I__1971\ : Span4Mux_h
    port map (
            O => \N__20245\,
            I => \N__20241\
        );

    \I__1970\ : CascadeMux
    port map (
            O => \N__20244\,
            I => \N__20238\
        );

    \I__1969\ : Span4Mux_v
    port map (
            O => \N__20241\,
            I => \N__20235\
        );

    \I__1968\ : InMux
    port map (
            O => \N__20238\,
            I => \N__20232\
        );

    \I__1967\ : Odrv4
    port map (
            O => \N__20235\,
            I => \VAC_CS\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__20232\,
            I => \VAC_CS\
        );

    \I__1965\ : IoInMux
    port map (
            O => \N__20227\,
            I => \N__20224\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__20224\,
            I => \N__20221\
        );

    \I__1963\ : IoSpan4Mux
    port map (
            O => \N__20221\,
            I => \N__20218\
        );

    \I__1962\ : Span4Mux_s2_h
    port map (
            O => \N__20218\,
            I => \N__20214\
        );

    \I__1961\ : CascadeMux
    port map (
            O => \N__20217\,
            I => \N__20211\
        );

    \I__1960\ : Span4Mux_h
    port map (
            O => \N__20214\,
            I => \N__20208\
        );

    \I__1959\ : InMux
    port map (
            O => \N__20211\,
            I => \N__20205\
        );

    \I__1958\ : Odrv4
    port map (
            O => \N__20208\,
            I => \VAC_SCLK\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__20205\,
            I => \VAC_SCLK\
        );

    \I__1956\ : CascadeMux
    port map (
            O => \N__20200\,
            I => \n19_adj_1622_cascade_\
        );

    \I__1955\ : InMux
    port map (
            O => \N__20197\,
            I => \N__20194\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__20194\,
            I => \N__20191\
        );

    \I__1953\ : Span4Mux_v
    port map (
            O => \N__20191\,
            I => \N__20186\
        );

    \I__1952\ : InMux
    port map (
            O => \N__20190\,
            I => \N__20181\
        );

    \I__1951\ : InMux
    port map (
            O => \N__20189\,
            I => \N__20181\
        );

    \I__1950\ : Odrv4
    port map (
            O => \N__20186\,
            I => buf_adcdata_vac_15
        );

    \I__1949\ : LocalMux
    port map (
            O => \N__20181\,
            I => buf_adcdata_vac_15
        );

    \I__1948\ : InMux
    port map (
            O => \N__20176\,
            I => \N__20173\
        );

    \I__1947\ : LocalMux
    port map (
            O => \N__20173\,
            I => \N__20170\
        );

    \I__1946\ : Span4Mux_v
    port map (
            O => \N__20170\,
            I => \N__20167\
        );

    \I__1945\ : Odrv4
    port map (
            O => \N__20167\,
            I => buf_data_iac_3
        );

    \I__1944\ : InMux
    port map (
            O => \N__20164\,
            I => \N__20161\
        );

    \I__1943\ : LocalMux
    port map (
            O => \N__20161\,
            I => \N__20158\
        );

    \I__1942\ : Span4Mux_v
    port map (
            O => \N__20158\,
            I => \N__20155\
        );

    \I__1941\ : Span4Mux_v
    port map (
            O => \N__20155\,
            I => \N__20152\
        );

    \I__1940\ : Odrv4
    port map (
            O => \N__20152\,
            I => buf_data_iac_21
        );

    \I__1939\ : CascadeMux
    port map (
            O => \N__20149\,
            I => \N__20146\
        );

    \I__1938\ : InMux
    port map (
            O => \N__20146\,
            I => \N__20139\
        );

    \I__1937\ : InMux
    port map (
            O => \N__20145\,
            I => \N__20136\
        );

    \I__1936\ : InMux
    port map (
            O => \N__20144\,
            I => \N__20133\
        );

    \I__1935\ : InMux
    port map (
            O => \N__20143\,
            I => \N__20130\
        );

    \I__1934\ : InMux
    port map (
            O => \N__20142\,
            I => \N__20127\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__20139\,
            I => \N__20120\
        );

    \I__1932\ : LocalMux
    port map (
            O => \N__20136\,
            I => \N__20120\
        );

    \I__1931\ : LocalMux
    port map (
            O => \N__20133\,
            I => \N__20120\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__20130\,
            I => \RTD.adress_7_N_1331_7\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__20127\,
            I => \RTD.adress_7_N_1331_7\
        );

    \I__1928\ : Odrv4
    port map (
            O => \N__20120\,
            I => \RTD.adress_7_N_1331_7\
        );

    \I__1927\ : InMux
    port map (
            O => \N__20113\,
            I => \N__20110\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__20110\,
            I => \N__20107\
        );

    \I__1925\ : Odrv4
    port map (
            O => \N__20107\,
            I => \RTD.n16\
        );

    \I__1924\ : CascadeMux
    port map (
            O => \N__20104\,
            I => \N__20099\
        );

    \I__1923\ : InMux
    port map (
            O => \N__20103\,
            I => \N__20093\
        );

    \I__1922\ : InMux
    port map (
            O => \N__20102\,
            I => \N__20093\
        );

    \I__1921\ : InMux
    port map (
            O => \N__20099\,
            I => \N__20088\
        );

    \I__1920\ : InMux
    port map (
            O => \N__20098\,
            I => \N__20088\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__20093\,
            I => \N__20085\
        );

    \I__1918\ : LocalMux
    port map (
            O => \N__20088\,
            I => \N__20082\
        );

    \I__1917\ : Odrv12
    port map (
            O => \N__20085\,
            I => \RTD.mode\
        );

    \I__1916\ : Odrv4
    port map (
            O => \N__20082\,
            I => \RTD.mode\
        );

    \I__1915\ : InMux
    port map (
            O => \N__20077\,
            I => \N__20074\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__20074\,
            I => \RTD.n10\
        );

    \I__1913\ : InMux
    port map (
            O => \N__20071\,
            I => \N__20065\
        );

    \I__1912\ : InMux
    port map (
            O => \N__20070\,
            I => \N__20065\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__20065\,
            I => \RTD.cfg_buf_2\
        );

    \I__1910\ : InMux
    port map (
            O => \N__20062\,
            I => \N__20056\
        );

    \I__1909\ : InMux
    port map (
            O => \N__20061\,
            I => \N__20056\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__20056\,
            I => \RTD.cfg_buf_4\
        );

    \I__1907\ : InMux
    port map (
            O => \N__20053\,
            I => \N__20047\
        );

    \I__1906\ : InMux
    port map (
            O => \N__20052\,
            I => \N__20047\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__20047\,
            I => \RTD.cfg_buf_7\
        );

    \I__1904\ : CascadeMux
    port map (
            O => \N__20044\,
            I => \N__20041\
        );

    \I__1903\ : InMux
    port map (
            O => \N__20041\,
            I => \N__20038\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__20038\,
            I => \RTD.n12\
        );

    \I__1901\ : InMux
    port map (
            O => \N__20035\,
            I => \N__20029\
        );

    \I__1900\ : InMux
    port map (
            O => \N__20034\,
            I => \N__20029\
        );

    \I__1899\ : LocalMux
    port map (
            O => \N__20029\,
            I => cfg_buf_1
        );

    \I__1898\ : InMux
    port map (
            O => \N__20026\,
            I => \N__20023\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__20023\,
            I => \N__20019\
        );

    \I__1896\ : CascadeMux
    port map (
            O => \N__20022\,
            I => \N__20016\
        );

    \I__1895\ : Span4Mux_v
    port map (
            O => \N__20019\,
            I => \N__20013\
        );

    \I__1894\ : InMux
    port map (
            O => \N__20016\,
            I => \N__20010\
        );

    \I__1893\ : Odrv4
    port map (
            O => \N__20013\,
            I => \buf_readRTD_7\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__20010\,
            I => \buf_readRTD_7\
        );

    \I__1891\ : InMux
    port map (
            O => \N__20005\,
            I => \N__20002\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__20002\,
            I => \RTD.n32\
        );

    \I__1889\ : InMux
    port map (
            O => \N__19999\,
            I => \N__19996\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__19996\,
            I => \N__19993\
        );

    \I__1887\ : Span4Mux_h
    port map (
            O => \N__19993\,
            I => \N__19989\
        );

    \I__1886\ : InMux
    port map (
            O => \N__19992\,
            I => \N__19986\
        );

    \I__1885\ : Odrv4
    port map (
            O => \N__19989\,
            I => adress_6
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__19986\,
            I => adress_6
        );

    \I__1883\ : InMux
    port map (
            O => \N__19981\,
            I => \N__19977\
        );

    \I__1882\ : InMux
    port map (
            O => \N__19980\,
            I => \N__19974\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__19977\,
            I => \N__19971\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__19974\,
            I => \RTD.adress_7\
        );

    \I__1879\ : Odrv12
    port map (
            O => \N__19971\,
            I => \RTD.adress_7\
        );

    \I__1878\ : InMux
    port map (
            O => \N__19966\,
            I => \N__19963\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__19963\,
            I => \N__19960\
        );

    \I__1876\ : Odrv12
    port map (
            O => \N__19960\,
            I => adress_0
        );

    \I__1875\ : SRMux
    port map (
            O => \N__19957\,
            I => \N__19954\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__19954\,
            I => \N__19950\
        );

    \I__1873\ : SRMux
    port map (
            O => \N__19953\,
            I => \N__19947\
        );

    \I__1872\ : Span4Mux_v
    port map (
            O => \N__19950\,
            I => \N__19942\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__19947\,
            I => \N__19942\
        );

    \I__1870\ : Span4Mux_v
    port map (
            O => \N__19942\,
            I => \N__19939\
        );

    \I__1869\ : Odrv4
    port map (
            O => \N__19939\,
            I => \RTD.n19855\
        );

    \I__1868\ : CascadeMux
    port map (
            O => \N__19936\,
            I => \RTD.adress_7_N_1331_7_cascade_\
        );

    \I__1867\ : InMux
    port map (
            O => \N__19933\,
            I => \N__19930\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__19930\,
            I => \N__19925\
        );

    \I__1865\ : InMux
    port map (
            O => \N__19929\,
            I => \N__19922\
        );

    \I__1864\ : InMux
    port map (
            O => \N__19928\,
            I => \N__19919\
        );

    \I__1863\ : Span4Mux_v
    port map (
            O => \N__19925\,
            I => \N__19912\
        );

    \I__1862\ : LocalMux
    port map (
            O => \N__19922\,
            I => \N__19912\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__19919\,
            I => \N__19912\
        );

    \I__1860\ : Span4Mux_v
    port map (
            O => \N__19912\,
            I => \N__19909\
        );

    \I__1859\ : Span4Mux_v
    port map (
            O => \N__19909\,
            I => \N__19906\
        );

    \I__1858\ : Sp12to4
    port map (
            O => \N__19906\,
            I => \N__19903\
        );

    \I__1857\ : Odrv12
    port map (
            O => \N__19903\,
            I => \RTD_DRDY\
        );

    \I__1856\ : CascadeMux
    port map (
            O => \N__19900\,
            I => \RTD.n11_cascade_\
        );

    \I__1855\ : CascadeMux
    port map (
            O => \N__19897\,
            I => \RTD.n19_cascade_\
        );

    \I__1854\ : CEMux
    port map (
            O => \N__19894\,
            I => \N__19885\
        );

    \I__1853\ : InMux
    port map (
            O => \N__19893\,
            I => \N__19872\
        );

    \I__1852\ : InMux
    port map (
            O => \N__19892\,
            I => \N__19872\
        );

    \I__1851\ : InMux
    port map (
            O => \N__19891\,
            I => \N__19872\
        );

    \I__1850\ : InMux
    port map (
            O => \N__19890\,
            I => \N__19872\
        );

    \I__1849\ : InMux
    port map (
            O => \N__19889\,
            I => \N__19872\
        );

    \I__1848\ : InMux
    port map (
            O => \N__19888\,
            I => \N__19872\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__19885\,
            I => \N__19867\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__19872\,
            I => \N__19867\
        );

    \I__1845\ : Odrv4
    port map (
            O => \N__19867\,
            I => n13151
        );

    \I__1844\ : CascadeMux
    port map (
            O => \N__19864\,
            I => \N__19860\
        );

    \I__1843\ : InMux
    port map (
            O => \N__19863\,
            I => \N__19854\
        );

    \I__1842\ : InMux
    port map (
            O => \N__19860\,
            I => \N__19854\
        );

    \I__1841\ : InMux
    port map (
            O => \N__19859\,
            I => \N__19851\
        );

    \I__1840\ : LocalMux
    port map (
            O => \N__19854\,
            I => \N__19848\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__19851\,
            I => \RTD.n1_adj_1393\
        );

    \I__1838\ : Odrv4
    port map (
            O => \N__19848\,
            I => \RTD.n1_adj_1393\
        );

    \I__1837\ : InMux
    port map (
            O => \N__19843\,
            I => \N__19840\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__19840\,
            I => \RTD.n19482\
        );

    \I__1835\ : CascadeMux
    port map (
            O => \N__19837\,
            I => \RTD.n19482_cascade_\
        );

    \I__1834\ : CascadeMux
    port map (
            O => \N__19834\,
            I => \RTD.n7285_cascade_\
        );

    \I__1833\ : CascadeMux
    port map (
            O => \N__19831\,
            I => \RTD.n21_cascade_\
        );

    \I__1832\ : InMux
    port map (
            O => \N__19828\,
            I => \N__19825\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__19825\,
            I => \N__19822\
        );

    \I__1830\ : Odrv12
    port map (
            O => \N__19822\,
            I => \RTD.n4\
        );

    \I__1829\ : CascadeMux
    port map (
            O => \N__19819\,
            I => \RTD.n20969_cascade_\
        );

    \I__1828\ : SRMux
    port map (
            O => \N__19816\,
            I => \N__19813\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__19813\,
            I => \N__19809\
        );

    \I__1826\ : SRMux
    port map (
            O => \N__19812\,
            I => \N__19806\
        );

    \I__1825\ : Span4Mux_h
    port map (
            O => \N__19809\,
            I => \N__19801\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__19806\,
            I => \N__19801\
        );

    \I__1823\ : Odrv4
    port map (
            O => \N__19801\,
            I => \RTD.n15050\
        );

    \I__1822\ : IoInMux
    port map (
            O => \N__19798\,
            I => \N__19795\
        );

    \I__1821\ : LocalMux
    port map (
            O => \N__19795\,
            I => \N__19792\
        );

    \I__1820\ : IoSpan4Mux
    port map (
            O => \N__19792\,
            I => \N__19789\
        );

    \I__1819\ : Span4Mux_s3_h
    port map (
            O => \N__19789\,
            I => \N__19786\
        );

    \I__1818\ : Span4Mux_v
    port map (
            O => \N__19786\,
            I => \N__19783\
        );

    \I__1817\ : Sp12to4
    port map (
            O => \N__19783\,
            I => \N__19780\
        );

    \I__1816\ : Odrv12
    port map (
            O => \N__19780\,
            I => \RTD_SDI\
        );

    \I__1815\ : CEMux
    port map (
            O => \N__19777\,
            I => \N__19774\
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__19774\,
            I => \N__19771\
        );

    \I__1813\ : Span4Mux_v
    port map (
            O => \N__19771\,
            I => \N__19768\
        );

    \I__1812\ : Span4Mux_h
    port map (
            O => \N__19768\,
            I => \N__19765\
        );

    \I__1811\ : Odrv4
    port map (
            O => \N__19765\,
            I => \RTD.n11704\
        );

    \I__1810\ : CascadeMux
    port map (
            O => \N__19762\,
            I => \RTD.n33_cascade_\
        );

    \I__1809\ : CascadeMux
    port map (
            O => \N__19759\,
            I => \N__19752\
        );

    \I__1808\ : CascadeMux
    port map (
            O => \N__19758\,
            I => \N__19746\
        );

    \I__1807\ : CascadeMux
    port map (
            O => \N__19757\,
            I => \N__19741\
        );

    \I__1806\ : CascadeMux
    port map (
            O => \N__19756\,
            I => \N__19738\
        );

    \I__1805\ : InMux
    port map (
            O => \N__19755\,
            I => \N__19729\
        );

    \I__1804\ : InMux
    port map (
            O => \N__19752\,
            I => \N__19726\
        );

    \I__1803\ : InMux
    port map (
            O => \N__19751\,
            I => \N__19723\
        );

    \I__1802\ : InMux
    port map (
            O => \N__19750\,
            I => \N__19720\
        );

    \I__1801\ : InMux
    port map (
            O => \N__19749\,
            I => \N__19717\
        );

    \I__1800\ : InMux
    port map (
            O => \N__19746\,
            I => \N__19712\
        );

    \I__1799\ : InMux
    port map (
            O => \N__19745\,
            I => \N__19712\
        );

    \I__1798\ : InMux
    port map (
            O => \N__19744\,
            I => \N__19703\
        );

    \I__1797\ : InMux
    port map (
            O => \N__19741\,
            I => \N__19703\
        );

    \I__1796\ : InMux
    port map (
            O => \N__19738\,
            I => \N__19703\
        );

    \I__1795\ : InMux
    port map (
            O => \N__19737\,
            I => \N__19703\
        );

    \I__1794\ : InMux
    port map (
            O => \N__19736\,
            I => \N__19692\
        );

    \I__1793\ : InMux
    port map (
            O => \N__19735\,
            I => \N__19692\
        );

    \I__1792\ : InMux
    port map (
            O => \N__19734\,
            I => \N__19692\
        );

    \I__1791\ : InMux
    port map (
            O => \N__19733\,
            I => \N__19692\
        );

    \I__1790\ : InMux
    port map (
            O => \N__19732\,
            I => \N__19692\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__19729\,
            I => \N__19689\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__19726\,
            I => \N__19674\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__19723\,
            I => \N__19674\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__19720\,
            I => \N__19674\
        );

    \I__1785\ : LocalMux
    port map (
            O => \N__19717\,
            I => \N__19674\
        );

    \I__1784\ : LocalMux
    port map (
            O => \N__19712\,
            I => \N__19674\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__19703\,
            I => \N__19674\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__19692\,
            I => \N__19674\
        );

    \I__1781\ : Span4Mux_v
    port map (
            O => \N__19689\,
            I => \N__19669\
        );

    \I__1780\ : Span4Mux_v
    port map (
            O => \N__19674\,
            I => \N__19669\
        );

    \I__1779\ : Odrv4
    port map (
            O => \N__19669\,
            I => n1_adj_1575
        );

    \I__1778\ : InMux
    port map (
            O => \N__19666\,
            I => \N__19663\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__19663\,
            I => \N__19660\
        );

    \I__1776\ : Odrv12
    port map (
            O => \N__19660\,
            I => \RTD.n16614\
        );

    \I__1775\ : CascadeMux
    port map (
            O => \N__19657\,
            I => \RTD.n16614_cascade_\
        );

    \I__1774\ : CascadeMux
    port map (
            O => \N__19654\,
            I => \N__19648\
        );

    \I__1773\ : CascadeMux
    port map (
            O => \N__19653\,
            I => \N__19645\
        );

    \I__1772\ : CascadeMux
    port map (
            O => \N__19652\,
            I => \N__19642\
        );

    \I__1771\ : CascadeMux
    port map (
            O => \N__19651\,
            I => \N__19637\
        );

    \I__1770\ : InMux
    port map (
            O => \N__19648\,
            I => \N__19626\
        );

    \I__1769\ : InMux
    port map (
            O => \N__19645\,
            I => \N__19626\
        );

    \I__1768\ : InMux
    port map (
            O => \N__19642\,
            I => \N__19626\
        );

    \I__1767\ : InMux
    port map (
            O => \N__19641\,
            I => \N__19626\
        );

    \I__1766\ : InMux
    port map (
            O => \N__19640\,
            I => \N__19626\
        );

    \I__1765\ : InMux
    port map (
            O => \N__19637\,
            I => \N__19623\
        );

    \I__1764\ : LocalMux
    port map (
            O => \N__19626\,
            I => n14465
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__19623\,
            I => n14465
        );

    \I__1762\ : InMux
    port map (
            O => \N__19618\,
            I => \N__19613\
        );

    \I__1761\ : InMux
    port map (
            O => \N__19617\,
            I => \N__19610\
        );

    \I__1760\ : InMux
    port map (
            O => \N__19616\,
            I => \N__19607\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__19613\,
            I => read_buf_8
        );

    \I__1758\ : LocalMux
    port map (
            O => \N__19610\,
            I => read_buf_8
        );

    \I__1757\ : LocalMux
    port map (
            O => \N__19607\,
            I => read_buf_8
        );

    \I__1756\ : CascadeMux
    port map (
            O => \N__19600\,
            I => \N__19597\
        );

    \I__1755\ : InMux
    port map (
            O => \N__19597\,
            I => \N__19592\
        );

    \I__1754\ : InMux
    port map (
            O => \N__19596\,
            I => \N__19589\
        );

    \I__1753\ : InMux
    port map (
            O => \N__19595\,
            I => \N__19586\
        );

    \I__1752\ : LocalMux
    port map (
            O => \N__19592\,
            I => read_buf_4
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__19589\,
            I => read_buf_4
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__19586\,
            I => read_buf_4
        );

    \I__1749\ : InMux
    port map (
            O => \N__19579\,
            I => \N__19569\
        );

    \I__1748\ : InMux
    port map (
            O => \N__19578\,
            I => \N__19569\
        );

    \I__1747\ : InMux
    port map (
            O => \N__19577\,
            I => \N__19563\
        );

    \I__1746\ : InMux
    port map (
            O => \N__19576\,
            I => \N__19563\
        );

    \I__1745\ : InMux
    port map (
            O => \N__19575\,
            I => \N__19553\
        );

    \I__1744\ : InMux
    port map (
            O => \N__19574\,
            I => \N__19553\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__19569\,
            I => \N__19547\
        );

    \I__1742\ : InMux
    port map (
            O => \N__19568\,
            I => \N__19544\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__19563\,
            I => \N__19541\
        );

    \I__1740\ : InMux
    port map (
            O => \N__19562\,
            I => \N__19530\
        );

    \I__1739\ : InMux
    port map (
            O => \N__19561\,
            I => \N__19530\
        );

    \I__1738\ : InMux
    port map (
            O => \N__19560\,
            I => \N__19530\
        );

    \I__1737\ : InMux
    port map (
            O => \N__19559\,
            I => \N__19530\
        );

    \I__1736\ : InMux
    port map (
            O => \N__19558\,
            I => \N__19530\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__19553\,
            I => \N__19527\
        );

    \I__1734\ : InMux
    port map (
            O => \N__19552\,
            I => \N__19520\
        );

    \I__1733\ : InMux
    port map (
            O => \N__19551\,
            I => \N__19520\
        );

    \I__1732\ : InMux
    port map (
            O => \N__19550\,
            I => \N__19520\
        );

    \I__1731\ : Odrv4
    port map (
            O => \N__19547\,
            I => n13279
        );

    \I__1730\ : LocalMux
    port map (
            O => \N__19544\,
            I => n13279
        );

    \I__1729\ : Odrv4
    port map (
            O => \N__19541\,
            I => n13279
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__19530\,
            I => n13279
        );

    \I__1727\ : Odrv4
    port map (
            O => \N__19527\,
            I => n13279
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__19520\,
            I => n13279
        );

    \I__1725\ : InMux
    port map (
            O => \N__19507\,
            I => \N__19500\
        );

    \I__1724\ : InMux
    port map (
            O => \N__19506\,
            I => \N__19500\
        );

    \I__1723\ : InMux
    port map (
            O => \N__19505\,
            I => \N__19497\
        );

    \I__1722\ : LocalMux
    port map (
            O => \N__19500\,
            I => read_buf_2
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__19497\,
            I => read_buf_2
        );

    \I__1720\ : CascadeMux
    port map (
            O => \N__19492\,
            I => \N__19488\
        );

    \I__1719\ : InMux
    port map (
            O => \N__19491\,
            I => \N__19484\
        );

    \I__1718\ : InMux
    port map (
            O => \N__19488\,
            I => \N__19479\
        );

    \I__1717\ : InMux
    port map (
            O => \N__19487\,
            I => \N__19479\
        );

    \I__1716\ : LocalMux
    port map (
            O => \N__19484\,
            I => read_buf_3
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__19479\,
            I => read_buf_3
        );

    \I__1714\ : CascadeMux
    port map (
            O => \N__19474\,
            I => \N__19469\
        );

    \I__1713\ : InMux
    port map (
            O => \N__19473\,
            I => \N__19461\
        );

    \I__1712\ : InMux
    port map (
            O => \N__19472\,
            I => \N__19461\
        );

    \I__1711\ : InMux
    port map (
            O => \N__19469\,
            I => \N__19448\
        );

    \I__1710\ : InMux
    port map (
            O => \N__19468\,
            I => \N__19448\
        );

    \I__1709\ : InMux
    port map (
            O => \N__19467\,
            I => \N__19448\
        );

    \I__1708\ : InMux
    port map (
            O => \N__19466\,
            I => \N__19448\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__19461\,
            I => \N__19444\
        );

    \I__1706\ : InMux
    port map (
            O => \N__19460\,
            I => \N__19437\
        );

    \I__1705\ : InMux
    port map (
            O => \N__19459\,
            I => \N__19437\
        );

    \I__1704\ : InMux
    port map (
            O => \N__19458\,
            I => \N__19437\
        );

    \I__1703\ : InMux
    port map (
            O => \N__19457\,
            I => \N__19434\
        );

    \I__1702\ : LocalMux
    port map (
            O => \N__19448\,
            I => \N__19427\
        );

    \I__1701\ : InMux
    port map (
            O => \N__19447\,
            I => \N__19424\
        );

    \I__1700\ : Span4Mux_v
    port map (
            O => \N__19444\,
            I => \N__19417\
        );

    \I__1699\ : LocalMux
    port map (
            O => \N__19437\,
            I => \N__19417\
        );

    \I__1698\ : LocalMux
    port map (
            O => \N__19434\,
            I => \N__19417\
        );

    \I__1697\ : InMux
    port map (
            O => \N__19433\,
            I => \N__19410\
        );

    \I__1696\ : InMux
    port map (
            O => \N__19432\,
            I => \N__19410\
        );

    \I__1695\ : InMux
    port map (
            O => \N__19431\,
            I => \N__19410\
        );

    \I__1694\ : InMux
    port map (
            O => \N__19430\,
            I => \N__19407\
        );

    \I__1693\ : Odrv12
    port map (
            O => \N__19427\,
            I => n11700
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__19424\,
            I => n11700
        );

    \I__1691\ : Odrv4
    port map (
            O => \N__19417\,
            I => n11700
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__19410\,
            I => n11700
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__19407\,
            I => n11700
        );

    \I__1688\ : CEMux
    port map (
            O => \N__19396\,
            I => \N__19393\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__19393\,
            I => \N__19390\
        );

    \I__1686\ : Span4Mux_h
    port map (
            O => \N__19390\,
            I => \N__19386\
        );

    \I__1685\ : CEMux
    port map (
            O => \N__19389\,
            I => \N__19383\
        );

    \I__1684\ : Odrv4
    port map (
            O => \N__19386\,
            I => \RTD.n11726\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__19383\,
            I => \RTD.n11726\
        );

    \I__1682\ : InMux
    port map (
            O => \N__19378\,
            I => \N__19373\
        );

    \I__1681\ : InMux
    port map (
            O => \N__19377\,
            I => \N__19370\
        );

    \I__1680\ : InMux
    port map (
            O => \N__19376\,
            I => \N__19367\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__19373\,
            I => read_buf_13
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__19370\,
            I => read_buf_13
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__19367\,
            I => read_buf_13
        );

    \I__1676\ : CascadeMux
    port map (
            O => \N__19360\,
            I => \N__19356\
        );

    \I__1675\ : InMux
    port map (
            O => \N__19359\,
            I => \N__19348\
        );

    \I__1674\ : InMux
    port map (
            O => \N__19356\,
            I => \N__19348\
        );

    \I__1673\ : InMux
    port map (
            O => \N__19355\,
            I => \N__19348\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__19348\,
            I => read_buf_9
        );

    \I__1671\ : InMux
    port map (
            O => \N__19345\,
            I => \N__19339\
        );

    \I__1670\ : InMux
    port map (
            O => \N__19344\,
            I => \N__19339\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__19339\,
            I => adress_1
        );

    \I__1668\ : InMux
    port map (
            O => \N__19336\,
            I => \N__19330\
        );

    \I__1667\ : InMux
    port map (
            O => \N__19335\,
            I => \N__19330\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__19330\,
            I => adress_2
        );

    \I__1665\ : CascadeMux
    port map (
            O => \N__19327\,
            I => \N__19323\
        );

    \I__1664\ : InMux
    port map (
            O => \N__19326\,
            I => \N__19318\
        );

    \I__1663\ : InMux
    port map (
            O => \N__19323\,
            I => \N__19318\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__19318\,
            I => adress_3
        );

    \I__1661\ : InMux
    port map (
            O => \N__19315\,
            I => \N__19309\
        );

    \I__1660\ : InMux
    port map (
            O => \N__19314\,
            I => \N__19309\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__19309\,
            I => \N__19306\
        );

    \I__1658\ : Odrv4
    port map (
            O => \N__19306\,
            I => adress_4
        );

    \I__1657\ : CascadeMux
    port map (
            O => \N__19303\,
            I => \N__19299\
        );

    \I__1656\ : InMux
    port map (
            O => \N__19302\,
            I => \N__19294\
        );

    \I__1655\ : InMux
    port map (
            O => \N__19299\,
            I => \N__19294\
        );

    \I__1654\ : LocalMux
    port map (
            O => \N__19294\,
            I => adress_5
        );

    \I__1653\ : CascadeMux
    port map (
            O => \N__19291\,
            I => \N__19287\
        );

    \I__1652\ : InMux
    port map (
            O => \N__19290\,
            I => \N__19283\
        );

    \I__1651\ : InMux
    port map (
            O => \N__19287\,
            I => \N__19280\
        );

    \I__1650\ : InMux
    port map (
            O => \N__19286\,
            I => \N__19277\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__19283\,
            I => read_buf_10
        );

    \I__1648\ : LocalMux
    port map (
            O => \N__19280\,
            I => read_buf_10
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__19277\,
            I => read_buf_10
        );

    \I__1646\ : InMux
    port map (
            O => \N__19270\,
            I => \N__19265\
        );

    \I__1645\ : CascadeMux
    port map (
            O => \N__19269\,
            I => \N__19262\
        );

    \I__1644\ : CascadeMux
    port map (
            O => \N__19268\,
            I => \N__19259\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__19265\,
            I => \N__19256\
        );

    \I__1642\ : InMux
    port map (
            O => \N__19262\,
            I => \N__19251\
        );

    \I__1641\ : InMux
    port map (
            O => \N__19259\,
            I => \N__19251\
        );

    \I__1640\ : Odrv4
    port map (
            O => \N__19256\,
            I => read_buf_11
        );

    \I__1639\ : LocalMux
    port map (
            O => \N__19251\,
            I => read_buf_11
        );

    \I__1638\ : CascadeMux
    port map (
            O => \N__19246\,
            I => \n11700_cascade_\
        );

    \I__1637\ : CascadeMux
    port map (
            O => \N__19243\,
            I => \N__19240\
        );

    \I__1636\ : InMux
    port map (
            O => \N__19240\,
            I => \N__19233\
        );

    \I__1635\ : InMux
    port map (
            O => \N__19239\,
            I => \N__19233\
        );

    \I__1634\ : InMux
    port map (
            O => \N__19238\,
            I => \N__19230\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__19233\,
            I => read_buf_14
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__19230\,
            I => read_buf_14
        );

    \I__1631\ : InMux
    port map (
            O => \N__19225\,
            I => \N__19219\
        );

    \I__1630\ : InMux
    port map (
            O => \N__19224\,
            I => \N__19219\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__19219\,
            I => read_buf_15
        );

    \I__1628\ : CascadeMux
    port map (
            O => \N__19216\,
            I => \N__19213\
        );

    \I__1627\ : InMux
    port map (
            O => \N__19213\,
            I => \N__19210\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__19210\,
            I => \N__19205\
        );

    \I__1625\ : InMux
    port map (
            O => \N__19209\,
            I => \N__19202\
        );

    \I__1624\ : InMux
    port map (
            O => \N__19208\,
            I => \N__19199\
        );

    \I__1623\ : Odrv12
    port map (
            O => \N__19205\,
            I => read_buf_1
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__19202\,
            I => read_buf_1
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__19199\,
            I => read_buf_1
        );

    \I__1620\ : InMux
    port map (
            O => \N__19192\,
            I => \N__19187\
        );

    \I__1619\ : InMux
    port map (
            O => \N__19191\,
            I => \N__19182\
        );

    \I__1618\ : InMux
    port map (
            O => \N__19190\,
            I => \N__19182\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__19187\,
            I => read_buf_0
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__19182\,
            I => read_buf_0
        );

    \I__1615\ : InMux
    port map (
            O => \N__19177\,
            I => \N__19172\
        );

    \I__1614\ : InMux
    port map (
            O => \N__19176\,
            I => \N__19167\
        );

    \I__1613\ : InMux
    port map (
            O => \N__19175\,
            I => \N__19167\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__19172\,
            I => read_buf_5
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__19167\,
            I => read_buf_5
        );

    \I__1610\ : CascadeMux
    port map (
            O => \N__19162\,
            I => \N__19158\
        );

    \I__1609\ : InMux
    port map (
            O => \N__19161\,
            I => \N__19154\
        );

    \I__1608\ : InMux
    port map (
            O => \N__19158\,
            I => \N__19149\
        );

    \I__1607\ : InMux
    port map (
            O => \N__19157\,
            I => \N__19149\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__19154\,
            I => read_buf_12
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__19149\,
            I => read_buf_12
        );

    \I__1604\ : CascadeMux
    port map (
            O => \N__19144\,
            I => \N__19141\
        );

    \I__1603\ : InMux
    port map (
            O => \N__19141\,
            I => \N__19135\
        );

    \I__1602\ : InMux
    port map (
            O => \N__19140\,
            I => \N__19135\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__19135\,
            I => \N__19131\
        );

    \I__1600\ : InMux
    port map (
            O => \N__19134\,
            I => \N__19128\
        );

    \I__1599\ : Odrv4
    port map (
            O => \N__19131\,
            I => read_buf_6
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__19128\,
            I => read_buf_6
        );

    \I__1597\ : InMux
    port map (
            O => \N__19123\,
            I => \N__19119\
        );

    \I__1596\ : CascadeMux
    port map (
            O => \N__19122\,
            I => \N__19116\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__19119\,
            I => \N__19112\
        );

    \I__1594\ : InMux
    port map (
            O => \N__19116\,
            I => \N__19109\
        );

    \I__1593\ : InMux
    port map (
            O => \N__19115\,
            I => \N__19106\
        );

    \I__1592\ : Odrv4
    port map (
            O => \N__19112\,
            I => read_buf_7
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__19109\,
            I => read_buf_7
        );

    \I__1590\ : LocalMux
    port map (
            O => \N__19106\,
            I => read_buf_7
        );

    \I__1589\ : IoInMux
    port map (
            O => \N__19099\,
            I => \N__19096\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__19096\,
            I => \N__19093\
        );

    \I__1587\ : IoSpan4Mux
    port map (
            O => \N__19093\,
            I => \N__19090\
        );

    \I__1586\ : Span4Mux_s3_h
    port map (
            O => \N__19090\,
            I => \N__19087\
        );

    \I__1585\ : Span4Mux_v
    port map (
            O => \N__19087\,
            I => \N__19084\
        );

    \I__1584\ : Span4Mux_v
    port map (
            O => \N__19084\,
            I => \N__19081\
        );

    \I__1583\ : Odrv4
    port map (
            O => \N__19081\,
            I => \RTD_CS\
        );

    \I__1582\ : CEMux
    port map (
            O => \N__19078\,
            I => \N__19075\
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__19075\,
            I => \N__19072\
        );

    \I__1580\ : Odrv12
    port map (
            O => \N__19072\,
            I => \RTD.n11673\
        );

    \I__1579\ : CascadeMux
    port map (
            O => \N__19069\,
            I => \n13279_cascade_\
        );

    \I__1578\ : CascadeMux
    port map (
            O => \N__19066\,
            I => \N__19063\
        );

    \I__1577\ : InMux
    port map (
            O => \N__19063\,
            I => \N__19060\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__19060\,
            I => \N__19057\
        );

    \I__1575\ : Span4Mux_h
    port map (
            O => \N__19057\,
            I => \N__19054\
        );

    \I__1574\ : Sp12to4
    port map (
            O => \N__19054\,
            I => \N__19051\
        );

    \I__1573\ : Span12Mux_v
    port map (
            O => \N__19051\,
            I => \N__19048\
        );

    \I__1572\ : Odrv12
    port map (
            O => \N__19048\,
            I => \RTD_SDO\
        );

    \I__1571\ : IoInMux
    port map (
            O => \N__19045\,
            I => \N__19042\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__19042\,
            I => \N__19039\
        );

    \I__1569\ : IoSpan4Mux
    port map (
            O => \N__19039\,
            I => \N__19036\
        );

    \I__1568\ : Span4Mux_s3_h
    port map (
            O => \N__19036\,
            I => \N__19033\
        );

    \I__1567\ : Span4Mux_v
    port map (
            O => \N__19033\,
            I => \N__19030\
        );

    \I__1566\ : Odrv4
    port map (
            O => \N__19030\,
            I => \RTD_SCLK\
        );

    \I__1565\ : CEMux
    port map (
            O => \N__19027\,
            I => \N__19024\
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__19024\,
            I => \N__19021\
        );

    \I__1563\ : Odrv4
    port map (
            O => \N__19021\,
            I => \RTD.n8\
        );

    \I__1562\ : IoInMux
    port map (
            O => \N__19018\,
            I => \N__19015\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__19015\,
            I => \N__19012\
        );

    \I__1560\ : IoSpan4Mux
    port map (
            O => \N__19012\,
            I => \N__19009\
        );

    \I__1559\ : IoSpan4Mux
    port map (
            O => \N__19009\,
            I => \N__19006\
        );

    \I__1558\ : Odrv4
    port map (
            O => \N__19006\,
            I => \ICE_SYSCLK\
        );

    \I__1557\ : IoInMux
    port map (
            O => \N__19003\,
            I => \N__19000\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__19000\,
            I => \N__18997\
        );

    \I__1555\ : IoSpan4Mux
    port map (
            O => \N__18997\,
            I => \N__18994\
        );

    \I__1554\ : Span4Mux_s3_v
    port map (
            O => \N__18994\,
            I => \N__18991\
        );

    \I__1553\ : Sp12to4
    port map (
            O => \N__18991\,
            I => \N__18988\
        );

    \I__1552\ : Span12Mux_h
    port map (
            O => \N__18988\,
            I => \N__18985\
        );

    \I__1551\ : Odrv12
    port map (
            O => \N__18985\,
            I => \ICE_GPMO_2\
        );

    \INVdds0_mclkcnt_i7_3772__i0C\ : INV
    port map (
            O => \INVdds0_mclkcnt_i7_3772__i0C_net\,
            I => \N__56030\
        );

    \INVdds0_mclk_294C\ : INV
    port map (
            O => \INVdds0_mclk_294C_net\,
            I => \N__56029\
        );

    \INVdata_cntvec_i0_i8C\ : INV
    port map (
            O => \INVdata_cntvec_i0_i8C_net\,
            I => \N__55186\
        );

    \INVdata_cntvec_i0_i0C\ : INV
    port map (
            O => \INVdata_cntvec_i0_i0C_net\,
            I => \N__55172\
        );

    \INVcomm_spi.data_valid_85C\ : INV
    port map (
            O => \INVcomm_spi.data_valid_85C_net\,
            I => \N__55130\
        );

    \INVcomm_spi.MISO_48_12187_12188_resetC\ : INV
    port map (
            O => \INVcomm_spi.MISO_48_12187_12188_resetC_net\,
            I => \N__55090\
        );

    \INVcomm_spi.imiso_83_12193_12194_resetC\ : INV
    port map (
            O => \INVcomm_spi.imiso_83_12193_12194_resetC_net\,
            I => \N__52368\
        );

    \INVdata_count_i0_i8C\ : INV
    port map (
            O => \INVdata_count_i0_i8C_net\,
            I => \N__55211\
        );

    \INVdata_count_i0_i0C\ : INV
    port map (
            O => \INVdata_count_i0_i0C_net\,
            I => \N__55198\
        );

    \INVcomm_spi.MISO_48_12187_12188_setC\ : INV
    port map (
            O => \INVcomm_spi.MISO_48_12187_12188_setC_net\,
            I => \N__55078\
        );

    \INVADC_VDC.genclk.t0on_i8C\ : INV
    port map (
            O => \INVADC_VDC.genclk.t0on_i8C_net\,
            I => \N__56022\
        );

    \INVADC_VDC.genclk.t0on_i0C\ : INV
    port map (
            O => \INVADC_VDC.genclk.t0on_i0C_net\,
            I => \N__56018\
        );

    \INVADC_VDC.genclk.div_state_i1C\ : INV
    port map (
            O => \INVADC_VDC.genclk.div_state_i1C_net\,
            I => \N__56023\
        );

    \INVacadc_skipcnt_i0_i9C\ : INV
    port map (
            O => \INVacadc_skipcnt_i0_i9C_net\,
            I => \N__55182\
        );

    \INVacadc_skipcnt_i0_i1C\ : INV
    port map (
            O => \INVacadc_skipcnt_i0_i1C_net\,
            I => \N__55167\
        );

    \INVacadc_skipcnt_i0_i0C\ : INV
    port map (
            O => \INVacadc_skipcnt_i0_i0C_net\,
            I => \N__55152\
        );

    \INVcomm_spi.bit_cnt_3767__i1C\ : INV
    port map (
            O => \INVcomm_spi.bit_cnt_3767__i1C_net\,
            I => \N__52414\
        );

    \INVcomm_spi.imiso_83_12193_12194_setC\ : INV
    port map (
            O => \INVcomm_spi.imiso_83_12193_12194_setC_net\,
            I => \N__52413\
        );

    \INVADC_VDC.genclk.t_clk_24C\ : INV
    port map (
            O => \INVADC_VDC.genclk.t_clk_24C_net\,
            I => \N__56016\
        );

    \INVacadc_trig_300C\ : INV
    port map (
            O => \INVacadc_trig_300C_net\,
            I => \N__55181\
        );

    \INVeis_state_i0C\ : INV
    port map (
            O => \INVeis_state_i0C_net\,
            I => \N__55117\
        );

    \INVADC_VDC.genclk.t0off_i8C\ : INV
    port map (
            O => \INVADC_VDC.genclk.t0off_i8C_net\,
            I => \N__56017\
        );

    \INVADC_VDC.genclk.t0off_i0C\ : INV
    port map (
            O => \INVADC_VDC.genclk.t0off_i0C_net\,
            I => \N__56015\
        );

    \INViac_raw_buf_vac_raw_buf_merged2WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged2WCLKN_net\,
            I => \N__55159\
        );

    \INViac_raw_buf_vac_raw_buf_merged7WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged7WCLKN_net\,
            I => \N__55246\
        );

    \INViac_raw_buf_vac_raw_buf_merged1WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged1WCLKN_net\,
            I => \N__55092\
        );

    \INViac_raw_buf_vac_raw_buf_merged6WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged6WCLKN_net\,
            I => \N__55243\
        );

    \INViac_raw_buf_vac_raw_buf_merged0WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged0WCLKN_net\,
            I => \N__55080\
        );

    \INViac_raw_buf_vac_raw_buf_merged5WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged5WCLKN_net\,
            I => \N__55236\
        );

    \INViac_raw_buf_vac_raw_buf_merged9WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged9WCLKN_net\,
            I => \N__55226\
        );

    \INViac_raw_buf_vac_raw_buf_merged4WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged4WCLKN_net\,
            I => \N__55215\
        );

    \INViac_raw_buf_vac_raw_buf_merged8WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged8WCLKN_net\,
            I => \N__55203\
        );

    \INViac_raw_buf_vac_raw_buf_merged10WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged10WCLKN_net\,
            I => \N__55111\
        );

    \INViac_raw_buf_vac_raw_buf_merged3WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged3WCLKN_net\,
            I => \N__55189\
        );

    \INViac_raw_buf_vac_raw_buf_merged11WCLKN\ : INV
    port map (
            O => \INViac_raw_buf_vac_raw_buf_merged11WCLKN_net\,
            I => \N__55132\
        );

    \IN_MUX_bfv_17_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_17_9_0_\
        );

    \IN_MUX_bfv_17_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n19454,
            carryinitout => \bfn_17_10_0_\
        );

    \IN_MUX_bfv_17_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n19462,
            carryinitout => \bfn_17_11_0_\
        );

    \IN_MUX_bfv_22_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_22_11_0_\
        );

    \IN_MUX_bfv_13_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_16_0_\
        );

    \IN_MUX_bfv_13_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \n19311_THRU_CRY_6_THRU_CO\,
            carryinitout => \bfn_13_17_0_\
        );

    \IN_MUX_bfv_13_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n19319,
            carryinitout => \bfn_13_18_0_\
        );

    \IN_MUX_bfv_18_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_12_0_\
        );

    \IN_MUX_bfv_18_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n19303,
            carryinitout => \bfn_18_13_0_\
        );

    \IN_MUX_bfv_15_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_17_0_\
        );

    \IN_MUX_bfv_15_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n19294,
            carryinitout => \bfn_15_18_0_\
        );

    \IN_MUX_bfv_12_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_12_0_\
        );

    \IN_MUX_bfv_12_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n19342,
            carryinitout => \bfn_12_13_0_\
        );

    \IN_MUX_bfv_16_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_16_15_0_\
        );

    \IN_MUX_bfv_16_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n19333,
            carryinitout => \bfn_16_16_0_\
        );

    \IN_MUX_bfv_11_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_3_0_\
        );

    \IN_MUX_bfv_11_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ADC_VDC.genclk.n19417\,
            carryinitout => \bfn_11_4_0_\
        );

    \IN_MUX_bfv_15_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_15_3_0_\
        );

    \IN_MUX_bfv_15_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ADC_VDC.genclk.n19432\,
            carryinitout => \bfn_15_4_0_\
        );

    \IN_MUX_bfv_13_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_6_0_\
        );

    \IN_MUX_bfv_11_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_7_0_\
        );

    \IN_MUX_bfv_11_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ADC_VDC.n19406\,
            carryinitout => \bfn_11_8_0_\
        );

    \IN_MUX_bfv_9_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_5_0_\
        );

    \IN_MUX_bfv_9_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ADC_VDC.n19371\,
            carryinitout => \bfn_9_6_0_\
        );

    \IN_MUX_bfv_9_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ADC_VDC.n19379\,
            carryinitout => \bfn_9_7_0_\
        );

    \IN_MUX_bfv_9_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ADC_VDC.n19387\,
            carryinitout => \bfn_9_8_0_\
        );

    \IN_MUX_bfv_9_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ADC_VDC.n19395\,
            carryinitout => \bfn_9_9_0_\
        );

    \IN_MUX_bfv_7_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_17_0_\
        );

    \IN_MUX_bfv_7_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_19_0_\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \RTD.SCLK_51_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010110000110110"
        )
    port map (
            in0 => \N__22257\,
            in1 => \N__22114\,
            in2 => \N__22410\,
            in3 => \N__20970\,
            lcout => \RTD_SCLK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41081\,
            ce => \N__19027\,
            sr => \_gnd_net_\
        );

    \RTD.i19108_4_lut_4_lut_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011110111111"
        )
    port map (
            in0 => \N__20969\,
            in1 => \N__22393\,
            in2 => \N__22132\,
            in3 => \N__22255\,
            lcout => \RTD.n8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i27_4_lut_4_lut_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010000110"
        )
    port map (
            in0 => \N__22254\,
            in1 => \N__22109\,
            in2 => \N__22409\,
            in3 => \N__20968\,
            lcout => \RTD.n11704\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i19151_4_lut_4_lut_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101001110101100"
        )
    port map (
            in0 => \N__20966\,
            in1 => \N__22394\,
            in2 => \N__22131\,
            in3 => \N__22253\,
            lcout => \RTD.n11726\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_3_lut_4_lut_adj_25_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010010010010"
        )
    port map (
            in0 => \N__22252\,
            in1 => \N__22105\,
            in2 => \N__22408\,
            in3 => \N__20967\,
            lcout => \RTD.n15050\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i19070_3_lut_3_lut_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010011001"
        )
    port map (
            in0 => \N__22113\,
            in1 => \N__22395\,
            in2 => \_gnd_net_\,
            in3 => \N__22256\,
            lcout => \RTD.n11673\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.CS_52_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011101010111"
        )
    port map (
            in0 => \N__20964\,
            in1 => \N__19666\,
            in2 => \N__22411\,
            in3 => \N__22258\,
            lcout => \RTD_CS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41131\,
            ce => \N__19078\,
            sr => \_gnd_net_\
        );

    \RTD.i1_4_lut_4_lut_adj_21_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100100000001"
        )
    port map (
            in0 => \N__22259\,
            in1 => \N__22118\,
            in2 => \N__20977\,
            in3 => \N__22403\,
            lcout => n13279,
            ltout => \n13279_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i14_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__19377\,
            in1 => \N__19238\,
            in2 => \N__19069\,
            in3 => \N__19744\,
            lcout => read_buf_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41143\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i7_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__22119\,
            in1 => \N__19447\,
            in2 => \N__20022\,
            in3 => \N__19123\,
            lcout => \buf_readRTD_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41143\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i1_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__19551\,
            in1 => \N__19191\,
            in2 => \N__19756\,
            in3 => \N__19208\,
            lcout => read_buf_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41143\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i6_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__19552\,
            in1 => \N__19177\,
            in2 => \N__19757\,
            in3 => \N__19134\,
            lcout => read_buf_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41143\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i0_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__19190\,
            in1 => \N__19737\,
            in2 => \N__19066\,
            in3 => \N__19550\,
            lcout => read_buf_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41143\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i11_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__19733\,
            in1 => \N__19286\,
            in2 => \N__19268\,
            in3 => \N__19558\,
            lcout => read_buf_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41080\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i13_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__19560\,
            in1 => \N__19376\,
            in2 => \N__19162\,
            in3 => \N__19736\,
            lcout => read_buf_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41080\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i5_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__19735\,
            in1 => \N__19175\,
            in2 => \N__19600\,
            in3 => \N__19561\,
            lcout => read_buf_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41080\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i8_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__19562\,
            in1 => \N__19616\,
            in2 => \N__19122\,
            in3 => \N__19732\,
            lcout => read_buf_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41080\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i12_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__19734\,
            in1 => \N__19157\,
            in2 => \N__19269\,
            in3 => \N__19559\,
            lcout => read_buf_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41080\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i0_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__22120\,
            in1 => \N__19192\,
            in2 => \N__21366\,
            in3 => \N__19458\,
            lcout => \buf_readRTD_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41080\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i5_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__19460\,
            in1 => \N__19176\,
            in2 => \N__20280\,
            in3 => \N__22122\,
            lcout => \buf_readRTD_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41080\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i12_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__22121\,
            in1 => \N__19161\,
            in2 => \N__25746\,
            in3 => \N__19459\,
            lcout => \buf_readRTD_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41080\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i6_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__19140\,
            in1 => \N__19473\,
            in2 => \N__29607\,
            in3 => \N__22129\,
            lcout => \buf_readRTD_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41130\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i7_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__19577\,
            in1 => \N__19115\,
            in2 => \N__19144\,
            in3 => \N__19755\,
            lcout => read_buf_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41130\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i2_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__19505\,
            in1 => \N__19576\,
            in2 => \N__19216\,
            in3 => \N__19751\,
            lcout => read_buf_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41130\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i11_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__19270\,
            in1 => \N__19472\,
            in2 => \N__21096\,
            in3 => \N__22128\,
            lcout => \buf_readRTD_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41130\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.bit_cnt_3771__i3_LC_3_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__20596\,
            in1 => \N__20566\,
            in2 => \N__20517\,
            in3 => \N__20620\,
            lcout => \RTD.bit_cnt_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41132\,
            ce => \N__19389\,
            sr => \N__19812\
        );

    \RTD.i1_4_lut_4_lut_adj_22_LC_3_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000010000000"
        )
    port map (
            in0 => \N__22246\,
            in1 => \N__22115\,
            in2 => \N__22402\,
            in3 => \N__20963\,
            lcout => n11700,
            ltout => \n11700_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i14_LC_3_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__22116\,
            in1 => \N__23415\,
            in2 => \N__19246\,
            in3 => \N__19239\,
            lcout => \buf_readRTD_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41115\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i15_LC_3_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__22117\,
            in1 => \N__19225\,
            in2 => \N__22452\,
            in3 => \N__19430\,
            lcout => \buf_readRTD_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41115\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i15_LC_3_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__19224\,
            in1 => \N__19749\,
            in2 => \N__19243\,
            in3 => \N__19568\,
            lcout => read_buf_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41115\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i1_LC_3_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__22093\,
            in1 => \N__19432\,
            in2 => \N__35325\,
            in3 => \N__19209\,
            lcout => \buf_readRTD_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41141\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i9_LC_3_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__19575\,
            in1 => \N__19618\,
            in2 => \N__19758\,
            in3 => \N__19355\,
            lcout => read_buf_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41141\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i10_LC_3_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__19359\,
            in1 => \N__19745\,
            in2 => \N__19291\,
            in3 => \N__19574\,
            lcout => read_buf_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41141\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i13_LC_3_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__19431\,
            in1 => \N__19378\,
            in2 => \N__22518\,
            in3 => \N__22095\,
            lcout => \buf_readRTD_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41141\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i9_LC_3_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__22094\,
            in1 => \N__19433\,
            in2 => \N__19360\,
            in3 => \N__23646\,
            lcout => \buf_readRTD_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41141\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adress_i1_LC_3_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__19344\,
            in1 => \N__19966\,
            in2 => \N__19651\,
            in3 => \N__19888\,
            lcout => adress_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41133\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adress_i2_LC_3_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__19889\,
            in1 => \N__19345\,
            in2 => \N__19652\,
            in3 => \N__19335\,
            lcout => adress_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41133\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adress_i3_LC_3_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__19336\,
            in1 => \N__19640\,
            in2 => \N__19327\,
            in3 => \N__19890\,
            lcout => adress_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41133\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adress_i4_LC_3_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__19891\,
            in1 => \N__19314\,
            in2 => \N__19653\,
            in3 => \N__19326\,
            lcout => adress_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41133\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adress_i5_LC_3_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__19315\,
            in1 => \N__19641\,
            in2 => \N__19303\,
            in3 => \N__19892\,
            lcout => adress_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41133\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adress_i6_LC_3_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__19893\,
            in1 => \N__19992\,
            in2 => \N__19654\,
            in3 => \N__19302\,
            lcout => adress_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41133\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i10_LC_3_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__19290\,
            in1 => \N__19457\,
            in2 => \N__23391\,
            in3 => \N__22127\,
            lcout => \buf_readRTD_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41133\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i12069_2_lut_LC_3_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__22260\,
            in1 => \N__22404\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n14465,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i8_LC_3_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__22123\,
            in1 => \N__21813\,
            in2 => \N__19474\,
            in3 => \N__19617\,
            lcout => \buf_readRTD_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41129\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i2_LC_3_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__19506\,
            in1 => \N__19466\,
            in2 => \N__33261\,
            in3 => \N__22124\,
            lcout => \buf_readRTD_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41129\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i4_LC_3_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__19595\,
            in1 => \N__19579\,
            in2 => \N__19492\,
            in3 => \N__19750\,
            lcout => read_buf_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41129\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i4_LC_3_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__19596\,
            in1 => \N__19468\,
            in2 => \N__33207\,
            in3 => \N__22126\,
            lcout => \buf_readRTD_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41129\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.read_buf_i3_LC_3_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__19487\,
            in1 => \N__19578\,
            in2 => \N__19759\,
            in3 => \N__19507\,
            lcout => read_buf_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41129\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.READ_DATA_i3_LC_3_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__19491\,
            in1 => \N__19467\,
            in2 => \N__33558\,
            in3 => \N__22125\,
            lcout => \buf_readRTD_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41129\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.bit_cnt_3771__i1_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20588\,
            in2 => \_gnd_net_\,
            in3 => \N__20615\,
            lcout => \RTD.bit_cnt_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41083\,
            ce => \N__19396\,
            sr => \N__19816\
        );

    \RTD.bit_cnt_3771__i0_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20587\,
            lcout => \RTD.bit_cnt_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41083\,
            ce => \N__19396\,
            sr => \N__19816\
        );

    \RTD.bit_cnt_3771__i2_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__20616\,
            in1 => \_gnd_net_\,
            in2 => \N__20595\,
            in3 => \N__20562\,
            lcout => \RTD.bit_cnt_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41083\,
            ce => \N__19396\,
            sr => \N__19816\
        );

    \RTD.MOSI_59_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__20927\,
            in1 => \N__19981\,
            in2 => \N__21004\,
            in3 => \N__22101\,
            lcout => \RTD_SDI\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41142\,
            ce => \N__19777\,
            sr => \N__19953\
        );

    \RTD.i1_3_lut_4_lut_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__22220\,
            in1 => \N__20544\,
            in2 => \N__20524\,
            in3 => \N__20925\,
            lcout => \RTD.n33\,
            ltout => \RTD.n33_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i24_3_lut_4_lut_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001000100"
        )
    port map (
            in0 => \N__20926\,
            in1 => \N__22221\,
            in2 => \N__19762\,
            in3 => \N__22100\,
            lcout => \RTD.n11_adj_1394\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i2_3_lut_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__20923\,
            in1 => \N__22353\,
            in2 => \_gnd_net_\,
            in3 => \N__22099\,
            lcout => n1_adj_1575,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_2_lut_adj_20_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22219\,
            in2 => \_gnd_net_\,
            in3 => \N__20924\,
            lcout => \RTD.n4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i31_3_lut_4_lut_3_lut_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__20894\,
            in1 => \N__22323\,
            in2 => \_gnd_net_\,
            in3 => \N__22191\,
            lcout => \RTD.n14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_2_lut_adj_24_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19928\,
            in2 => \_gnd_net_\,
            in3 => \N__20144\,
            lcout => \RTD.n16614\,
            ltout => \RTD.n16614_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i2_3_lut_adj_19_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110101"
        )
    port map (
            in0 => \N__20895\,
            in1 => \_gnd_net_\,
            in2 => \N__19657\,
            in3 => \N__21903\,
            lcout => \RTD.n11712\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_2_lut_adj_26_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__22324\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19859\,
            lcout => \RTD.n19855\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i19027_3_lut_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111111"
        )
    port map (
            in0 => \N__20896\,
            in1 => \N__20102\,
            in2 => \_gnd_net_\,
            in3 => \N__19843\,
            lcout => \RTD.n21091\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i16891_3_lut_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__22192\,
            in1 => \N__20518\,
            in2 => \_gnd_net_\,
            in3 => \N__20540\,
            lcout => \RTD.n19482\,
            ltout => \RTD.n19482_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adc_state_3__I_0_66_Mux_0_i7_4_lut_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010111010101"
        )
    port map (
            in0 => \N__20897\,
            in1 => \N__20103\,
            in2 => \N__19837\,
            in3 => \N__22030\,
            lcout => \RTD.n7_adj_1395\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_2_lut_3_lut_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__22190\,
            in1 => \N__21983\,
            in2 => \_gnd_net_\,
            in3 => \N__20893\,
            lcout => \RTD.n1_adj_1393\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i18129_2_lut_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22193\,
            in2 => \_gnd_net_\,
            in3 => \N__21989\,
            lcout => \RTD.n7285\,
            ltout => \RTD.n7285_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_4_lut_adj_13_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__20914\,
            in1 => \N__19929\,
            in2 => \N__19834\,
            in3 => \N__20142\,
            lcout => OPEN,
            ltout => \RTD.n21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_4_lut_adj_14_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011001000"
        )
    port map (
            in0 => \N__22350\,
            in1 => \N__20098\,
            in2 => \N__19831\,
            in3 => \N__21990\,
            lcout => \RTD.n16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i18734_4_lut_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101000"
        )
    port map (
            in0 => \N__19828\,
            in1 => \N__22351\,
            in2 => \N__20104\,
            in3 => \N__20005\,
            lcout => OPEN,
            ltout => \RTD.n20969_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adc_state_i2_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__22352\,
            in1 => \N__20475\,
            in2 => \N__19819\,
            in3 => \N__21991\,
            lcout => adc_state_2_adj_1474,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41134\,
            ce => \N__20683\,
            sr => \_gnd_net_\
        );

    \RTD.i1_2_lut_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__20519\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20545\,
            lcout => \RTD.n32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i4916_2_lut_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22194\,
            in2 => \_gnd_net_\,
            in3 => \N__20913\,
            lcout => \RTD.n1_adj_1392\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adress_i7_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011000000"
        )
    port map (
            in0 => \N__20143\,
            in1 => \N__19999\,
            in2 => \N__22261\,
            in3 => \N__20944\,
            lcout => \RTD.adress_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41082\,
            ce => \N__19894\,
            sr => \N__19957\
        );

    \RTD.adress_i0_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110001011111"
        )
    port map (
            in0 => \N__20943\,
            in1 => \N__19980\,
            in2 => \N__20149\,
            in3 => \N__22248\,
            lcout => adress_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41082\,
            ce => \N__19894\,
            sr => \N__19957\
        );

    \RTD.i7_4_lut_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__20077\,
            in1 => \N__21202\,
            in2 => \N__20044\,
            in3 => \N__20797\,
            lcout => \RTD.adress_7_N_1331_7\,
            ltout => \RTD.adress_7_N_1331_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_2_lut_adj_16_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110101"
        )
    port map (
            in0 => \N__20941\,
            in1 => \_gnd_net_\,
            in2 => \N__19936\,
            in3 => \_gnd_net_\,
            lcout => \RTD.n11\,
            ltout => \RTD.n11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i34_4_lut_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101101010001"
        )
    port map (
            in0 => \N__22247\,
            in1 => \N__19933\,
            in2 => \N__19900\,
            in3 => \N__20942\,
            lcout => OPEN,
            ltout => \RTD.n19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i35_4_lut_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011000"
        )
    port map (
            in0 => \N__22361\,
            in1 => \N__19863\,
            in2 => \N__19897\,
            in3 => \N__22026\,
            lcout => n13151,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i22_4_lut_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111000000"
        )
    port map (
            in0 => \N__20730\,
            in1 => \N__22360\,
            in2 => \N__19864\,
            in3 => \N__20790\,
            lcout => n13162,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.mode_53_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100001000"
        )
    port map (
            in0 => \N__20965\,
            in1 => \N__20145\,
            in2 => \N__21910\,
            in3 => \N__20113\,
            lcout => \RTD.mode\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41116\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i2_4_lut_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__23819\,
            in1 => \N__20061\,
            in2 => \N__42075\,
            in3 => \N__20070\,
            lcout => \RTD.n10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i2_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__20071\,
            in1 => \N__21155\,
            in2 => \N__23823\,
            in3 => \N__21184\,
            lcout => \RTD.cfg_buf_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41116\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i4_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__21185\,
            in1 => \N__20062\,
            in2 => \N__42074\,
            in3 => \N__21157\,
            lcout => \RTD.cfg_buf_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41116\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i7_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__20053\,
            in1 => \N__21156\,
            in2 => \N__24194\,
            in3 => \N__21187\,
            lcout => \RTD.cfg_buf_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41116\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i4_4_lut_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__23697\,
            in1 => \N__20052\,
            in2 => \N__24195\,
            in3 => \N__20034\,
            lcout => \RTD.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i1_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__20035\,
            in1 => \N__21154\,
            in2 => \N__23698\,
            in3 => \N__21183\,
            lcout => cfg_buf_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41116\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i5_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__21186\,
            in1 => \N__21214\,
            in2 => \N__41436\,
            in3 => \N__21158\,
            lcout => \RTD.cfg_buf_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41116\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_7_i19_3_lut_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23581\,
            in1 => \N__20189\,
            in2 => \_gnd_net_\,
            in3 => \N__56901\,
            lcout => OPEN,
            ltout => \n19_adj_1622_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19365_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011001100"
        )
    port map (
            in0 => \N__20026\,
            in1 => \N__57503\,
            in2 => \N__20200\,
            in3 => \N__47737\,
            lcout => n21961,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i15_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__48315\,
            in1 => \N__20190\,
            in2 => \N__48533\,
            in3 => \N__21238\,
            lcout => buf_adcdata_vac_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55174\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_3_i30_3_lut_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20176\,
            in1 => \N__21022\,
            in2 => \_gnd_net_\,
            in3 => \N__56347\,
            lcout => n30_adj_1612,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i3_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__50908\,
            in1 => \N__48999\,
            in2 => \N__49041\,
            in3 => \N__21042\,
            lcout => buf_adcdata_iac_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55174\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18784_2_lut_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20164\,
            in2 => \_gnd_net_\,
            in3 => \N__56902\,
            lcout => n20937,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i2_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__50907\,
            in1 => \N__48998\,
            in2 => \N__21322\,
            in3 => \N__22490\,
            lcout => buf_adcdata_iac_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55174\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i18_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__48505\,
            in1 => \N__48321\,
            in2 => \N__21298\,
            in3 => \N__23852\,
            lcout => buf_adcdata_vac_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55190\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i21_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__48506\,
            in1 => \N__48322\,
            in2 => \N__21346\,
            in3 => \N__21839\,
            lcout => buf_adcdata_vac_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55190\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i9_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__21251\,
            in1 => \N__50935\,
            in2 => \N__21447\,
            in3 => \N__50516\,
            lcout => cmd_rdadctmp_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55190\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i11_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__49025\,
            in1 => \N__50934\,
            in2 => \N__21321\,
            in3 => \N__50515\,
            lcout => cmd_rdadctmp_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55190\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19423_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__56904\,
            in1 => \N__24690\,
            in2 => \N__57538\,
            in3 => \N__27873\,
            lcout => n22039,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i29_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__37878\,
            in1 => \N__21338\,
            in2 => \N__20305\,
            in3 => \N__48286\,
            lcout => cmd_rdadctmp_29_adj_1414,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55204\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i28_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__48285\,
            in1 => \N__20300\,
            in2 => \N__21276\,
            in3 => \N__37877\,
            lcout => cmd_rdadctmp_28_adj_1415,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55204\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i20_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__48284\,
            in1 => \N__48492\,
            in2 => \N__25706\,
            in3 => \N__20304\,
            lcout => buf_adcdata_vac_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55204\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i7_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__22818\,
            in1 => \N__48287\,
            in2 => \N__21583\,
            in3 => \N__37872\,
            lcout => cmd_rdadctmp_7_adj_1436,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55216\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19516_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__21403\,
            in1 => \N__57446\,
            in2 => \N__20290\,
            in3 => \N__47823\,
            lcout => n22117,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_199_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000110"
        )
    port map (
            in0 => \N__48203\,
            in1 => \N__29855\,
            in2 => \N__20244\,
            in3 => \N__29782\,
            lcout => n14_adj_1577,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_104_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29854\,
            in2 => \_gnd_net_\,
            in3 => \N__29781\,
            lcout => n20573,
            ltout => \n20573_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.CS_37_LC_5_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100100011"
        )
    port map (
            in0 => \N__22982\,
            in1 => \N__20263\,
            in2 => \N__20257\,
            in3 => \N__48205\,
            lcout => \VAC_CS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55227\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.SCLK_35_LC_5_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000011100100"
        )
    port map (
            in0 => \N__48204\,
            in1 => \N__29856\,
            in2 => \N__20217\,
            in3 => \N__29783\,
            lcout => \VAC_SCLK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55227\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i12_LC_5_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__48961\,
            in1 => \N__50954\,
            in2 => \N__21801\,
            in3 => \N__33462\,
            lcout => buf_adcdata_iac_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55237\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i22_LC_5_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__50493\,
            in1 => \N__21777\,
            in2 => \N__50965\,
            in3 => \N__24446\,
            lcout => cmd_rdadctmp_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55237\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i20_LC_5_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__21794\,
            in1 => \N__50956\,
            in2 => \N__21759\,
            in3 => \N__50494\,
            lcout => cmd_rdadctmp_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55237\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i14_LC_5_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__48962\,
            in1 => \N__50955\,
            in2 => \N__24453\,
            in3 => \N__29576\,
            lcout => buf_adcdata_iac_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55237\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i13_LC_5_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__50880\,
            in1 => \N__48967\,
            in2 => \N__21781\,
            in3 => \N__25808\,
            lcout => buf_adcdata_iac_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55240\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18773_2_lut_LC_5_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__56911\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20407\,
            lcout => n21001,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i11_LC_5_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__48966\,
            in1 => \N__50881\,
            in2 => \N__21760\,
            in3 => \N__33534\,
            lcout => buf_adcdata_iac_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55240\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_354_Mux_7_i15_4_lut_LC_5_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__54723\,
            in1 => \N__30079\,
            in2 => \N__52192\,
            in3 => \N__42435\,
            lcout => \data_index_9_N_212_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.bit_cnt_i3_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111100011110000"
        )
    port map (
            in0 => \N__20430\,
            in1 => \N__23232\,
            in2 => \N__23209\,
            in3 => \N__20453\,
            lcout => bit_cnt_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55082\,
            ce => \N__28907\,
            sr => \N__20740\
        );

    \CLK_DDS.bit_cnt_i2_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__23231\,
            in1 => \_gnd_net_\,
            in2 => \N__20457\,
            in3 => \N__20429\,
            lcout => bit_cnt_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55082\,
            ce => \N__28907\,
            sr => \N__20740\
        );

    \CLK_DDS.bit_cnt_i1_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20449\,
            in2 => \_gnd_net_\,
            in3 => \N__23230\,
            lcout => bit_cnt_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55082\,
            ce => \N__28907\,
            sr => \N__20740\
        );

    \CLK_DDS.dds_state_i0_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100010100000101"
        )
    port map (
            in0 => \N__28612\,
            in1 => \N__20413\,
            in2 => \N__28908\,
            in3 => \N__23191\,
            lcout => dds_state_0_adj_1447,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55087\,
            ce => \N__20640\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.i19109_4_lut_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011110"
        )
    port map (
            in0 => \N__28593\,
            in1 => \N__28865\,
            in2 => \N__28678\,
            in3 => \N__28746\,
            lcout => \CLK_DDS.n9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.dds_state_i1_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__28749\,
            in1 => \N__28594\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => dds_state_1_adj_1446,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55095\,
            ce => \N__20641\,
            sr => \N__28973\
        );

    \RTD.i2_3_lut_adj_18_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__20614\,
            in1 => \N__20586\,
            in2 => \_gnd_net_\,
            in3 => \N__20561\,
            lcout => \RTD.n17638\,
            ltout => \RTD.n17638_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i19033_3_lut_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20520\,
            in2 => \N__20482\,
            in3 => \N__22222\,
            lcout => OPEN,
            ltout => \RTD.n21063_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adc_state_3__I_0_66_Mux_0_i14_4_lut_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100010001000"
        )
    port map (
            in0 => \N__20479\,
            in1 => \N__22102\,
            in2 => \N__20461\,
            in3 => \N__20928\,
            lcout => \RTD.n17676\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.i3_3_lut_4_lut_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__28748\,
            in1 => \N__28591\,
            in2 => \N__20458\,
            in3 => \N__20431\,
            lcout => n8_adj_1409,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.i1_3_lut_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001000100"
        )
    port map (
            in0 => \N__28592\,
            in1 => \N__28866\,
            in2 => \_gnd_net_\,
            in3 => \N__28747\,
            lcout => \CLK_DDS.n16711\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.adc_state_i1_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101010000"
        )
    port map (
            in0 => \N__22387\,
            in1 => \N__20731\,
            in2 => \N__20719\,
            in3 => \N__20940\,
            lcout => \RTD.adc_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41099\,
            ce => \N__20679\,
            sr => \_gnd_net_\
        );

    \RTD.adc_state_i3_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010110111011"
        )
    port map (
            in0 => \N__22354\,
            in1 => \N__20710\,
            in2 => \N__20704\,
            in3 => \N__22104\,
            lcout => \RTD.adc_state_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41099\,
            ce => \N__20679\,
            sr => \_gnd_net_\
        );

    \RTD.adc_state_i0_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__22388\,
            in1 => \N__20695\,
            in2 => \_gnd_net_\,
            in3 => \N__20689\,
            lcout => \RTD.adc_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41099\,
            ce => \N__20679\,
            sr => \_gnd_net_\
        );

    \RTD.cfg_tmp_i1_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101011000000"
        )
    port map (
            in0 => \N__20932\,
            in1 => \N__20983\,
            in2 => \N__22130\,
            in3 => \N__23682\,
            lcout => \RTD.cfg_tmp_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41098\,
            ce => \N__20767\,
            sr => \N__20752\
        );

    \RTD.cfg_tmp_i2_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010010100000"
        )
    port map (
            in0 => \N__22032\,
            in1 => \N__23827\,
            in2 => \N__20668\,
            in3 => \N__20937\,
            lcout => \RTD.cfg_tmp_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41098\,
            ce => \N__20767\,
            sr => \N__20752\
        );

    \RTD.cfg_tmp_i3_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010100000"
        )
    port map (
            in0 => \N__20933\,
            in1 => \N__20659\,
            in2 => \N__23785\,
            in3 => \N__22036\,
            lcout => \RTD.cfg_tmp_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41098\,
            ce => \N__20767\,
            sr => \N__20752\
        );

    \RTD.cfg_tmp_i4_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100010001000"
        )
    port map (
            in0 => \N__22033\,
            in1 => \N__20653\,
            in2 => \N__42076\,
            in3 => \N__20938\,
            lcout => \RTD.cfg_tmp_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41098\,
            ce => \N__20767\,
            sr => \N__20752\
        );

    \RTD.cfg_tmp_i5_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110000100000"
        )
    port map (
            in0 => \N__20934\,
            in1 => \N__22035\,
            in2 => \N__41437\,
            in3 => \N__20647\,
            lcout => \RTD.cfg_tmp_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41098\,
            ce => \N__20767\,
            sr => \N__20752\
        );

    \RTD.cfg_tmp_i6_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100010001000"
        )
    port map (
            in0 => \N__22034\,
            in1 => \N__21016\,
            in2 => \N__29329\,
            in3 => \N__20939\,
            lcout => \RTD.cfg_tmp_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41098\,
            ce => \N__20767\,
            sr => \N__20752\
        );

    \RTD.cfg_tmp_i7_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010100000"
        )
    port map (
            in0 => \N__20935\,
            in1 => \N__21010\,
            in2 => \N__24199\,
            in3 => \N__22037\,
            lcout => \RTD.cfg_tmp_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41098\,
            ce => \N__20767\,
            sr => \N__20752\
        );

    \RTD.cfg_tmp_i0_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100010001000"
        )
    port map (
            in0 => \N__22031\,
            in1 => \N__20994\,
            in2 => \N__23737\,
            in3 => \N__20936\,
            lcout => \RTD.cfg_tmp_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41098\,
            ce => \N__20767\,
            sr => \N__20752\
        );

    \RTD.i1_3_lut_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011111111"
        )
    port map (
            in0 => \N__20945\,
            in1 => \_gnd_net_\,
            in2 => \N__22389\,
            in3 => \N__21152\,
            lcout => n18586,
            ltout => \n18586_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i0_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010100000"
        )
    port map (
            in0 => \N__20806\,
            in1 => \N__23732\,
            in2 => \N__20809\,
            in3 => \N__21153\,
            lcout => cfg_buf_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41079\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i1_4_lut_adj_23_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__23733\,
            in1 => \N__21114\,
            in2 => \N__29325\,
            in3 => \N__20805\,
            lcout => \RTD.n9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i18127_2_lut_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__22223\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22355\,
            lcout => OPEN,
            ltout => \RTD.n20722_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i30_4_lut_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000001010"
        )
    port map (
            in0 => \N__20791\,
            in1 => \N__20779\,
            in2 => \N__20770\,
            in3 => \N__22025\,
            lcout => \RTD.n13198\,
            ltout => \RTD.n13198_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i12587_2_lut_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__20755\,
            in3 => \N__22359\,
            lcout => \RTD.n14984\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i3_4_lut_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111111110110"
        )
    port map (
            in0 => \N__41426\,
            in1 => \N__21213\,
            in2 => \N__23777\,
            in3 => \N__21195\,
            lcout => \RTD.n11_adj_1396\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i3_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__21196\,
            in1 => \N__21159\,
            in2 => \N__23778\,
            in3 => \N__21181\,
            lcout => \RTD.cfg_buf_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41097\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.cfg_buf_i6_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__21182\,
            in1 => \N__21115\,
            in2 => \N__29318\,
            in3 => \N__21160\,
            lcout => \RTD.cfg_buf_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__41097\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19496_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__23767\,
            in1 => \N__57310\,
            in2 => \N__21103\,
            in3 => \N__56903\,
            lcout => OPEN,
            ltout => \n22099_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22099_bdd_4_lut_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__57311\,
            in1 => \N__21065\,
            in2 => \N__21079\,
            in3 => \N__23290\,
            lcout => OPEN,
            ltout => \n22102_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18255_3_lut_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__47820\,
            in1 => \N__29524\,
            in2 => \N__21076\,
            in3 => \_gnd_net_\,
            lcout => n20850,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i19_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__48319\,
            in1 => \N__48495\,
            in2 => \N__21277\,
            in3 => \N__21069\,
            lcout => buf_adcdata_vac_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55146\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_3_i19_3_lut_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23179\,
            in1 => \N__21474\,
            in2 => \_gnd_net_\,
            in3 => \N__56905\,
            lcout => OPEN,
            ltout => \n19_adj_1610_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_3_i22_3_lut_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47741\,
            in2 => \N__21049\,
            in3 => \N__21038\,
            lcout => n22_adj_1611,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i0_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__50906\,
            in1 => \N__48997\,
            in2 => \N__21451\,
            in3 => \N__23450\,
            lcout => buf_adcdata_iac_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55146\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i21_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__21557\,
            in1 => \N__48320\,
            in2 => \N__24142\,
            in3 => \N__37870\,
            lcout => cmd_rdadctmp_21_adj_1422,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55146\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i26_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__37874\,
            in1 => \N__24235\,
            in2 => \N__48346\,
            in3 => \N__21290\,
            lcout => cmd_rdadctmp_26_adj_1417,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55161\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i30_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__22619\,
            in1 => \N__48325\,
            in2 => \N__21345\,
            in3 => \N__37876\,
            lcout => cmd_rdadctmp_30_adj_1413,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55161\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i10_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__21314\,
            in1 => \N__21252\,
            in2 => \N__50910\,
            in3 => \N__50514\,
            lcout => cmd_rdadctmp_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55161\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i24_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__24251\,
            in1 => \N__48323\,
            in2 => \N__21237\,
            in3 => \N__37873\,
            lcout => cmd_rdadctmp_24_adj_1419,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55161\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i27_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__21269\,
            in1 => \N__48324\,
            in2 => \N__21297\,
            in3 => \N__37875\,
            lcout => cmd_rdadctmp_27_adj_1416,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55161\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i1_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__48990\,
            in1 => \N__50936\,
            in2 => \N__23627\,
            in3 => \N__21253\,
            lcout => buf_adcdata_iac_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55161\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i23_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__48196\,
            in1 => \N__21230\,
            in2 => \N__21420\,
            in3 => \N__37840\,
            lcout => cmd_rdadctmp_23_adj_1420,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55176\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18241_3_lut_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__21672\,
            in1 => \N__24268\,
            in2 => \_gnd_net_\,
            in3 => \N__57485\,
            lcout => n20836,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i11_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__48195\,
            in1 => \N__22838\,
            in2 => \N__22566\,
            in3 => \N__37838\,
            lcout => cmd_rdadctmp_11_adj_1432,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55176\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i3_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__48493\,
            in1 => \N__48197\,
            in2 => \N__22845\,
            in3 => \N__21473\,
            lcout => buf_adcdata_vac_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55176\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i14_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__48194\,
            in1 => \N__48494\,
            in2 => \N__21421\,
            in3 => \N__22677\,
            lcout => buf_adcdata_vac_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55176\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i8_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__24286\,
            in1 => \N__50953\,
            in2 => \N__21446\,
            in3 => \N__50513\,
            lcout => cmd_rdadctmp_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55176\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i22_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__37839\,
            in1 => \N__21413\,
            in2 => \N__21568\,
            in3 => \N__48198\,
            lcout => cmd_rdadctmp_22_adj_1421,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55176\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i8_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__48439\,
            in1 => \N__21387\,
            in2 => \N__48265\,
            in3 => \N__22726\,
            lcout => buf_adcdata_vac_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55191\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_5_i19_3_lut_LC_6_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__21533\,
            in1 => \N__23350\,
            in2 => \_gnd_net_\,
            in3 => \N__56907\,
            lcout => n19_adj_1487,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_0_i19_3_lut_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__56908\,
            in1 => \N__26635\,
            in2 => \_gnd_net_\,
            in3 => \N__21386\,
            lcout => OPEN,
            ltout => \n19_adj_1479_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19393_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010101010"
        )
    port map (
            in0 => \N__57448\,
            in1 => \N__21373\,
            in2 => \N__21349\,
            in3 => \N__47821\,
            lcout => n21973,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_6_i23_3_lut_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__55962\,
            in1 => \N__56906\,
            in2 => \_gnd_net_\,
            in3 => \N__36664\,
            lcout => OPEN,
            ltout => \n23_adj_1512_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18247_4_lut_LC_6_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__56909\,
            in1 => \N__57449\,
            in2 => \N__21586\,
            in3 => \N__45235\,
            lcout => n20842,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i4_LC_6_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__21513\,
            in1 => \N__48113\,
            in2 => \N__22879\,
            in3 => \N__37785\,
            lcout => cmd_rdadctmp_4_adj_1439,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55205\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i6_LC_6_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__37787\,
            in1 => \N__21579\,
            in2 => \N__48202\,
            in3 => \N__21502\,
            lcout => cmd_rdadctmp_6_adj_1437,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55205\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i13_LC_6_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__48437\,
            in1 => \N__48112\,
            in2 => \N__21541\,
            in3 => \N__21567\,
            lcout => buf_adcdata_vac_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55205\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i5_LC_6_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__37786\,
            in1 => \N__21501\,
            in2 => \N__21517\,
            in3 => \N__48117\,
            lcout => cmd_rdadctmp_5_adj_1438,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55205\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19061_2_lut_LC_6_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21493\,
            in2 => \_gnd_net_\,
            in3 => \N__56910\,
            lcout => n21109,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i18_LC_6_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__50491\,
            in1 => \N__21696\,
            in2 => \N__50909\,
            in3 => \N__21725\,
            lcout => cmd_rdadctmp_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55205\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i17_LC_6_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__21695\,
            in1 => \N__50830\,
            in2 => \N__45139\,
            in3 => \N__50492\,
            lcout => cmd_rdadctmp_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55205\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i21_LC_6_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__21776\,
            in1 => \N__50856\,
            in2 => \N__21802\,
            in3 => \N__50496\,
            lcout => cmd_rdadctmp_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55217\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i19_LC_6_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__21752\,
            in1 => \N__50855\,
            in2 => \N__21732\,
            in3 => \N__50495\,
            lcout => cmd_rdadctmp_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55217\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i10_LC_6_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__48892\,
            in1 => \N__50960\,
            in2 => \N__21736\,
            in3 => \N__25961\,
            lcout => buf_adcdata_iac_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55228\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18806_2_lut_LC_6_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21709\,
            in2 => \_gnd_net_\,
            in3 => \N__56912\,
            lcout => n21285,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i9_LC_6_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__48873\,
            in1 => \N__50821\,
            in2 => \N__21700\,
            in3 => \N__21671\,
            lcout => buf_adcdata_iac_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55238\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pll_main.i19651_1_lut_LC_7_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56040\,
            lcout => \DDS_MCLK1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.bit_cnt_i0_LC_7_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111101000000"
        )
    port map (
            in0 => \N__28776\,
            in1 => \N__28607\,
            in2 => \N__28942\,
            in3 => \N__23233\,
            lcout => bit_cnt_0_adj_1449,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55076\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.CS_28_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001110111"
        )
    port map (
            in0 => \N__28876\,
            in1 => \N__28773\,
            in2 => \_gnd_net_\,
            in3 => \N__28613\,
            lcout => \DDS_CS1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55083\,
            ce => \N__23269\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.SCLK_27_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010011010001"
        )
    port map (
            in0 => \N__28750\,
            in1 => \N__28617\,
            in2 => \N__21603\,
            in3 => \N__28880\,
            lcout => \DDS_SCK1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55096\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RTD.i2_2_lut_3_lut_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__22333\,
            in1 => \N__22195\,
            in2 => \_gnd_net_\,
            in3 => \N__22103\,
            lcout => \RTD.n20487\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.dds_state_i2_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28941\,
            in2 => \_gnd_net_\,
            in3 => \N__28736\,
            lcout => dds_state_2_adj_1445,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55113\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18248_4_lut_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010001000"
        )
    port map (
            in0 => \N__21889\,
            in1 => \N__57187\,
            in2 => \N__31339\,
            in3 => \N__56982\,
            lcout => n20843,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.MOSI_31_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__28940\,
            in1 => \N__27726\,
            in2 => \_gnd_net_\,
            in3 => \N__21867\,
            lcout => \DDS_MOSI1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55113\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i1_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__45331\,
            in1 => \N__52195\,
            in2 => \N__44146\,
            in3 => \N__23681\,
            lcout => \buf_cfgRTD_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55113\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_217_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__41365\,
            in1 => \N__51298\,
            in2 => \_gnd_net_\,
            in3 => \N__54093\,
            lcout => n14_adj_1516,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22141_bdd_4_lut_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100010"
        )
    port map (
            in0 => \N__22704\,
            in1 => \N__23404\,
            in2 => \N__23542\,
            in3 => \N__57191\,
            lcout => n20828,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22153_bdd_4_lut_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100010"
        )
    port map (
            in0 => \N__21852\,
            in1 => \N__22501\,
            in2 => \N__23374\,
            in3 => \N__57188\,
            lcout => n22156,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19541_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__56886\,
            in1 => \N__23717\,
            in2 => \N__21823\,
            in3 => \N__57192\,
            lcout => OPEN,
            ltout => \n22183_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22183_bdd_4_lut_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__23326\,
            in1 => \N__22596\,
            in2 => \N__22543\,
            in3 => \N__57190\,
            lcout => n20772,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22165_bdd_4_lut_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100010"
        )
    port map (
            in0 => \N__22652\,
            in1 => \N__23635\,
            in2 => \N__23524\,
            in3 => \N__57189\,
            lcout => n20814,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_2_i30_3_lut_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__22465\,
            in1 => \_gnd_net_\,
            in2 => \N__22540\,
            in3 => \N__56271\,
            lcout => n30_adj_1615,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19521_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__41425\,
            in1 => \N__57182\,
            in2 => \N__22525\,
            in3 => \N__56865\,
            lcout => n22153,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i0_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__48524\,
            in1 => \N__48179\,
            in2 => \N__22807\,
            in3 => \N__23477\,
            lcout => buf_adcdata_vac_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55134\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_2_i19_3_lut_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23308\,
            in1 => \N__22424\,
            in2 => \_gnd_net_\,
            in3 => \N__56867\,
            lcout => OPEN,
            ltout => \n19_adj_1613_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_2_i22_3_lut_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__22491\,
            in1 => \_gnd_net_\,
            in2 => \N__22468\,
            in3 => \N__47742\,
            lcout => n22_adj_1614,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19501_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__56866\,
            in1 => \N__24175\,
            in2 => \N__22459\,
            in3 => \N__57181\,
            lcout => n22135,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i2_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__48178\,
            in1 => \N__48525\,
            in2 => \N__22570\,
            in3 => \N__22425\,
            lcout => buf_adcdata_vac_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55134\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i22_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__48508\,
            in1 => \N__48176\,
            in2 => \N__22627\,
            in3 => \N__22703\,
            lcout => buf_adcdata_vac_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55147\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_6_i19_3_lut_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__56883\,
            in1 => \N__23560\,
            in2 => \_gnd_net_\,
            in3 => \N__22673\,
            lcout => n19_adj_1482,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i17_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__48173\,
            in1 => \N__48509\,
            in2 => \N__22656\,
            in3 => \N__24234\,
            lcout => buf_adcdata_vac_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55147\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i31_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__22605\,
            in1 => \N__48177\,
            in2 => \N__22626\,
            in3 => \N__37844\,
            lcout => cmd_rdadctmp_31_adj_1412,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55147\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i23_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__48174\,
            in1 => \N__48510\,
            in2 => \N__24338\,
            in3 => \N__22606\,
            lcout => buf_adcdata_vac_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55147\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i16_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__48507\,
            in1 => \N__48175\,
            in2 => \N__22597\,
            in3 => \N__24255\,
            lcout => buf_adcdata_vac_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55147\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i18_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__37834\,
            in1 => \N__22740\,
            in2 => \N__48262\,
            in3 => \N__24110\,
            lcout => cmd_rdadctmp_18_adj_1425,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55162\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i1_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__48478\,
            in1 => \N__48181\,
            in2 => \N__22783\,
            in3 => \N__23960\,
            lcout => buf_adcdata_vac_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55162\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i9_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__48180\,
            in1 => \N__48479\,
            in2 => \N__35276\,
            in3 => \N__22741\,
            lcout => buf_adcdata_vac_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55162\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i10_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__22559\,
            in1 => \N__48182\,
            in2 => \N__22782\,
            in3 => \N__37832\,
            lcout => cmd_rdadctmp_10_adj_1433,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55162\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i19_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__37835\,
            in1 => \N__24111\,
            in2 => \N__48263\,
            in3 => \N__24020\,
            lcout => cmd_rdadctmp_19_adj_1424,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55162\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i12_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__47948\,
            in1 => \N__48183\,
            in2 => \N__22846\,
            in3 => \N__37833\,
            lcout => cmd_rdadctmp_12_adj_1431,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55162\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i8_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__37836\,
            in1 => \N__22796\,
            in2 => \N__48264\,
            in3 => \N__22825\,
            lcout => cmd_rdadctmp_8_adj_1435,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55162\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i9_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__22775\,
            in1 => \N__48184\,
            in2 => \N__22803\,
            in3 => \N__37837\,
            lcout => cmd_rdadctmp_9_adj_1434,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55162\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i0_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__22905\,
            in1 => \N__48223\,
            in2 => \N__22765\,
            in3 => \N__37779\,
            lcout => cmd_rdadctmp_0_adj_1443,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55177\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n21973_bdd_4_lut_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100010"
        )
    port map (
            in0 => \N__27838\,
            in1 => \N__22747\,
            in2 => \N__24420\,
            in3 => \N__47822\,
            lcout => n21976,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i17_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__37781\,
            in1 => \N__22725\,
            in2 => \N__48281\,
            in3 => \N__22739\,
            lcout => cmd_rdadctmp_17_adj_1426,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55177\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i16_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__22724\,
            in1 => \N__48224\,
            in2 => \N__45205\,
            in3 => \N__37780\,
            lcout => cmd_rdadctmp_16_adj_1427,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55177\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i2_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__37783\,
            in1 => \N__22897\,
            in2 => \N__48282\,
            in3 => \N__22887\,
            lcout => cmd_rdadctmp_2_adj_1441,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55177\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i1_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__22896\,
            in1 => \N__48225\,
            in2 => \N__22909\,
            in3 => \N__37782\,
            lcout => cmd_rdadctmp_1_adj_1442,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55177\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i3_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__37784\,
            in1 => \N__22888\,
            in2 => \N__48283\,
            in3 => \N__22875\,
            lcout => cmd_rdadctmp_3_adj_1440,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55177\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i1_3_lut_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__48040\,
            in1 => \N__22993\,
            in2 => \_gnd_net_\,
            in3 => \N__22864\,
            lcout => n12643,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.adc_state_i2_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011000100010"
        )
    port map (
            in0 => \N__29766\,
            in1 => \N__29845\,
            in2 => \_gnd_net_\,
            in3 => \N__48042\,
            lcout => \DTRIG_N_910_adj_1444\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55192\,
            ce => \N__22951\,
            sr => \_gnd_net_\
        );

    \ADC_VAC.adc_state_i1_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011110101"
        )
    port map (
            in0 => \N__48041\,
            in1 => \_gnd_net_\,
            in2 => \N__29858\,
            in3 => \N__29767\,
            lcout => adc_state_1_adj_1410,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55192\,
            ce => \N__22951\,
            sr => \_gnd_net_\
        );

    \ADC_VAC.i1_4_lut_adj_4_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000010100"
        )
    port map (
            in0 => \N__48039\,
            in1 => \N__29765\,
            in2 => \N__29857\,
            in3 => \N__22994\,
            lcout => \ADC_VAC.n12556\,
            ltout => \ADC_VAC.n12556_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i12432_2_lut_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22855\,
            in3 => \N__29841\,
            lcout => \ADC_VAC.n14829\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_118_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29764\,
            in2 => \_gnd_net_\,
            in3 => \N__29837\,
            lcout => n20540,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i1_2_lut_adj_3_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__29787\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22852\,
            lcout => \ADC_VAC.n20668\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i1_4_lut_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111101111"
        )
    port map (
            in0 => \N__29846\,
            in1 => \N__48035\,
            in2 => \N__22999\,
            in3 => \N__30141\,
            lcout => \ADC_VAC.n20667\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i18152_4_lut_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23104\,
            in1 => \N__23118\,
            in2 => \N__22927\,
            in3 => \N__23133\,
            lcout => OPEN,
            ltout => \ADC_VAC.n20747_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i18168_4_lut_LC_7_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__23070\,
            in1 => \N__22941\,
            in2 => \N__23017\,
            in3 => \N__23052\,
            lcout => OPEN,
            ltout => \ADC_VAC.n20763_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i19024_4_lut_LC_7_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__48037\,
            in1 => \N__23085\,
            in2 => \N__23014\,
            in3 => \N__29791\,
            lcout => OPEN,
            ltout => \ADC_VAC.n21031_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.adc_state_i0_LC_7_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000001110100"
        )
    port map (
            in0 => \N__29792\,
            in1 => \N__29862\,
            in2 => \N__23011\,
            in3 => \N__48038\,
            lcout => adc_state_0_adj_1411,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55206\,
            ce => \N__23008\,
            sr => \_gnd_net_\
        );

    \ADC_VAC.i30_4_lut_LC_7_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000110000001"
        )
    port map (
            in0 => \N__30142\,
            in1 => \N__29847\,
            in2 => \N__29793\,
            in3 => \N__22998\,
            lcout => OPEN,
            ltout => \ADC_VAC.n17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i19101_2_lut_LC_7_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22954\,
            in3 => \N__48036\,
            lcout => \ADC_VAC.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.bit_cnt_i0_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22942\,
            in2 => \_gnd_net_\,
            in3 => \N__22930\,
            lcout => \ADC_VAC.bit_cnt_0\,
            ltout => OPEN,
            carryin => \bfn_7_17_0_\,
            carryout => \ADC_VAC.n19357\,
            clk => \N__55218\,
            ce => \N__23041\,
            sr => \N__23029\
        );

    \ADC_VAC.bit_cnt_i1_LC_7_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22926\,
            in2 => \_gnd_net_\,
            in3 => \N__22912\,
            lcout => \ADC_VAC.bit_cnt_1\,
            ltout => OPEN,
            carryin => \ADC_VAC.n19357\,
            carryout => \ADC_VAC.n19358\,
            clk => \N__55218\,
            ce => \N__23041\,
            sr => \N__23029\
        );

    \ADC_VAC.bit_cnt_i2_LC_7_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23134\,
            in2 => \_gnd_net_\,
            in3 => \N__23122\,
            lcout => \ADC_VAC.bit_cnt_2\,
            ltout => OPEN,
            carryin => \ADC_VAC.n19358\,
            carryout => \ADC_VAC.n19359\,
            clk => \N__55218\,
            ce => \N__23041\,
            sr => \N__23029\
        );

    \ADC_VAC.bit_cnt_i3_LC_7_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23119\,
            in2 => \_gnd_net_\,
            in3 => \N__23107\,
            lcout => \ADC_VAC.bit_cnt_3\,
            ltout => OPEN,
            carryin => \ADC_VAC.n19359\,
            carryout => \ADC_VAC.n19360\,
            clk => \N__55218\,
            ce => \N__23041\,
            sr => \N__23029\
        );

    \ADC_VAC.bit_cnt_i4_LC_7_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23103\,
            in2 => \_gnd_net_\,
            in3 => \N__23089\,
            lcout => \ADC_VAC.bit_cnt_4\,
            ltout => OPEN,
            carryin => \ADC_VAC.n19360\,
            carryout => \ADC_VAC.n19361\,
            clk => \N__55218\,
            ce => \N__23041\,
            sr => \N__23029\
        );

    \ADC_VAC.bit_cnt_i5_LC_7_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23086\,
            in2 => \_gnd_net_\,
            in3 => \N__23074\,
            lcout => \ADC_VAC.bit_cnt_5\,
            ltout => OPEN,
            carryin => \ADC_VAC.n19361\,
            carryout => \ADC_VAC.n19362\,
            clk => \N__55218\,
            ce => \N__23041\,
            sr => \N__23029\
        );

    \ADC_VAC.bit_cnt_i6_LC_7_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23071\,
            in2 => \_gnd_net_\,
            in3 => \N__23059\,
            lcout => \ADC_VAC.bit_cnt_6\,
            ltout => OPEN,
            carryin => \ADC_VAC.n19362\,
            carryout => \ADC_VAC.n19363\,
            clk => \N__55218\,
            ce => \N__23041\,
            sr => \N__23029\
        );

    \ADC_VAC.bit_cnt_i7_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23053\,
            in2 => \_gnd_net_\,
            in3 => \N__23056\,
            lcout => \ADC_VAC.bit_cnt_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55218\,
            ce => \N__23041\,
            sr => \N__23029\
        );

    \ADC_IAC.i1_3_lut_LC_7_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__25007\,
            in1 => \N__50645\,
            in2 => \_gnd_net_\,
            in3 => \N__24657\,
            lcout => n12542,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.adc_state_i2_LC_7_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001110001000"
        )
    port map (
            in0 => \N__50647\,
            in1 => \N__29999\,
            in2 => \_gnd_net_\,
            in3 => \N__29930\,
            lcout => \DTRIG_N_910\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55229\,
            ce => \N__24955\,
            sr => \_gnd_net_\
        );

    \ADC_IAC.adc_state_i1_LC_7_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001010101"
        )
    port map (
            in0 => \N__29931\,
            in1 => \_gnd_net_\,
            in2 => \N__30013\,
            in3 => \N__50648\,
            lcout => adc_state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55229\,
            ce => \N__24955\,
            sr => \_gnd_net_\
        );

    \ADC_IAC.i1_2_lut_LC_7_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29990\,
            in2 => \_gnd_net_\,
            in3 => \N__29927\,
            lcout => n20553,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i1_4_lut_adj_6_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010010"
        )
    port map (
            in0 => \N__29928\,
            in1 => \N__25008\,
            in2 => \N__30012\,
            in3 => \N__50646\,
            lcout => \ADC_IAC.n12459\,
            ltout => \ADC_IAC.n12459_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i12394_2_lut_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23155\,
            in3 => \N__29995\,
            lcout => \ADC_IAC.n14791\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_83_LC_7_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29994\,
            in2 => \_gnd_net_\,
            in3 => \N__29929\,
            lcout => n20543,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.bit_cnt_i0_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24745\,
            in2 => \_gnd_net_\,
            in3 => \N__23152\,
            lcout => \ADC_IAC.bit_cnt_0\,
            ltout => OPEN,
            carryin => \bfn_7_19_0_\,
            carryout => \ADC_IAC.n19350\,
            clk => \N__55239\,
            ce => \N__23254\,
            sr => \N__23239\
        );

    \ADC_IAC.bit_cnt_i1_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24783\,
            in2 => \_gnd_net_\,
            in3 => \N__23149\,
            lcout => \ADC_IAC.bit_cnt_1\,
            ltout => OPEN,
            carryin => \ADC_IAC.n19350\,
            carryout => \ADC_IAC.n19351\,
            clk => \N__55239\,
            ce => \N__23254\,
            sr => \N__23239\
        );

    \ADC_IAC.bit_cnt_i2_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24769\,
            in2 => \_gnd_net_\,
            in3 => \N__23146\,
            lcout => \ADC_IAC.bit_cnt_2\,
            ltout => OPEN,
            carryin => \ADC_IAC.n19351\,
            carryout => \ADC_IAC.n19352\,
            clk => \N__55239\,
            ce => \N__23254\,
            sr => \N__23239\
        );

    \ADC_IAC.bit_cnt_i3_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24796\,
            in2 => \_gnd_net_\,
            in3 => \N__23143\,
            lcout => \ADC_IAC.bit_cnt_3\,
            ltout => OPEN,
            carryin => \ADC_IAC.n19352\,
            carryout => \ADC_IAC.n19353\,
            clk => \N__55239\,
            ce => \N__23254\,
            sr => \N__23239\
        );

    \ADC_IAC.bit_cnt_i4_LC_7_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24808\,
            in2 => \_gnd_net_\,
            in3 => \N__23140\,
            lcout => \ADC_IAC.bit_cnt_4\,
            ltout => OPEN,
            carryin => \ADC_IAC.n19353\,
            carryout => \ADC_IAC.n19354\,
            clk => \N__55239\,
            ce => \N__23254\,
            sr => \N__23239\
        );

    \ADC_IAC.bit_cnt_i5_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25041\,
            in2 => \_gnd_net_\,
            in3 => \N__23137\,
            lcout => \ADC_IAC.bit_cnt_5\,
            ltout => OPEN,
            carryin => \ADC_IAC.n19354\,
            carryout => \ADC_IAC.n19355\,
            clk => \N__55239\,
            ce => \N__23254\,
            sr => \N__23239\
        );

    \ADC_IAC.bit_cnt_i6_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24757\,
            in2 => \_gnd_net_\,
            in3 => \N__23260\,
            lcout => \ADC_IAC.bit_cnt_6\,
            ltout => OPEN,
            carryin => \ADC_IAC.n19355\,
            carryout => \ADC_IAC.n19356\,
            clk => \N__55239\,
            ce => \N__23254\,
            sr => \N__23239\
        );

    \ADC_IAC.bit_cnt_i7_LC_7_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24730\,
            in2 => \_gnd_net_\,
            in3 => \N__23257\,
            lcout => \ADC_IAC.bit_cnt_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55239\,
            ce => \N__23254\,
            sr => \N__23239\
        );

    \ADC_VDC.i1_2_lut_adj_42_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34588\,
            in2 => \_gnd_net_\,
            in3 => \N__34361\,
            lcout => \ADC_VDC.n20345\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19022_2_lut_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23229\,
            in2 => \_gnd_net_\,
            in3 => \N__23205\,
            lcout => n21206,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i9_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__34365\,
            in1 => \N__25078\,
            in2 => \N__26884\,
            in3 => \N__26509\,
            lcout => cmd_rdadctmp_9_adj_1463,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32904\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i3_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__28361\,
            in1 => \N__34629\,
            in2 => \N__23172\,
            in3 => \N__25222\,
            lcout => buf_adcdata_vdc_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32904\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i7_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__34364\,
            in1 => \N__26528\,
            in2 => \N__26883\,
            in3 => \N__25122\,
            lcout => cmd_rdadctmp_7_adj_1465,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32904\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i10_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__25077\,
            in1 => \N__34366\,
            in2 => \N__26988\,
            in3 => \N__26850\,
            lcout => cmd_rdadctmp_10_adj_1462,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32904\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i6_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__34363\,
            in1 => \N__25121\,
            in2 => \N__26882\,
            in3 => \N__25149\,
            lcout => cmd_rdadctmp_6_adj_1466,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32904\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.i23_4_lut_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110110011001"
        )
    port map (
            in0 => \N__28943\,
            in1 => \N__28775\,
            in2 => \N__28677\,
            in3 => \N__28611\,
            lcout => \CLK_DDS.n9_adj_1386\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i5_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__34362\,
            in1 => \N__25148\,
            in2 => \N__26881\,
            in3 => \N__26569\,
            lcout => cmd_rdadctmp_5_adj_1467,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32904\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i15_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__26450\,
            in1 => \N__34367\,
            in2 => \N__25252\,
            in3 => \N__26851\,
            lcout => cmd_rdadctmp_15_adj_1457,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32904\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i14_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__34370\,
            in1 => \N__25287\,
            in2 => \N__25248\,
            in3 => \N__26888\,
            lcout => cmd_rdadctmp_14_adj_1458,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32886\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i0_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__28362\,
            in1 => \N__34631\,
            in2 => \N__23499\,
            in3 => \N__25318\,
            lcout => buf_adcdata_vdc_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32886\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i18_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__34371\,
            in1 => \N__25193\,
            in2 => \N__26485\,
            in3 => \N__26889\,
            lcout => cmd_rdadctmp_18_adj_1454,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32886\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i1_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__28364\,
            in1 => \N__34633\,
            in2 => \N__23985\,
            in3 => \N__25303\,
            lcout => buf_adcdata_vdc_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32886\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i19_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__34372\,
            in1 => \N__26915\,
            in2 => \N__25198\,
            in3 => \N__26890\,
            lcout => cmd_rdadctmp_19_adj_1453,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32886\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i10_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__28363\,
            in1 => \N__34632\,
            in2 => \N__24072\,
            in3 => \N__25444\,
            lcout => buf_adcdata_vdc_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32886\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i21_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__34373\,
            in1 => \N__25463\,
            in2 => \N__26773\,
            in3 => \N__26891\,
            lcout => cmd_rdadctmp_21_adj_1451,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32886\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i13_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__25286\,
            in1 => \N__26363\,
            in2 => \N__26895\,
            in3 => \N__34374\,
            lcout => cmd_rdadctmp_13_adj_1459,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32886\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i22_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101000001010"
        )
    port map (
            in0 => \N__25424\,
            in1 => \N__34369\,
            in2 => \N__26896\,
            in3 => \N__25464\,
            lcout => cmd_rdadctmp_22_adj_1450,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32872\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i21_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__25519\,
            in1 => \N__34640\,
            in2 => \N__23367\,
            in3 => \N__28397\,
            lcout => buf_adcdata_vdc_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32908\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i20_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__34636\,
            in1 => \N__28419\,
            in2 => \N__25668\,
            in3 => \N__25534\,
            lcout => buf_adcdata_vdc_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32908\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i13_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__28414\,
            in1 => \N__34637\,
            in2 => \N__23343\,
            in3 => \N__25378\,
            lcout => buf_adcdata_vdc_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32908\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i18_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__34635\,
            in1 => \N__28418\,
            in2 => \N__23874\,
            in3 => \N__25564\,
            lcout => buf_adcdata_vdc_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32908\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i16_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__28415\,
            in1 => \N__34638\,
            in2 => \N__23325\,
            in3 => \N__25333\,
            lcout => buf_adcdata_vdc_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32908\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i2_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__25270\,
            in1 => \N__28420\,
            in2 => \N__23307\,
            in3 => \N__34641\,
            lcout => buf_adcdata_vdc_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32908\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i19_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__28416\,
            in1 => \N__34639\,
            in2 => \N__23286\,
            in3 => \N__25549\,
            lcout => buf_adcdata_vdc_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32908\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i15_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__34634\,
            in1 => \N__28417\,
            in2 => \N__23577\,
            in3 => \N__25348\,
            lcout => buf_adcdata_vdc_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32908\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i14_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111100100000"
        )
    port map (
            in0 => \N__25363\,
            in1 => \N__34627\,
            in2 => \N__28398\,
            in3 => \N__23553\,
            lcout => buf_adcdata_vdc_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32885\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i22_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__34625\,
            in1 => \N__28390\,
            in2 => \N__23541\,
            in3 => \N__25504\,
            lcout => buf_adcdata_vdc_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32885\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i17_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__28388\,
            in1 => \N__34626\,
            in2 => \N__23523\,
            in3 => \N__25579\,
            lcout => buf_adcdata_vdc_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32885\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_0_i19_3_lut_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23500\,
            in1 => \N__23478\,
            in2 => \_gnd_net_\,
            in3 => \N__56960\,
            lcout => OPEN,
            ltout => \n19_adj_1477_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_0_i22_3_lut_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23457\,
            in2 => \N__23431\,
            in3 => \N__47774\,
            lcout => n22_adj_1476,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19506_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__29317\,
            in1 => \N__57183\,
            in2 => \N__23428\,
            in3 => \N__56959\,
            lcout => n22141,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i23_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__28389\,
            in1 => \N__27055\,
            in2 => \N__24309\,
            in3 => \N__34628\,
            lcout => buf_adcdata_vdc_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32885\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19388_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__56885\,
            in1 => \N__23398\,
            in2 => \N__57465\,
            in3 => \N__23805\,
            lcout => OPEN,
            ltout => \n21931_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n21931_bdd_4_lut_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__23878\,
            in1 => \N__23857\,
            in2 => \N__23830\,
            in3 => \N__57345\,
            lcout => n21934,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i2_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__52190\,
            in1 => \N__45329\,
            in2 => \N__38729\,
            in3 => \N__23806\,
            lcout => \buf_cfgRTD_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55114\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i3_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__45330\,
            in1 => \N__52191\,
            in2 => \N__43760\,
            in3 => \N__23763\,
            lcout => \buf_cfgRTD_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55114\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i0_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__52189\,
            in1 => \N__45328\,
            in2 => \N__43504\,
            in3 => \N__23718\,
            lcout => \buf_cfgRTD_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55114\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12100_2_lut_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__54721\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54091\,
            lcout => n14490,
            ltout => \n14490_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i1_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__57346\,
            in1 => \N__35991\,
            in2 => \N__23701\,
            in3 => \N__30939\,
            lcout => comm_cmd_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55114\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19526_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__23680\,
            in1 => \N__57341\,
            in2 => \N__23659\,
            in3 => \N__56884\,
            lcout => n22165,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_1_i22_3_lut_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__47743\,
            in1 => \N__23629\,
            in2 => \_gnd_net_\,
            in3 => \N__23941\,
            lcout => OPEN,
            ltout => \n22_adj_1618_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_1_i30_3_lut_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23596\,
            in2 => \N__23584\,
            in3 => \N__56345\,
            lcout => n30_adj_1619,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18186_4_lut_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110110101000"
        )
    port map (
            in0 => \N__57186\,
            in1 => \N__56685\,
            in2 => \N__24004\,
            in3 => \N__41449\,
            lcout => OPEN,
            ltout => \n20781_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_2__bdd_4_lut_19360_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__23932\,
            in1 => \N__47744\,
            in2 => \N__23989\,
            in3 => \N__56346\,
            lcout => n21943,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_1_i19_3_lut_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__23986\,
            in1 => \N__23961\,
            in2 => \_gnd_net_\,
            in3 => \N__56684\,
            lcout => n19_adj_1617,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19536_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__56683\,
            in1 => \N__41899\,
            in2 => \N__30463\,
            in3 => \N__57184\,
            lcout => OPEN,
            ltout => \n22171_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22171_bdd_4_lut_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__57185\,
            in1 => \N__50299\,
            in2 => \N__23935\,
            in3 => \N__31537\,
            lcout => n20775,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15210_2_lut_3_lut_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__30803\,
            in1 => \N__51284\,
            in2 => \_gnd_net_\,
            in3 => \N__54092\,
            lcout => n14_adj_1523,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_2__bdd_4_lut_19433_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__23923\,
            in1 => \N__47789\,
            in2 => \N__23911\,
            in3 => \N__56338\,
            lcout => OPEN,
            ltout => \n22051_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22051_bdd_4_lut_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__56339\,
            in1 => \N__24205\,
            in2 => \N__23899\,
            in3 => \N__23896\,
            lcout => n22054,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n21967_bdd_4_lut_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__56340\,
            in1 => \N__23887\,
            in2 => \N__26008\,
            in3 => \N__25612\,
            lcout => n21970,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i25_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__37869\,
            in1 => \N__24256\,
            in2 => \N__48280\,
            in3 => \N__24230\,
            lcout => cmd_rdadctmp_25_adj_1418,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55135\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i20_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__24128\,
            in1 => \N__48219\,
            in2 => \N__24031\,
            in3 => \N__37868\,
            lcout => cmd_rdadctmp_20_adj_1423,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55135\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22039_bdd_4_lut_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__27613\,
            in1 => \N__24214\,
            in2 => \N__32272\,
            in3 => \N__57440\,
            lcout => n22042,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i7_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__45727\,
            in1 => \N__45327\,
            in2 => \_gnd_net_\,
            in3 => \N__24166\,
            lcout => \buf_cfgRTD_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55148\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i12_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__24090\,
            in1 => \N__48480\,
            in2 => \N__24138\,
            in3 => \N__48217\,
            lcout => buf_adcdata_vac_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55148\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i10_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__48216\,
            in1 => \N__24112\,
            in2 => \N__48511\,
            in3 => \N__24045\,
            lcout => buf_adcdata_vac_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55148\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_4_i19_3_lut_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26734\,
            in1 => \N__24089\,
            in2 => \_gnd_net_\,
            in3 => \N__56725\,
            lcout => n19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_2_i19_3_lut_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__24076\,
            in1 => \N__24044\,
            in2 => \_gnd_net_\,
            in3 => \N__56726\,
            lcout => n19_adj_1505,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i11_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__48438\,
            in1 => \N__48218\,
            in2 => \N__24030\,
            in3 => \N__25893\,
            lcout => buf_adcdata_vac_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55163\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_7_i26_3_lut_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__31306\,
            in1 => \N__56639\,
            in2 => \_gnd_net_\,
            in3 => \N__30100\,
            lcout => OPEN,
            ltout => \n26_adj_1511_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18239_4_lut_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__56641\,
            in1 => \N__24394\,
            in2 => \N__24376\,
            in3 => \N__57436\,
            lcout => OPEN,
            ltout => \n20834_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_2__bdd_4_lut_19442_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__56334\,
            in1 => \N__29032\,
            in2 => \N__24373\,
            in3 => \N__47753\,
            lcout => OPEN,
            ltout => \n22057_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22057_bdd_4_lut_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001010"
        )
    port map (
            in0 => \N__27892\,
            in1 => \N__24292\,
            in2 => \N__24370\,
            in3 => \N__56335\,
            lcout => n22060,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19020_2_lut_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24367\,
            in2 => \_gnd_net_\,
            in3 => \N__56640\,
            lcout => n21261,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22135_bdd_4_lut_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111010100100"
        )
    port map (
            in0 => \N__24355\,
            in1 => \N__24342\,
            in2 => \N__57524\,
            in3 => \N__24310\,
            lcout => n20831,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i7_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__50500\,
            in1 => \N__24279\,
            in2 => \N__24562\,
            in3 => \N__50921\,
            lcout => cmd_rdadctmp_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55178\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i21_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__50919\,
            in1 => \N__48975\,
            in2 => \N__24646\,
            in3 => \N__27287\,
            lcout => buf_adcdata_iac_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55178\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_1_i16_3_lut_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__31932\,
            in1 => \N__32239\,
            in2 => \_gnd_net_\,
            in3 => \N__56698\,
            lcout => n16_adj_1507,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i8_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__54718\,
            in1 => \N__24433\,
            in2 => \N__52167\,
            in3 => \N__42382\,
            lcout => data_index_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55178\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i6_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__50920\,
            in1 => \N__24558\,
            in2 => \N__24718\,
            in3 => \N__50501\,
            lcout => cmd_rdadctmp_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55178\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_354_Mux_8_i15_4_lut_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__54717\,
            in1 => \N__24432\,
            in2 => \N__52166\,
            in3 => \N__42381\,
            lcout => \data_index_9_N_212_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_6__I_0_368_i8_2_lut_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57388\,
            in2 => \_gnd_net_\,
            in3 => \N__47748\,
            lcout => n8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i19_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__50759\,
            in1 => \N__48968\,
            in2 => \N__24616\,
            in3 => \N__26069\,
            lcout => buf_adcdata_iac_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55193\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i23_LC_8_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__50469\,
            in1 => \N__24454\,
            in2 => \N__50837\,
            in3 => \N__25856\,
            lcout => cmd_rdadctmp_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55193\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6362_3_lut_LC_8_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43487\,
            in1 => \N__42396\,
            in2 => \_gnd_net_\,
            in3 => \N__43300\,
            lcout => n8_adj_1534,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i7_LC_8_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__54724\,
            in1 => \N__30078\,
            in2 => \N__52170\,
            in3 => \N__42439\,
            lcout => data_index_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55193\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i8_LC_8_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__50746\,
            in1 => \N__48894\,
            in2 => \N__45138\,
            in3 => \N__24413\,
            lcout => buf_adcdata_iac_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55207\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i27_LC_8_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__50415\,
            in1 => \N__27757\,
            in2 => \N__50834\,
            in3 => \N__24611\,
            lcout => cmd_rdadctmp_27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55207\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i1_LC_8_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101000001010"
        )
    port map (
            in0 => \N__24666\,
            in1 => \N__24574\,
            in2 => \N__50470\,
            in3 => \N__50749\,
            lcout => cmd_rdadctmp_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55207\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i5_LC_8_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__50417\,
            in1 => \N__24886\,
            in2 => \N__50836\,
            in3 => \N__24711\,
            lcout => cmd_rdadctmp_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55207\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i22_LC_8_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__48893\,
            in1 => \N__50747\,
            in2 => \N__24904\,
            in3 => \N__24683\,
            lcout => buf_adcdata_iac_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55207\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i2_LC_8_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__50416\,
            in1 => \N__24667\,
            in2 => \N__50835\,
            in3 => \N__24870\,
            lcout => cmd_rdadctmp_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55207\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i30_LC_8_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__24899\,
            in1 => \N__50748\,
            in2 => \N__24644\,
            in3 => \N__50418\,
            lcout => cmd_rdadctmp_30,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55207\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.CS_37_LC_8_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010001010101"
        )
    port map (
            in0 => \N__24820\,
            in1 => \N__50714\,
            in2 => \N__25012\,
            in3 => \N__24658\,
            lcout => \IAC_CS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55219\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i29_LC_8_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__50712\,
            in1 => \N__50458\,
            in2 => \N__24645\,
            in3 => \N__28157\,
            lcout => cmd_rdadctmp_29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55219\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i28_LC_8_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__50454\,
            in1 => \N__50715\,
            in2 => \N__28161\,
            in3 => \N__24612\,
            lcout => cmd_rdadctmp_28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55219\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i0_LC_8_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__50711\,
            in1 => \N__50457\,
            in2 => \N__24595\,
            in3 => \N__24573\,
            lcout => cmd_rdadctmp_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55219\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i31_LC_8_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__50455\,
            in1 => \N__50716\,
            in2 => \N__26292\,
            in3 => \N__24903\,
            lcout => cmd_rdadctmp_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55219\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i4_LC_8_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__50713\,
            in1 => \N__50459\,
            in2 => \N__24859\,
            in3 => \N__24885\,
            lcout => cmd_rdadctmp_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55219\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i3_LC_8_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__50456\,
            in1 => \N__24855\,
            in2 => \N__24874\,
            in3 => \N__50717\,
            lcout => cmd_rdadctmp_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55219\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_207_LC_8_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000110"
        )
    port map (
            in0 => \N__50710\,
            in1 => \N__30005\,
            in2 => \N__24837\,
            in3 => \N__29936\,
            lcout => n14_adj_1581,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i1_2_lut_adj_5_LC_8_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29934\,
            in2 => \_gnd_net_\,
            in3 => \N__24814\,
            lcout => \ADC_IAC.n20670\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i1_4_lut_LC_8_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101111101111"
        )
    port map (
            in0 => \N__50649\,
            in1 => \N__30003\,
            in2 => \N__24997\,
            in3 => \N__30139\,
            lcout => \ADC_IAC.n20669\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i18158_4_lut_LC_8_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24807\,
            in1 => \N__24795\,
            in2 => \N__24784\,
            in3 => \N__24768\,
            lcout => OPEN,
            ltout => \ADC_IAC.n20753_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i18170_4_lut_LC_8_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__24756\,
            in1 => \N__24744\,
            in2 => \N__24733\,
            in3 => \N__24729\,
            lcout => OPEN,
            ltout => \ADC_IAC.n20765_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i18788_4_lut_LC_8_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__25042\,
            in1 => \N__50651\,
            in2 => \N__25027\,
            in3 => \N__29933\,
            lcout => OPEN,
            ltout => \ADC_IAC.n21007_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.adc_state_i0_LC_8_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000111110000"
        )
    port map (
            in0 => \N__29935\,
            in1 => \N__50724\,
            in2 => \N__25024\,
            in3 => \N__30004\,
            lcout => adc_state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55230\,
            ce => \N__25021\,
            sr => \_gnd_net_\
        );

    \ADC_IAC.i30_4_lut_LC_8_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110000000101"
        )
    port map (
            in0 => \N__30140\,
            in1 => \N__24989\,
            in2 => \N__30014\,
            in3 => \N__29932\,
            lcout => OPEN,
            ltout => \ADC_IAC.n17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.i19104_2_lut_LC_8_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110101111"
        )
    port map (
            in0 => \N__50650\,
            in1 => \_gnd_net_\,
            in2 => \N__24958\,
            in3 => \_gnd_net_\,
            lcout => \ADC_IAC.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i23_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000101110"
        )
    port map (
            in0 => \N__25429\,
            in1 => \N__34121\,
            in2 => \N__25401\,
            in3 => \N__26308\,
            lcout => \ADC_VDC.cmd_rdadctmp_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32806\,
            ce => \N__26545\,
            sr => \N__24946\
        );

    \comm_spi.RESET_I_0_102_2_lut_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48744\,
            in2 => \_gnd_net_\,
            in3 => \N__55474\,
            lcout => \comm_spi.data_tx_7__N_772\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadcbuf_i0_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24931\,
            in2 => \N__26611\,
            in3 => \_gnd_net_\,
            lcout => \ADC_VDC.cmd_rdadcbuf_0\,
            ltout => OPEN,
            carryin => \bfn_9_5_0_\,
            carryout => \ADC_VDC.n19364\,
            clk => \N__32842\,
            ce => \N__29162\,
            sr => \N__29103\
        );

    \ADC_VDC.cmd_rdadcbuf_i1_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24925\,
            in2 => \N__26410\,
            in3 => \N__24919\,
            lcout => \ADC_VDC.cmd_rdadcbuf_1\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19364\,
            carryout => \ADC_VDC.n19365\,
            clk => \N__32842\,
            ce => \N__29162\,
            sr => \N__29103\
        );

    \ADC_VDC.cmd_rdadcbuf_i2_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26388\,
            in2 => \N__24916\,
            in3 => \N__24907\,
            lcout => \ADC_VDC.cmd_rdadcbuf_2\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19365\,
            carryout => \ADC_VDC.n19366\,
            clk => \N__32842\,
            ce => \N__29162\,
            sr => \N__29103\
        );

    \ADC_VDC.cmd_rdadcbuf_i3_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25168\,
            in2 => \N__26590\,
            in3 => \N__25162\,
            lcout => \ADC_VDC.cmd_rdadcbuf_3\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19366\,
            carryout => \ADC_VDC.n19367\,
            clk => \N__32842\,
            ce => \N__29162\,
            sr => \N__29103\
        );

    \ADC_VDC.cmd_rdadcbuf_i4_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25159\,
            in2 => \N__26568\,
            in3 => \N__25153\,
            lcout => \ADC_VDC.cmd_rdadcbuf_4\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19367\,
            carryout => \ADC_VDC.n19368\,
            clk => \N__32842\,
            ce => \N__29162\,
            sr => \N__29103\
        );

    \ADC_VDC.cmd_rdadcbuf_i5_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25132\,
            in2 => \N__25150\,
            in3 => \N__25126\,
            lcout => \ADC_VDC.cmd_rdadcbuf_5\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19368\,
            carryout => \ADC_VDC.n19369\,
            clk => \N__32842\,
            ce => \N__29162\,
            sr => \N__29103\
        );

    \ADC_VDC.cmd_rdadcbuf_i6_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25105\,
            in2 => \N__25123\,
            in3 => \N__25099\,
            lcout => \ADC_VDC.cmd_rdadcbuf_6\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19369\,
            carryout => \ADC_VDC.n19370\,
            clk => \N__32842\,
            ce => \N__29162\,
            sr => \N__29103\
        );

    \ADC_VDC.cmd_rdadcbuf_i7_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25096\,
            in2 => \N__26533\,
            in3 => \N__25090\,
            lcout => \ADC_VDC.cmd_rdadcbuf_7\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19370\,
            carryout => \ADC_VDC.n19371\,
            clk => \N__32842\,
            ce => \N__29162\,
            sr => \N__29103\
        );

    \ADC_VDC.cmd_rdadcbuf_i8_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25087\,
            in2 => \N__26508\,
            in3 => \N__25081\,
            lcout => \ADC_VDC.cmd_rdadcbuf_8\,
            ltout => OPEN,
            carryin => \bfn_9_6_0_\,
            carryout => \ADC_VDC.n19372\,
            clk => \N__32903\,
            ce => \N__29179\,
            sr => \N__29108\
        );

    \ADC_VDC.cmd_rdadcbuf_i9_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25076\,
            in2 => \N__25063\,
            in3 => \N__25054\,
            lcout => \ADC_VDC.cmd_rdadcbuf_9\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19372\,
            carryout => \ADC_VDC.n19373\,
            clk => \N__32903\,
            ce => \N__29179\,
            sr => \N__29108\
        );

    \ADC_VDC.cmd_rdadcbuf_i10_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25051\,
            in2 => \N__26984\,
            in3 => \N__25045\,
            lcout => \ADC_VDC.cmd_rdadcbuf_10\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19373\,
            carryout => \ADC_VDC.n19374\,
            clk => \N__32903\,
            ce => \N__29179\,
            sr => \N__29108\
        );

    \ADC_VDC.cmd_rdadcbuf_i11_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25317\,
            in2 => \N__26959\,
            in3 => \N__25306\,
            lcout => cmd_rdadcbuf_11,
            ltout => OPEN,
            carryin => \ADC_VDC.n19374\,
            carryout => \ADC_VDC.n19375\,
            clk => \N__32903\,
            ce => \N__29179\,
            sr => \N__29108\
        );

    \ADC_VDC.cmd_rdadcbuf_i12_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25302\,
            in2 => \N__26365\,
            in3 => \N__25291\,
            lcout => cmd_rdadcbuf_12,
            ltout => OPEN,
            carryin => \ADC_VDC.n19375\,
            carryout => \ADC_VDC.n19376\,
            clk => \N__32903\,
            ce => \N__29179\,
            sr => \N__29108\
        );

    \ADC_VDC.cmd_rdadcbuf_i13_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25266\,
            in2 => \N__25288\,
            in3 => \N__25255\,
            lcout => cmd_rdadcbuf_13,
            ltout => OPEN,
            carryin => \ADC_VDC.n19376\,
            carryout => \ADC_VDC.n19377\,
            clk => \N__32903\,
            ce => \N__29179\,
            sr => \N__29108\
        );

    \ADC_VDC.cmd_rdadcbuf_i14_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25221\,
            in2 => \N__25247\,
            in3 => \N__25210\,
            lcout => cmd_rdadcbuf_14,
            ltout => OPEN,
            carryin => \ADC_VDC.n19377\,
            carryout => \ADC_VDC.n19378\,
            clk => \N__32903\,
            ce => \N__29179\,
            sr => \N__29108\
        );

    \ADC_VDC.cmd_rdadcbuf_i15_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26670\,
            in2 => \N__26451\,
            in3 => \N__25207\,
            lcout => cmd_rdadcbuf_15,
            ltout => OPEN,
            carryin => \ADC_VDC.n19378\,
            carryout => \ADC_VDC.n19379\,
            clk => \N__32903\,
            ce => \N__29179\,
            sr => \N__29108\
        );

    \ADC_VDC.cmd_rdadcbuf_i16_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27087\,
            in2 => \N__26428\,
            in3 => \N__25204\,
            lcout => cmd_rdadcbuf_16,
            ltout => OPEN,
            carryin => \bfn_9_7_0_\,
            carryout => \ADC_VDC.n19380\,
            clk => \N__32896\,
            ce => \N__29191\,
            sr => \N__29104\
        );

    \ADC_VDC.cmd_rdadcbuf_i17_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27102\,
            in2 => \N__26481\,
            in3 => \N__25201\,
            lcout => cmd_rdadcbuf_17,
            ltout => OPEN,
            carryin => \ADC_VDC.n19380\,
            carryout => \ADC_VDC.n19381\,
            clk => \N__32896\,
            ce => \N__29191\,
            sr => \N__29104\
        );

    \ADC_VDC.cmd_rdadcbuf_i18_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27114\,
            in2 => \N__25197\,
            in3 => \N__25174\,
            lcout => cmd_rdadcbuf_18,
            ltout => OPEN,
            carryin => \ADC_VDC.n19381\,
            carryout => \ADC_VDC.n19382\,
            clk => \N__32896\,
            ce => \N__29191\,
            sr => \N__29104\
        );

    \ADC_VDC.cmd_rdadcbuf_i19_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26646\,
            in2 => \N__26919\,
            in3 => \N__25171\,
            lcout => cmd_rdadcbuf_19,
            ltout => OPEN,
            carryin => \ADC_VDC.n19382\,
            carryout => \ADC_VDC.n19383\,
            clk => \N__32896\,
            ce => \N__29191\,
            sr => \N__29104\
        );

    \ADC_VDC.cmd_rdadcbuf_i20_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26658\,
            in2 => \N__26769\,
            in3 => \N__25468\,
            lcout => cmd_rdadcbuf_20,
            ltout => OPEN,
            carryin => \ADC_VDC.n19383\,
            carryout => \ADC_VDC.n19384\,
            clk => \N__32896\,
            ce => \N__29191\,
            sr => \N__29104\
        );

    \ADC_VDC.cmd_rdadcbuf_i21_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25443\,
            in2 => \N__25465\,
            in3 => \N__25432\,
            lcout => cmd_rdadcbuf_21,
            ltout => OPEN,
            carryin => \ADC_VDC.n19384\,
            carryout => \ADC_VDC.n19385\,
            clk => \N__32896\,
            ce => \N__29191\,
            sr => \N__29104\
        );

    \ADC_VDC.cmd_rdadcbuf_i22_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26709\,
            in2 => \N__25428\,
            in3 => \N__25405\,
            lcout => cmd_rdadcbuf_22,
            ltout => OPEN,
            carryin => \ADC_VDC.n19385\,
            carryout => \ADC_VDC.n19386\,
            clk => \N__32896\,
            ce => \N__29191\,
            sr => \N__29104\
        );

    \ADC_VDC.cmd_rdadcbuf_i23_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26745\,
            in2 => \N__25402\,
            in3 => \N__25381\,
            lcout => cmd_rdadcbuf_23,
            ltout => OPEN,
            carryin => \ADC_VDC.n19386\,
            carryout => \ADC_VDC.n19387\,
            clk => \N__32896\,
            ce => \N__29191\,
            sr => \N__29104\
        );

    \ADC_VDC.cmd_rdadcbuf_i24_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25377\,
            in2 => \_gnd_net_\,
            in3 => \N__25366\,
            lcout => cmd_rdadcbuf_24,
            ltout => OPEN,
            carryin => \bfn_9_8_0_\,
            carryout => \ADC_VDC.n19388\,
            clk => \N__32894\,
            ce => \N__29186\,
            sr => \N__29113\
        );

    \ADC_VDC.cmd_rdadcbuf_i25_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25362\,
            in2 => \_gnd_net_\,
            in3 => \N__25351\,
            lcout => cmd_rdadcbuf_25,
            ltout => OPEN,
            carryin => \ADC_VDC.n19388\,
            carryout => \ADC_VDC.n19389\,
            clk => \N__32894\,
            ce => \N__29186\,
            sr => \N__29113\
        );

    \ADC_VDC.cmd_rdadcbuf_i26_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25347\,
            in2 => \_gnd_net_\,
            in3 => \N__25336\,
            lcout => cmd_rdadcbuf_26,
            ltout => OPEN,
            carryin => \ADC_VDC.n19389\,
            carryout => \ADC_VDC.n19390\,
            clk => \N__32894\,
            ce => \N__29186\,
            sr => \N__29113\
        );

    \ADC_VDC.cmd_rdadcbuf_i27_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25332\,
            in2 => \_gnd_net_\,
            in3 => \N__25321\,
            lcout => cmd_rdadcbuf_27,
            ltout => OPEN,
            carryin => \ADC_VDC.n19390\,
            carryout => \ADC_VDC.n19391\,
            clk => \N__32894\,
            ce => \N__29186\,
            sr => \N__29113\
        );

    \ADC_VDC.cmd_rdadcbuf_i28_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25578\,
            in2 => \_gnd_net_\,
            in3 => \N__25567\,
            lcout => cmd_rdadcbuf_28,
            ltout => OPEN,
            carryin => \ADC_VDC.n19391\,
            carryout => \ADC_VDC.n19392\,
            clk => \N__32894\,
            ce => \N__29186\,
            sr => \N__29113\
        );

    \ADC_VDC.cmd_rdadcbuf_i29_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25563\,
            in2 => \_gnd_net_\,
            in3 => \N__25552\,
            lcout => cmd_rdadcbuf_29,
            ltout => OPEN,
            carryin => \ADC_VDC.n19392\,
            carryout => \ADC_VDC.n19393\,
            clk => \N__32894\,
            ce => \N__29186\,
            sr => \N__29113\
        );

    \ADC_VDC.cmd_rdadcbuf_i30_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25548\,
            in2 => \_gnd_net_\,
            in3 => \N__25537\,
            lcout => cmd_rdadcbuf_30,
            ltout => OPEN,
            carryin => \ADC_VDC.n19393\,
            carryout => \ADC_VDC.n19394\,
            clk => \N__32894\,
            ce => \N__29186\,
            sr => \N__29113\
        );

    \ADC_VDC.cmd_rdadcbuf_i31_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25533\,
            in2 => \_gnd_net_\,
            in3 => \N__25522\,
            lcout => cmd_rdadcbuf_31,
            ltout => OPEN,
            carryin => \ADC_VDC.n19394\,
            carryout => \ADC_VDC.n19395\,
            clk => \N__32894\,
            ce => \N__29186\,
            sr => \N__29113\
        );

    \ADC_VDC.cmd_rdadcbuf_i32_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25518\,
            in2 => \_gnd_net_\,
            in3 => \N__25507\,
            lcout => cmd_rdadcbuf_32,
            ltout => OPEN,
            carryin => \bfn_9_9_0_\,
            carryout => \ADC_VDC.n19396\,
            clk => \N__32884\,
            ce => \N__29190\,
            sr => \N__29109\
        );

    \ADC_VDC.cmd_rdadcbuf_i33_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25503\,
            in2 => \_gnd_net_\,
            in3 => \N__25492\,
            lcout => cmd_rdadcbuf_33,
            ltout => OPEN,
            carryin => \ADC_VDC.n19396\,
            carryout => \ADC_VDC.n19397\,
            clk => \N__32884\,
            ce => \N__29190\,
            sr => \N__29109\
        );

    \ADC_VDC.add_23_36_lut_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27047\,
            in2 => \_gnd_net_\,
            in3 => \N__25489\,
            lcout => \ADC_VDC.cmd_rdadcbuf_35_N_1130_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n21943_bdd_4_lut_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__56272\,
            in1 => \N__25486\,
            in2 => \N__27940\,
            in3 => \N__25477\,
            lcout => OPEN,
            ltout => \n21946_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_0__i0_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__54099\,
            in1 => \_gnd_net_\,
            in2 => \N__25471\,
            in3 => \N__36255\,
            lcout => comm_buf_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55104\,
            ce => \N__27504\,
            sr => \N__27453\
        );

    \i15211_2_lut_3_lut_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__43461\,
            in1 => \N__51219\,
            in2 => \_gnd_net_\,
            in3 => \N__54097\,
            lcout => n14_adj_1524,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15203_2_lut_3_lut_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__38650\,
            in1 => \N__51218\,
            in2 => \_gnd_net_\,
            in3 => \N__54096\,
            lcout => n14_adj_1551,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15205_2_lut_3_lut_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__42623\,
            in1 => \N__51220\,
            in2 => \_gnd_net_\,
            in3 => \N__54098\,
            lcout => n14_adj_1525,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_0__i7_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54103\,
            in1 => \N__36896\,
            in2 => \_gnd_net_\,
            in3 => \N__25597\,
            lcout => comm_buf_0_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55115\,
            ce => \N__27512\,
            sr => \N__27465\
        );

    \comm_buf_0__i6_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35810\,
            in1 => \N__25588\,
            in2 => \_gnd_net_\,
            in3 => \N__54105\,
            lcout => comm_buf_0_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55115\,
            ce => \N__27512\,
            sr => \N__27465\
        );

    \comm_buf_0__i4_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54102\,
            in1 => \N__35668\,
            in2 => \_gnd_net_\,
            in3 => \N__25720\,
            lcout => comm_buf_0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55115\,
            ce => \N__27512\,
            sr => \N__27465\
        );

    \comm_buf_0__i3_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__35563\,
            in1 => \N__54104\,
            in2 => \_gnd_net_\,
            in3 => \N__41230\,
            lcout => comm_buf_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55115\,
            ce => \N__27512\,
            sr => \N__27465\
        );

    \comm_cmd_0__bdd_4_lut_19413_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010101010"
        )
    port map (
            in0 => \N__56562\,
            in1 => \N__38936\,
            in2 => \N__41656\,
            in3 => \N__57443\,
            lcout => OPEN,
            ltout => \n22015_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22015_bdd_4_lut_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011000010"
        )
    port map (
            in0 => \N__44031\,
            in1 => \N__57444\,
            in2 => \N__25582\,
            in3 => \N__36925\,
            lcout => n20871,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18223_3_lut_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__56563\,
            in1 => \N__31198\,
            in2 => \_gnd_net_\,
            in3 => \N__47311\,
            lcout => OPEN,
            ltout => \n20818_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18225_4_lut_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010111000"
        )
    port map (
            in0 => \N__25639\,
            in1 => \N__57445\,
            in2 => \N__25624\,
            in3 => \N__56567\,
            lcout => OPEN,
            ltout => \n20820_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_2__bdd_4_lut_19408_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__56344\,
            in1 => \N__25621\,
            in2 => \N__25615\,
            in3 => \N__47746\,
            lcout => n21967,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_0__i1_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__35995\,
            in1 => \N__54106\,
            in2 => \_gnd_net_\,
            in3 => \N__25606\,
            lcout => comm_buf_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55124\,
            ce => \N__27517\,
            sr => \N__27469\
        );

    \i36_4_lut_4_lut_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010010010101110"
        )
    port map (
            in0 => \N__56343\,
            in1 => \N__57442\,
            in2 => \N__56699\,
            in3 => \N__47745\,
            lcout => n30,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19398_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__56635\,
            in1 => \N__26100\,
            in2 => \N__28134\,
            in3 => \N__57242\,
            lcout => OPEN,
            ltout => \n22003_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22003_bdd_4_lut_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001111100000"
        )
    port map (
            in0 => \N__27587\,
            in1 => \N__57250\,
            in2 => \N__25600\,
            in3 => \N__33864\,
            lcout => n22006,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i24_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__50512\,
            in1 => \N__25982\,
            in2 => \N__25873\,
            in3 => \N__50882\,
            lcout => cmd_rdadctmp_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55136\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i0_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__30943\,
            in1 => \N__56637\,
            in2 => \N__30993\,
            in3 => \N__36259\,
            lcout => comm_cmd_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55136\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_4_lut_adj_101_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__56636\,
            in1 => \N__57241\,
            in2 => \N__45381\,
            in3 => \N__47747\,
            lcout => n20624,
            ltout => \n20624_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_90_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111101000101"
        )
    port map (
            in0 => \N__52168\,
            in1 => \N__49239\,
            in2 => \N__25765\,
            in3 => \N__54722\,
            lcout => n11417,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19057_2_lut_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__31357\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56634\,
            lcout => n20936,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.i4_4_lut_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__55695\,
            in1 => \N__25910\,
            in2 => \N__25937\,
            in3 => \N__43677\,
            lcout => OPEN,
            ltout => \SIG_DDS.n10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.dds_state_i0_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000000010110011"
        )
    port map (
            in0 => \N__25774\,
            in1 => \N__55655\,
            in2 => \N__25762\,
            in3 => \N__55696\,
            lcout => dds_state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55149\,
            ce => \N__45538\,
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__42045\,
            in1 => \N__57386\,
            in2 => \N__25759\,
            in3 => \N__56642\,
            lcout => n22207,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_2__bdd_4_lut_19428_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__56374\,
            in1 => \N__47752\,
            in2 => \N__28999\,
            in3 => \N__56336\,
            lcout => OPEN,
            ltout => \n22027_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22027_bdd_4_lut_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__56337\,
            in1 => \N__25729\,
            in2 => \N__25723\,
            in3 => \N__25645\,
            lcout => n22030,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22207_bdd_4_lut_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001000100"
        )
    port map (
            in0 => \N__57387\,
            in1 => \N__25710\,
            in2 => \N__25675\,
            in3 => \N__25651\,
            lcout => n20801,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.bit_cnt_i3_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__43687\,
            in1 => \N__25912\,
            in2 => \N__25939\,
            in3 => \N__25786\,
            lcout => \SIG_DDS.bit_cnt_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55164\,
            ce => \N__55672\,
            sr => \N__43711\
        );

    \SIG_DDS.bit_cnt_i1_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25930\,
            in2 => \_gnd_net_\,
            in3 => \N__43685\,
            lcout => \SIG_DDS.bit_cnt_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55164\,
            ce => \N__55672\,
            sr => \N__43711\
        );

    \i18250_3_lut_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__25968\,
            in1 => \N__31945\,
            in2 => \_gnd_net_\,
            in3 => \N__57391\,
            lcout => n20845,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.bit_cnt_i2_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101111110100000"
        )
    port map (
            in0 => \N__43686\,
            in1 => \_gnd_net_\,
            in2 => \N__25938\,
            in3 => \N__25911\,
            lcout => \SIG_DDS.bit_cnt_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55164\,
            ce => \N__55672\,
            sr => \N__43711\
        );

    \mux_129_Mux_3_i16_3_lut_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__56694\,
            in1 => \N__31827\,
            in2 => \_gnd_net_\,
            in3 => \N__36713\,
            lcout => n16_adj_1500,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_3_i19_3_lut_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__26698\,
            in1 => \N__25889\,
            in2 => \_gnd_net_\,
            in3 => \N__56693\,
            lcout => n19_adj_1501,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i15_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__48969\,
            in1 => \N__50801\,
            in2 => \N__25872\,
            in3 => \N__31979\,
            lcout => buf_adcdata_iac_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55179\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_adj_261_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__54719\,
            in1 => \N__39187\,
            in2 => \N__25840\,
            in3 => \N__53536\,
            lcout => n10503,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22117_bdd_4_lut_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100010"
        )
    port map (
            in0 => \N__28237\,
            in1 => \N__25831\,
            in2 => \N__25819\,
            in3 => \N__47824\,
            lcout => n22120,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.i18704_2_lut_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__25785\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55887\,
            lcout => \SIG_DDS.n21292\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i5_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__42144\,
            in1 => \N__39236\,
            in2 => \_gnd_net_\,
            in3 => \N__26096\,
            lcout => \VAC_OSR0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55179\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19467_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__28085\,
            in1 => \N__57370\,
            in2 => \N__26070\,
            in3 => \N__56686\,
            lcout => n22075,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i17_LC_9_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__26027\,
            in1 => \N__27777\,
            in2 => \N__50937\,
            in3 => \N__48960\,
            lcout => buf_adcdata_iac_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55194\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \trig_dds0_304_LC_9_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__52111\,
            in1 => \N__26047\,
            in2 => \N__53005\,
            in3 => \N__54720\,
            lcout => trig_dds0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55194\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19556_LC_9_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__28050\,
            in1 => \N__57389\,
            in2 => \N__26031\,
            in3 => \N__56802\,
            lcout => OPEN,
            ltout => \n22201_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22201_bdd_4_lut_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__57390\,
            in1 => \N__32336\,
            in2 => \N__26011\,
            in3 => \N__27571\,
            lcout => n20805,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_start_329_LC_9_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__43474\,
            in1 => \N__29879\,
            in2 => \_gnd_net_\,
            in3 => \N__30442\,
            lcout => eis_start,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55194\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i16_LC_9_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__48959\,
            in1 => \N__50884\,
            in2 => \N__27993\,
            in3 => \N__25992\,
            lcout => buf_adcdata_iac_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55194\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i25_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__27773\,
            in1 => \N__50951\,
            in2 => \N__25993\,
            in3 => \N__50453\,
            lcout => cmd_rdadctmp_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55208\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19447_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__26207\,
            in1 => \N__57484\,
            in2 => \N__26262\,
            in3 => \N__56801\,
            lcout => n22045,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i23_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__50949\,
            in1 => \N__48911\,
            in2 => \N__26293\,
            in3 => \N__26258\,
            lcout => buf_adcdata_iac_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55208\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_rst_I_0_1_lut_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32101\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \AC_ADC_SYNC\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i8_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__45765\,
            in1 => \N__39237\,
            in2 => \_gnd_net_\,
            in3 => \N__26208\,
            lcout => \VAC_FLT1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55208\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i18_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__48910\,
            in1 => \N__50950\,
            in2 => \N__27756\,
            in3 => \N__27800\,
            lcout => buf_adcdata_iac_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55208\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.SCLK_35_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101000011100100"
        )
    port map (
            in0 => \N__50723\,
            in1 => \N__30021\,
            in2 => \N__26184\,
            in3 => \N__29950\,
            lcout => \IAC_SCLK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55220\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i11_3_lut_LC_10_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__27013\,
            in1 => \N__28276\,
            in2 => \_gnd_net_\,
            in3 => \N__27022\,
            lcout => \ADC_VDC.n18394\,
            ltout => \ADC_VDC.n18394_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i15984_3_lut_LC_10_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34773\,
            in2 => \N__26167\,
            in3 => \N__34114\,
            lcout => \ADC_VDC.n18397\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \EIS_SYNCCLK_I_0_1_lut_LC_10_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26164\,
            lcout => \IAC_CLK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i37_4_lut_LC_10_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011001000110"
        )
    port map (
            in0 => \N__34770\,
            in1 => \N__34876\,
            in2 => \N__34148\,
            in3 => \N__30679\,
            lcout => OPEN,
            ltout => \ADC_VDC.n31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_4_lut_adj_36_LC_10_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111111100"
        )
    port map (
            in0 => \N__28285\,
            in1 => \N__34589\,
            in2 => \N__26335\,
            in3 => \N__34299\,
            lcout => \ADC_VDC.n20514\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.adc_state_1__bdd_4_lut_4_lut_LC_10_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010110001101100"
        )
    port map (
            in0 => \N__34771\,
            in1 => \N__34120\,
            in2 => \N__34630\,
            in3 => \N__26307\,
            lcout => OPEN,
            ltout => \ADC_VDC.n21925_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.n21925_bdd_4_lut_4_lut_LC_10_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010011110100"
        )
    port map (
            in0 => \N__34593\,
            in1 => \N__30649\,
            in2 => \N__26332\,
            in3 => \N__34772\,
            lcout => OPEN,
            ltout => \ADC_VDC.n21928_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.adc_state_i1_LC_10_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__26329\,
            in1 => \N__34594\,
            in2 => \N__26323\,
            in3 => \N__34355\,
            lcout => \ADC_VDC.adc_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32846\,
            ce => \N__26320\,
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_2_lut_3_lut_LC_10_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__32515\,
            in1 => \N__32551\,
            in2 => \_gnd_net_\,
            in3 => \N__30667\,
            lcout => OPEN,
            ltout => \ADC_VDC.n6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i4_4_lut_LC_10_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__32470\,
            in1 => \N__32641\,
            in2 => \N__26311\,
            in3 => \N__32599\,
            lcout => \ADC_VDC.n10519\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i3_LC_10_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__34259\,
            in1 => \N__26798\,
            in2 => \N__26389\,
            in3 => \N__26586\,
            lcout => cmd_rdadctmp_3_adj_1469,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32880\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_3_lut_4_lut_adj_40_LC_10_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110000000000"
        )
    port map (
            in0 => \N__34096\,
            in1 => \N__34257\,
            in2 => \N__34751\,
            in3 => \N__34503\,
            lcout => n12853,
            ltout => \n12853_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i1_LC_10_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__34258\,
            in1 => \N__26610\,
            in2 => \N__26296\,
            in3 => \N__26408\,
            lcout => cmd_rdadctmp_1_adj_1471,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32880\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i0_LC_10_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__26797\,
            in1 => \N__26609\,
            in2 => \N__34879\,
            in3 => \N__34260\,
            lcout => cmd_rdadctmp_0_adj_1472,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32880\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_4_lut_4_lut_4_lut_LC_10_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010100000"
        )
    port map (
            in0 => \N__34255\,
            in1 => \N__34723\,
            in2 => \N__34564\,
            in3 => \N__34094\,
            lcout => \ADC_VDC.n13060\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i4_LC_10_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__26585\,
            in1 => \N__26564\,
            in2 => \N__26836\,
            in3 => \N__34261\,
            lcout => cmd_rdadctmp_4_adj_1468,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32880\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_4_lut_adj_43_LC_10_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000011100000"
        )
    port map (
            in0 => \N__34256\,
            in1 => \N__34724\,
            in2 => \N__34565\,
            in3 => \N__34095\,
            lcout => \ADC_VDC.n12885\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i8_LC_10_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__26504\,
            in1 => \N__26532\,
            in2 => \N__26837\,
            in3 => \N__34262\,
            lcout => cmd_rdadctmp_8_adj_1464,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32880\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i17_LC_10_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__34303\,
            in1 => \N__26427\,
            in2 => \N__26879\,
            in3 => \N__26480\,
            lcout => cmd_rdadctmp_17_adj_1455,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32912\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i16_LC_10_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__26426\,
            in1 => \N__34306\,
            in2 => \N__26458\,
            in3 => \N__26842\,
            lcout => cmd_rdadctmp_16_adj_1456,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32912\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i2_LC_10_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__34304\,
            in1 => \N__26387\,
            in2 => \N__26880\,
            in3 => \N__26409\,
            lcout => cmd_rdadctmp_2_adj_1470,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32912\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i12_LC_10_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__26958\,
            in1 => \N__34305\,
            in2 => \N__26364\,
            in3 => \N__26841\,
            lcout => cmd_rdadctmp_12_adj_1460,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32912\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i11_LC_10_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__34302\,
            in1 => \N__26957\,
            in2 => \N__26878\,
            in3 => \N__26989\,
            lcout => cmd_rdadctmp_11_adj_1461,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32912\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i19078_2_lut_LC_10_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34584\,
            in2 => \_gnd_net_\,
            in3 => \N__34301\,
            lcout => OPEN,
            ltout => \ADC_VDC.n21673_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.SCLK_46_LC_10_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001011100010"
        )
    port map (
            in0 => \N__26931\,
            in1 => \N__30613\,
            in2 => \N__26941\,
            in3 => \N__34141\,
            lcout => \VDC_SCLK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32912\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadctmp_i20_LC_10_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__26768\,
            in1 => \N__26920\,
            in2 => \N__34393\,
            in3 => \N__26846\,
            lcout => cmd_rdadctmp_20_adj_1452,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32912\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i12_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__34567\,
            in1 => \N__28369\,
            in2 => \N__26727\,
            in3 => \N__26746\,
            lcout => buf_adcdata_vdc_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32871\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i11_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__28365\,
            in1 => \N__34571\,
            in2 => \N__26691\,
            in3 => \N__26710\,
            lcout => buf_adcdata_vdc_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32871\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i4_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__34568\,
            in1 => \N__28370\,
            in2 => \N__26674\,
            in3 => \N__51342\,
            lcout => buf_adcdata_vdc_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32871\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i9_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__28368\,
            in1 => \N__34573\,
            in2 => \N__35301\,
            in3 => \N__26659\,
            lcout => buf_adcdata_vdc_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32871\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i8_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__34570\,
            in1 => \N__28371\,
            in2 => \N__26628\,
            in3 => \N__26647\,
            lcout => buf_adcdata_vdc_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32871\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i7_LC_10_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__28367\,
            in1 => \N__34572\,
            in2 => \N__47898\,
            in3 => \N__27115\,
            lcout => buf_adcdata_vdc_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32871\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i6_LC_10_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__34569\,
            in1 => \N__27103\,
            in2 => \N__40881\,
            in3 => \N__28372\,
            lcout => buf_adcdata_vdc_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32871\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.ADC_DATA_i5_LC_10_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__28366\,
            in1 => \N__34574\,
            in2 => \N__27091\,
            in3 => \N__38319\,
            lcout => buf_adcdata_vdc_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32871\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_3_lut_4_lut_4_lut_LC_10_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010100010"
        )
    port map (
            in0 => \N__34385\,
            in1 => \N__34774\,
            in2 => \N__34642\,
            in3 => \N__34149\,
            lcout => \ADC_VDC.n13020\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i18765_3_lut_LC_10_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000010001"
        )
    port map (
            in0 => \N__27048\,
            in1 => \N__34624\,
            in2 => \_gnd_net_\,
            in3 => \N__27076\,
            lcout => OPEN,
            ltout => \ADC_VDC.n21106_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.cmd_rdadcbuf_i34_LC_10_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__34386\,
            in1 => \N__27067\,
            in2 => \N__27058\,
            in3 => \N__34150\,
            lcout => cmd_rdadcbuf_34,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32913\,
            ce => \N__27031\,
            sr => \_gnd_net_\
        );

    \ADC_VDC.i9_4_lut_LC_10_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__29202\,
            in1 => \N__28497\,
            in2 => \N__28516\,
            in3 => \N__28434\,
            lcout => \ADC_VDC.n21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i7_4_lut_LC_10_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29235\,
            in1 => \N__28530\,
            in2 => \N__29257\,
            in3 => \N__29220\,
            lcout => \ADC_VDC.n19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_3__i0_LC_10_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__27004\,
            in1 => \N__54086\,
            in2 => \_gnd_net_\,
            in3 => \N__36242\,
            lcout => comm_buf_3_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55088\,
            ce => \N__27259\,
            sr => \N__27250\
        );

    \comm_buf_3__i7_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54085\,
            in1 => \N__36898\,
            in2 => \_gnd_net_\,
            in3 => \N__27226\,
            lcout => comm_buf_3_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55088\,
            ce => \N__27259\,
            sr => \N__27250\
        );

    \comm_buf_3__i6_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__35798\,
            in1 => \N__54089\,
            in2 => \_gnd_net_\,
            in3 => \N__27208\,
            lcout => comm_buf_3_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55088\,
            ce => \N__27259\,
            sr => \N__27250\
        );

    \comm_buf_3__i5_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__54084\,
            in1 => \_gnd_net_\,
            in2 => \N__27190\,
            in3 => \N__37995\,
            lcout => comm_buf_3_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55088\,
            ce => \N__27259\,
            sr => \N__27250\
        );

    \comm_buf_3__i4_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__35640\,
            in1 => \N__54088\,
            in2 => \_gnd_net_\,
            in3 => \N__27175\,
            lcout => comm_buf_3_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55088\,
            ce => \N__27259\,
            sr => \N__27250\
        );

    \comm_buf_3__i3_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__54083\,
            in1 => \N__27157\,
            in2 => \_gnd_net_\,
            in3 => \N__35558\,
            lcout => comm_buf_3_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55088\,
            ce => \N__27259\,
            sr => \N__27250\
        );

    \comm_buf_3__i2_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__35441\,
            in1 => \N__54087\,
            in2 => \_gnd_net_\,
            in3 => \N__27148\,
            lcout => comm_buf_3_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55088\,
            ce => \N__27259\,
            sr => \N__27250\
        );

    \comm_buf_3__i1_LC_10_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__54082\,
            in1 => \N__35977\,
            in2 => \_gnd_net_\,
            in3 => \N__27133\,
            lcout => comm_buf_3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55088\,
            ce => \N__27259\,
            sr => \N__27250\
        );

    \i18988_2_lut_4_lut_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__50096\,
            in1 => \N__49539\,
            in2 => \N__49957\,
            in3 => \N__53530\,
            lcout => OPEN,
            ltout => \n21143_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19_4_lut_adj_293_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000011010101"
        )
    port map (
            in0 => \N__54079\,
            in1 => \N__51643\,
            in2 => \N__27118\,
            in3 => \N__51685\,
            lcout => OPEN,
            ltout => \n12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_294_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49914\,
            in2 => \N__27262\,
            in3 => \N__49869\,
            lcout => n12116,
            ltout => \n12116_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12359_2_lut_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27253\,
            in3 => \N__54701\,
            lcout => n14756,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_279_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__50095\,
            in1 => \N__53529\,
            in2 => \_gnd_net_\,
            in3 => \N__49947\,
            lcout => OPEN,
            ltout => \n25_adj_1592_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_288_LC_10_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__49538\,
            in1 => \N__46077\,
            in2 => \N__27238\,
            in3 => \N__51642\,
            lcout => OPEN,
            ltout => \n11944_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_289_LC_10_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__46429\,
            in1 => \N__49870\,
            in2 => \N__27235\,
            in3 => \N__37515\,
            lcout => n11941,
            ltout => \n11941_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12338_2_lut_LC_10_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__27232\,
            in3 => \N__54700\,
            lcout => n14735,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19331_LC_10_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001100100"
        )
    port map (
            in0 => \N__57408\,
            in1 => \N__56797\,
            in2 => \N__41926\,
            in3 => \N__32100\,
            lcout => OPEN,
            ltout => \n21919_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n21919_bdd_4_lut_LC_10_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011000010"
        )
    port map (
            in0 => \N__38175\,
            in1 => \N__57409\,
            in2 => \N__27229\,
            in3 => \N__38623\,
            lcout => n21922,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18199_3_lut_LC_10_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__31176\,
            in1 => \N__56798\,
            in2 => \_gnd_net_\,
            in3 => \N__47274\,
            lcout => OPEN,
            ltout => \n20794_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18201_4_lut_LC_10_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011110000"
        )
    port map (
            in0 => \N__56800\,
            in1 => \N__27373\,
            in2 => \N__27358\,
            in3 => \N__57410\,
            lcout => OPEN,
            ltout => \n20796_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_2__bdd_4_lut_LC_10_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110001000"
        )
    port map (
            in0 => \N__56308\,
            in1 => \N__27355\,
            in2 => \N__27349\,
            in3 => \N__47694\,
            lcout => OPEN,
            ltout => \n22213_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22213_bdd_4_lut_LC_10_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101100"
        )
    port map (
            in0 => \N__27346\,
            in1 => \N__30157\,
            in2 => \N__27334\,
            in3 => \N__56309\,
            lcout => OPEN,
            ltout => \n22216_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_0__i2_LC_10_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54101\,
            in2 => \N__27331\,
            in3 => \N__35450\,
            lcout => comm_buf_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55105\,
            ce => \N__27505\,
            sr => \N__27454\
        );

    \i19000_4_lut_4_lut_LC_10_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101011101111"
        )
    port map (
            in0 => \N__56799\,
            in1 => \N__47508\,
            in2 => \N__56342\,
            in3 => \N__57407\,
            lcout => n21071,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19336_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__27328\,
            in1 => \N__47578\,
            in2 => \N__27313\,
            in3 => \N__57462\,
            lcout => OPEN,
            ltout => \n21907_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n21907_bdd_4_lut_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__47579\,
            in1 => \N__28174\,
            in2 => \N__27304\,
            in3 => \N__45067\,
            lcout => n21910,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19418_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__29715\,
            in1 => \N__57463\,
            in2 => \N__27300\,
            in3 => \N__56638\,
            lcout => OPEN,
            ltout => \n22033_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22033_bdd_4_lut_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__57464\,
            in1 => \N__32310\,
            in2 => \N__27265\,
            in3 => \N__29393\,
            lcout => OPEN,
            ltout => \n22036_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18228_3_lut_LC_10_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47580\,
            in2 => \N__27544\,
            in3 => \N__27541\,
            lcout => OPEN,
            ltout => \n20823_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1537450_i1_3_lut_LC_10_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27529\,
            in2 => \N__27523\,
            in3 => \N__56274\,
            lcout => OPEN,
            ltout => \n30_adj_1514_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_0__i5_LC_10_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__38022\,
            in1 => \_gnd_net_\,
            in2 => \N__27520\,
            in3 => \N__54100\,
            lcout => comm_buf_0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55116\,
            ce => \N__27513\,
            sr => \N__27464\
        );

    \CLK_DDS.tmp_buf_i10_LC_10_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__28795\,
            in1 => \N__28947\,
            in2 => \N__27628\,
            in3 => \N__30187\,
            lcout => \CLK_DDS.tmp_buf_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55125\,
            ce => \N__28551\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i11_LC_10_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__29556\,
            in1 => \N__28954\,
            in2 => \N__27418\,
            in3 => \N__28799\,
            lcout => \CLK_DDS.tmp_buf_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55125\,
            ce => \N__28551\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i12_LC_10_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__28796\,
            in1 => \N__27588\,
            in2 => \N__27409\,
            in3 => \N__28950\,
            lcout => \CLK_DDS.tmp_buf_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55125\,
            ce => \N__28551\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i13_LC_10_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__28951\,
            in1 => \N__28800\,
            in2 => \N__27400\,
            in3 => \N__29401\,
            lcout => \CLK_DDS.tmp_buf_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55125\,
            ce => \N__28551\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i14_LC_10_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__28797\,
            in1 => \N__28948\,
            in2 => \N__27391\,
            in3 => \N__27608\,
            lcout => \CLK_DDS.tmp_buf_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55125\,
            ce => \N__28551\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i15_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__28952\,
            in1 => \N__28801\,
            in2 => \N__27382\,
            in3 => \N__27920\,
            lcout => tmp_buf_15_adj_1448,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55125\,
            ce => \N__28551\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i9_LC_10_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__28798\,
            in1 => \N__28949\,
            in2 => \N__27570\,
            in3 => \N__27619\,
            lcout => \CLK_DDS.tmp_buf_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55125\,
            ce => \N__28551\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i8_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__28953\,
            in1 => \N__28802\,
            in2 => \N__27640\,
            in3 => \N__27964\,
            lcout => \CLK_DDS.tmp_buf_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55125\,
            ce => \N__28551\,
            sr => \_gnd_net_\
        );

    \buf_dds1_i14_LC_10_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__46017\,
            in1 => \N__40786\,
            in2 => \N__45914\,
            in3 => \N__27609\,
            lcout => buf_dds1_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55137\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i12_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__27589\,
            in1 => \N__45901\,
            in2 => \N__46708\,
            in3 => \N__46016\,
            lcout => buf_dds1_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55137\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i15_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__46018\,
            in1 => \N__30814\,
            in2 => \N__45915\,
            in3 => \N__27921\,
            lcout => buf_dds1_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55137\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i11_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__29555\,
            in1 => \N__45900\,
            in2 => \N__43806\,
            in3 => \N__46015\,
            lcout => buf_dds1_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55137\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \trig_dds1_305_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110000001100100"
        )
    port map (
            in0 => \N__52169\,
            in1 => \N__54699\,
            in2 => \N__28654\,
            in3 => \N__45937\,
            lcout => trig_dds1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55137\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i9_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__46019\,
            in1 => \N__44085\,
            in2 => \N__45916\,
            in3 => \N__27566\,
            lcout => buf_dds1_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55137\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_stop_328_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__44084\,
            in1 => \N__29887\,
            in2 => \_gnd_net_\,
            in3 => \N__38935\,
            lcout => eis_stop,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55137\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i0_LC_10_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__28974\,
            in1 => \N__28804\,
            in2 => \N__27730\,
            in3 => \N__27826\,
            lcout => \CLK_DDS.tmp_buf_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55150\,
            ce => \N__28555\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i1_LC_10_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__28803\,
            in1 => \N__28978\,
            in2 => \N__27706\,
            in3 => \N__31933\,
            lcout => \CLK_DDS.tmp_buf_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55150\,
            ce => \N__28555\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i2_LC_10_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__28975\,
            in1 => \N__28805\,
            in2 => \N__27697\,
            in3 => \N__32017\,
            lcout => \CLK_DDS.tmp_buf_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55150\,
            ce => \N__28555\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i3_LC_10_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__31828\,
            in1 => \N__28979\,
            in2 => \N__27688\,
            in3 => \N__28810\,
            lcout => \CLK_DDS.tmp_buf_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55150\,
            ce => \N__28555\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i4_LC_10_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__28976\,
            in1 => \N__28806\,
            in2 => \N__27679\,
            in3 => \N__36143\,
            lcout => \CLK_DDS.tmp_buf_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55150\,
            ce => \N__28555\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i5_LC_10_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__28980\,
            in1 => \N__28808\,
            in2 => \N__27667\,
            in3 => \N__29508\,
            lcout => \CLK_DDS.tmp_buf_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55150\,
            ce => \N__28555\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i6_LC_10_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__28977\,
            in1 => \N__28807\,
            in2 => \N__27658\,
            in3 => \N__36115\,
            lcout => \CLK_DDS.tmp_buf_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55150\,
            ce => \N__28555\,
            sr => \_gnd_net_\
        );

    \CLK_DDS.tmp_buf_i7_LC_10_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__28981\,
            in1 => \N__28809\,
            in2 => \N__27649\,
            in3 => \N__42544\,
            lcout => \CLK_DDS.tmp_buf_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55150\,
            ce => \N__28555\,
            sr => \_gnd_net_\
        );

    \buf_dds0_i3_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__45692\,
            in1 => \N__36397\,
            in2 => \N__52172\,
            in3 => \N__36717\,
            lcout => buf_dds0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55165\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i14_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__32258\,
            in1 => \_gnd_net_\,
            in2 => \N__41545\,
            in3 => \N__45691\,
            lcout => buf_dds0_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55165\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i0_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__39330\,
            in1 => \N__41356\,
            in2 => \N__52171\,
            in3 => \N__35856\,
            lcout => \acadc_skipCount_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55165\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i13_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__44846\,
            in1 => \N__39329\,
            in2 => \_gnd_net_\,
            in3 => \N__30205\,
            lcout => \acadc_skipCount_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55165\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22045_bdd_4_lut_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__27922\,
            in1 => \N__27901\,
            in2 => \N__45595\,
            in3 => \N__57502\,
            lcout => n22048,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i7_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__41544\,
            in1 => \N__39219\,
            in2 => \_gnd_net_\,
            in3 => \N__27857\,
            lcout => \VAC_FLT0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55165\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_0_i16_3_lut_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__27824\,
            in1 => \N__40374\,
            in2 => \_gnd_net_\,
            in3 => \N__56921\,
            lcout => n16_adj_1480,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i0_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__45840\,
            in1 => \N__27825\,
            in2 => \N__41364\,
            in3 => \N__46020\,
            lcout => buf_dds1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55165\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i8_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__27963\,
            in1 => \N__45911\,
            in2 => \N__43533\,
            in3 => \N__46021\,
            lcout => buf_dds1_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19511_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__28013\,
            in1 => \N__56913\,
            in2 => \N__27801\,
            in3 => \N__57489\,
            lcout => n22147,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i26_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__27746\,
            in1 => \N__50883\,
            in2 => \N__27778\,
            in3 => \N__50479\,
            lcout => cmd_rdadctmp_26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i9_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__52112\,
            in1 => \N__32337\,
            in2 => \N__44148\,
            in3 => \N__45673\,
            lcout => buf_dds0_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55180\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_5_i23_3_lut_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__30045\,
            in1 => \N__56914\,
            in2 => \_gnd_net_\,
            in3 => \N__30204\,
            lcout => n23_adj_1513,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i20_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__48953\,
            in1 => \N__50948\,
            in2 => \N__28162\,
            in3 => \N__28121\,
            lcout => buf_adcdata_iac_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55195\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i4_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__52108\,
            in1 => \N__39240\,
            in2 => \N__28086\,
            in3 => \N__43817\,
            lcout => \IAC_FLT1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55195\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i2_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__39238\,
            in1 => \N__52109\,
            in2 => \N__44149\,
            in3 => \N__28046\,
            lcout => \IAC_OSR1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55195\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i13_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__44850\,
            in1 => \N__32300\,
            in2 => \_gnd_net_\,
            in3 => \N__45677\,
            lcout => buf_dds0_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55195\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i3_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__39239\,
            in1 => \N__52110\,
            in2 => \N__38733\,
            in3 => \N__28014\,
            lcout => \IAC_FLT0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55195\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_0__bdd_4_lut_19551_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__28211\,
            in1 => \N__57541\,
            in2 => \N__27992\,
            in3 => \N__56967\,
            lcout => OPEN,
            ltout => \n22189_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22189_bdd_4_lut_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__57542\,
            in1 => \N__27959\,
            in2 => \N__27943\,
            in3 => \N__43413\,
            lcout => n20769,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_5_i16_3_lut_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__29509\,
            in1 => \N__43066\,
            in2 => \_gnd_net_\,
            in3 => \N__56968\,
            lcout => n16_adj_1489,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i1_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__52162\,
            in1 => \N__39241\,
            in2 => \N__43534\,
            in3 => \N__28212\,
            lcout => \IAC_OSR0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55209\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.t0off_i0_LC_11_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30349\,
            in2 => \_gnd_net_\,
            in3 => \N__28195\,
            lcout => \ADC_VDC.genclk.t0off_0\,
            ltout => OPEN,
            carryin => \bfn_11_3_0_\,
            carryout => \ADC_VDC.genclk.n19410\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__30532\,
            sr => \N__37444\
        );

    \ADC_VDC.genclk.t0off_i1_LC_11_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30379\,
            in2 => \N__52809\,
            in3 => \N__28192\,
            lcout => \ADC_VDC.genclk.t0off_1\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19410\,
            carryout => \ADC_VDC.genclk.n19411\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__30532\,
            sr => \N__37444\
        );

    \ADC_VDC.genclk.t0off_i2_LC_11_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52754\,
            in2 => \N__30322\,
            in3 => \N__28189\,
            lcout => \ADC_VDC.genclk.t0off_2\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19411\,
            carryout => \ADC_VDC.genclk.n19412\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__30532\,
            sr => \N__37444\
        );

    \ADC_VDC.genclk.t0off_i3_LC_11_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30232\,
            in2 => \N__52810\,
            in3 => \N__28186\,
            lcout => \ADC_VDC.genclk.t0off_3\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19412\,
            carryout => \ADC_VDC.genclk.n19413\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__30532\,
            sr => \N__37444\
        );

    \ADC_VDC.genclk.t0off_i4_LC_11_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52758\,
            in2 => \N__30367\,
            in3 => \N__28183\,
            lcout => \ADC_VDC.genclk.t0off_4\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19413\,
            carryout => \ADC_VDC.genclk.n19414\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__30532\,
            sr => \N__37444\
        );

    \ADC_VDC.genclk.t0off_i5_LC_11_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30246\,
            in2 => \N__52811\,
            in3 => \N__28180\,
            lcout => \ADC_VDC.genclk.t0off_5\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19414\,
            carryout => \ADC_VDC.genclk.n19415\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__30532\,
            sr => \N__37444\
        );

    \ADC_VDC.genclk.t0off_i6_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52762\,
            in2 => \N__30394\,
            in3 => \N__28177\,
            lcout => \ADC_VDC.genclk.t0off_6\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19415\,
            carryout => \ADC_VDC.genclk.n19416\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__30532\,
            sr => \N__37444\
        );

    \ADC_VDC.genclk.t0off_i7_LC_11_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30306\,
            in2 => \N__52812\,
            in3 => \N__28264\,
            lcout => \ADC_VDC.genclk.t0off_7\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19416\,
            carryout => \ADC_VDC.genclk.n19417\,
            clk => \INVADC_VDC.genclk.t0off_i0C_net\,
            ce => \N__30532\,
            sr => \N__37444\
        );

    \ADC_VDC.genclk.t0off_i8_LC_11_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30259\,
            in2 => \N__52750\,
            in3 => \N__28261\,
            lcout => \ADC_VDC.genclk.t0off_8\,
            ltout => OPEN,
            carryin => \bfn_11_4_0_\,
            carryout => \ADC_VDC.genclk.n19418\,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__30528\,
            sr => \N__37445\
        );

    \ADC_VDC.genclk.t0off_i9_LC_11_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52667\,
            in2 => \N__30583\,
            in3 => \N__28258\,
            lcout => \ADC_VDC.genclk.t0off_9\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19418\,
            carryout => \ADC_VDC.genclk.n19419\,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__30528\,
            sr => \N__37445\
        );

    \ADC_VDC.genclk.t0off_i10_LC_11_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30292\,
            in2 => \N__52747\,
            in3 => \N__28255\,
            lcout => \ADC_VDC.genclk.t0off_10\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19419\,
            carryout => \ADC_VDC.genclk.n19420\,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__30528\,
            sr => \N__37445\
        );

    \ADC_VDC.genclk.t0off_i11_LC_11_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52655\,
            in2 => \N__30553\,
            in3 => \N__28252\,
            lcout => \ADC_VDC.genclk.t0off_11\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19420\,
            carryout => \ADC_VDC.genclk.n19421\,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__30528\,
            sr => \N__37445\
        );

    \ADC_VDC.genclk.t0off_i12_LC_11_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30334\,
            in2 => \N__52748\,
            in3 => \N__28249\,
            lcout => \ADC_VDC.genclk.t0off_12\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19421\,
            carryout => \ADC_VDC.genclk.n19422\,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__30528\,
            sr => \N__37445\
        );

    \ADC_VDC.genclk.t0off_i13_LC_11_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52659\,
            in2 => \N__30274\,
            in3 => \N__28246\,
            lcout => \ADC_VDC.genclk.t0off_13\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19422\,
            carryout => \ADC_VDC.genclk.n19423\,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__30528\,
            sr => \N__37445\
        );

    \ADC_VDC.genclk.t0off_i14_LC_11_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30595\,
            in2 => \N__52749\,
            in3 => \N__28243\,
            lcout => \ADC_VDC.genclk.t0off_14\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19423\,
            carryout => \ADC_VDC.genclk.n19424\,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__30528\,
            sr => \N__37445\
        );

    \ADC_VDC.genclk.t0off_i15_LC_11_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__30567\,
            in1 => \N__52663\,
            in2 => \_gnd_net_\,
            in3 => \N__28240\,
            lcout => \ADC_VDC.genclk.t0off_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADC_VDC.genclk.t0off_i8C_net\,
            ce => \N__30528\,
            sr => \N__37445\
        );

    \ADC_VDC.i1_3_lut_4_lut_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001000"
        )
    port map (
            in0 => \N__34290\,
            in1 => \N__34742\,
            in2 => \N__34147\,
            in3 => \N__34490\,
            lcout => n13073,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.adc_state_i3_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010010000001100"
        )
    port map (
            in0 => \N__34113\,
            in1 => \N__34292\,
            in2 => \N__34562\,
            in3 => \N__34745\,
            lcout => adc_state_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32861\,
            ce => \N__30508\,
            sr => \_gnd_net_\
        );

    \ADC_VDC.i12542_2_lut_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29134\,
            in2 => \_gnd_net_\,
            in3 => \N__34289\,
            lcout => \ADC_VDC.n14900\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_2_lut_adj_31_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__34291\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34489\,
            lcout => OPEN,
            ltout => \ADC_VDC.n20618_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_4_lut_adj_38_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011001100"
        )
    port map (
            in0 => \N__34112\,
            in1 => \N__30475\,
            in2 => \N__28300\,
            in3 => \N__30469\,
            lcout => \ADC_VDC.n47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.adc_state_i0_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001011110"
        )
    port map (
            in0 => \N__34300\,
            in1 => \N__34844\,
            in2 => \N__34563\,
            in3 => \N__34716\,
            lcout => \ADC_VDC.adc_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32873\,
            ce => \N__28297\,
            sr => \_gnd_net_\
        );

    \ADC_VDC.i15997_3_lut_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001011010"
        )
    port map (
            in0 => \N__34845\,
            in1 => \_gnd_net_\,
            in2 => \N__34746\,
            in3 => \N__34151\,
            lcout => \ADC_VDC.n12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_2_lut_adj_30_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34712\,
            in2 => \_gnd_net_\,
            in3 => \N__34122\,
            lcout => \ADC_VDC.n7_adj_1403\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i18107_2_lut_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__34846\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34152\,
            lcout => \ADC_VDC.n20702\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i8_4_lut_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__28464\,
            in1 => \N__29271\,
            in2 => \N__28483\,
            in3 => \N__28449\,
            lcout => \ADC_VDC.n20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CLK_DDS.i19065_4_lut_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100111001100"
        )
    port map (
            in0 => \N__28909\,
            in1 => \N__28774\,
            in2 => \N__28664\,
            in3 => \N__28621\,
            lcout => \CLK_DDS.n12722\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.avg_cnt_i0_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28531\,
            in2 => \_gnd_net_\,
            in3 => \N__28519\,
            lcout => \ADC_VDC.avg_cnt_0\,
            ltout => OPEN,
            carryin => \bfn_11_7_0_\,
            carryout => \ADC_VDC.n19399\,
            clk => \N__32895\,
            ce => \N__29178\,
            sr => \N__29095\
        );

    \ADC_VDC.avg_cnt_i1_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28515\,
            in2 => \_gnd_net_\,
            in3 => \N__28501\,
            lcout => \ADC_VDC.avg_cnt_1\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19399\,
            carryout => \ADC_VDC.n19400\,
            clk => \N__32895\,
            ce => \N__29178\,
            sr => \N__29095\
        );

    \ADC_VDC.avg_cnt_i2_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28498\,
            in2 => \_gnd_net_\,
            in3 => \N__28486\,
            lcout => \ADC_VDC.avg_cnt_2\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19400\,
            carryout => \ADC_VDC.n19401\,
            clk => \N__32895\,
            ce => \N__29178\,
            sr => \N__29095\
        );

    \ADC_VDC.avg_cnt_i3_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28482\,
            in2 => \_gnd_net_\,
            in3 => \N__28468\,
            lcout => \ADC_VDC.avg_cnt_3\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19401\,
            carryout => \ADC_VDC.n19402\,
            clk => \N__32895\,
            ce => \N__29178\,
            sr => \N__29095\
        );

    \ADC_VDC.avg_cnt_i4_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28465\,
            in2 => \_gnd_net_\,
            in3 => \N__28453\,
            lcout => \ADC_VDC.avg_cnt_4\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19402\,
            carryout => \ADC_VDC.n19403\,
            clk => \N__32895\,
            ce => \N__29178\,
            sr => \N__29095\
        );

    \ADC_VDC.avg_cnt_i5_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28450\,
            in2 => \_gnd_net_\,
            in3 => \N__28438\,
            lcout => \ADC_VDC.avg_cnt_5\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19403\,
            carryout => \ADC_VDC.n19404\,
            clk => \N__32895\,
            ce => \N__29178\,
            sr => \N__29095\
        );

    \ADC_VDC.avg_cnt_i6_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28435\,
            in2 => \_gnd_net_\,
            in3 => \N__28423\,
            lcout => \ADC_VDC.avg_cnt_6\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19404\,
            carryout => \ADC_VDC.n19405\,
            clk => \N__32895\,
            ce => \N__29178\,
            sr => \N__29095\
        );

    \ADC_VDC.avg_cnt_i7_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29272\,
            in2 => \_gnd_net_\,
            in3 => \N__29260\,
            lcout => \ADC_VDC.avg_cnt_7\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19405\,
            carryout => \ADC_VDC.n19406\,
            clk => \N__32895\,
            ce => \N__29178\,
            sr => \N__29095\
        );

    \ADC_VDC.avg_cnt_i8_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29253\,
            in2 => \_gnd_net_\,
            in3 => \N__29239\,
            lcout => \ADC_VDC.avg_cnt_8\,
            ltout => OPEN,
            carryin => \bfn_11_8_0_\,
            carryout => \ADC_VDC.n19407\,
            clk => \N__32893\,
            ce => \N__29177\,
            sr => \N__29099\
        );

    \ADC_VDC.avg_cnt_i9_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29236\,
            in2 => \_gnd_net_\,
            in3 => \N__29224\,
            lcout => \ADC_VDC.avg_cnt_9\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19407\,
            carryout => \ADC_VDC.n19408\,
            clk => \N__32893\,
            ce => \N__29177\,
            sr => \N__29099\
        );

    \ADC_VDC.avg_cnt_i10_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29221\,
            in2 => \_gnd_net_\,
            in3 => \N__29209\,
            lcout => \ADC_VDC.avg_cnt_10\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19408\,
            carryout => \ADC_VDC.n19409\,
            clk => \N__32893\,
            ce => \N__29177\,
            sr => \N__29099\
        );

    \ADC_VDC.avg_cnt_i11_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29203\,
            in2 => \_gnd_net_\,
            in3 => \N__29206\,
            lcout => \ADC_VDC.avg_cnt_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32893\,
            ce => \N__29177\,
            sr => \N__29099\
        );

    \mux_128_Mux_7_i23_3_lut_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__29356\,
            in1 => \N__56956\,
            in2 => \_gnd_net_\,
            in3 => \N__36598\,
            lcout => OPEN,
            ltout => \n23_adj_1510_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18238_4_lut_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__56957\,
            in1 => \N__57393\,
            in2 => \N__29035\,
            in3 => \N__41692\,
            lcout => n20833,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18215_4_lut_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010001000"
        )
    port map (
            in0 => \N__57392\,
            in1 => \N__29017\,
            in2 => \N__31150\,
            in3 => \N__56958\,
            lcout => n20810,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i7_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29377\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => buf_control_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55084\,
            ce => \N__29344\,
            sr => \N__40641\
        );

    \i18851_2_lut_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__57394\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51286\,
            lcout => OPEN,
            ltout => \n21050_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18824_4_lut_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__54674\,
            in1 => \N__47696\,
            in2 => \N__29347\,
            in3 => \N__56169\,
            lcout => n21049,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_81_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__54672\,
            in1 => \N__51285\,
            in2 => \_gnd_net_\,
            in3 => \N__54080\,
            lcout => n20081,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_287_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000001000"
        )
    port map (
            in0 => \N__54081\,
            in1 => \N__49236\,
            in2 => \N__40621\,
            in3 => \N__54673\,
            lcout => n11905,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_150_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__53509\,
            in1 => \N__44400\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n10508,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i6_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__41527\,
            in1 => \N__45310\,
            in2 => \_gnd_net_\,
            in3 => \N__29296\,
            lcout => \buf_cfgRTD_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55089\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15009_2_lut_3_lut_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000000"
        )
    port map (
            in0 => \N__29421\,
            in1 => \_gnd_net_\,
            in2 => \N__29437\,
            in3 => \N__29448\,
            lcout => \comm_state_3_N_428_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_245_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010001000"
        )
    port map (
            in0 => \N__54656\,
            in1 => \N__49237\,
            in2 => \N__51297\,
            in3 => \N__44356\,
            lcout => n11882,
            ltout => \n11882_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i4_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__35662\,
            in1 => \N__30989\,
            in2 => \N__29275\,
            in3 => \N__29449\,
            lcout => comm_cmd_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55089\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_302_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__29447\,
            in1 => \N__29420\,
            in2 => \_gnd_net_\,
            in3 => \N__29432\,
            lcout => n20602,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i6_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__29436\,
            in1 => \N__30990\,
            in2 => \N__35811\,
            in3 => \N__30928\,
            lcout => comm_cmd_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55089\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i2_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__30999\,
            in1 => \N__30929\,
            in2 => \N__47701\,
            in3 => \N__35449\,
            lcout => comm_cmd_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55097\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i5_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__30930\,
            in1 => \N__31000\,
            in2 => \N__38023\,
            in3 => \N__29422\,
            lcout => comm_cmd_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55097\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_3_lut_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51293\,
            in2 => \N__53531\,
            in3 => \N__46588\,
            lcout => OPEN,
            ltout => \n8_adj_1522_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_237_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010000000"
        )
    port map (
            in0 => \N__29482\,
            in1 => \N__49238\,
            in2 => \N__29407\,
            in3 => \N__54657\,
            lcout => n12214,
            ltout => \n12214_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i2_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__54659\,
            in1 => \N__35448\,
            in2 => \N__29404\,
            in3 => \N__35082\,
            lcout => comm_buf_6_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55097\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i3_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__33075\,
            in1 => \N__54661\,
            in2 => \N__35568\,
            in3 => \N__29471\,
            lcout => comm_buf_6_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55097\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i13_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010111001100"
        )
    port map (
            in0 => \N__54658\,
            in1 => \N__29397\,
            in2 => \N__44851\,
            in3 => \N__45912\,
            lcout => buf_dds1_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55097\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i1_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__47172\,
            in1 => \N__54660\,
            in2 => \N__35978\,
            in3 => \N__29470\,
            lcout => comm_buf_6_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55097\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22075_bdd_4_lut_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__29557\,
            in1 => \N__29536\,
            in2 => \N__43104\,
            in3 => \N__57441\,
            lcout => n22078,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i5_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001110101010"
        )
    port map (
            in0 => \N__29498\,
            in1 => \N__54665\,
            in2 => \N__50137\,
            in3 => \N__45891\,
            lcout => buf_dds1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55106\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i0_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__54662\,
            in1 => \N__36254\,
            in2 => \N__38076\,
            in3 => \N__29472\,
            lcout => comm_buf_6_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55106\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_adj_236_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50097\,
            in2 => \_gnd_net_\,
            in3 => \N__54094\,
            lcout => n7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i7_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__54664\,
            in1 => \N__36895\,
            in2 => \N__33960\,
            in3 => \N__29476\,
            lcout => comm_buf_6_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55106\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i6_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__29475\,
            in1 => \N__54667\,
            in2 => \N__33166\,
            in3 => \N__35806\,
            lcout => comm_buf_6_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55106\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i5_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__54663\,
            in1 => \N__38259\,
            in2 => \N__38016\,
            in3 => \N__29474\,
            lcout => comm_buf_6_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55106\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_6__i4_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__29473\,
            in1 => \N__46734\,
            in2 => \N__35663\,
            in3 => \N__54666\,
            lcout => comm_buf_6_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55106\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14137_4_lut_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111100010011"
        )
    port map (
            in0 => \N__31489\,
            in1 => \N__32155\,
            in2 => \N__30462\,
            in3 => \N__38899\,
            lcout => OPEN,
            ltout => \n16539_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_state_i0_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101000010001"
        )
    port map (
            in0 => \N__37582\,
            in1 => \N__32159\,
            in2 => \N__29650\,
            in3 => \N__31837\,
            lcout => eis_state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeis_state_i0C_net\,
            ce => \N__30406\,
            sr => \N__32099\
        );

    \i24_4_lut_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110111001100010"
        )
    port map (
            in0 => \N__37581\,
            in1 => \N__32158\,
            in2 => \N__39122\,
            in3 => \N__46976\,
            lcout => OPEN,
            ltout => \n17_adj_1601_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_state_i1_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011110010"
        )
    port map (
            in0 => \N__39106\,
            in1 => \N__37583\,
            in2 => \N__29647\,
            in3 => \N__29644\,
            lcout => eis_state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeis_state_i0C_net\,
            ce => \N__30406\,
            sr => \N__32099\
        );

    \i1_2_lut_adj_211_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30454\,
            in2 => \_gnd_net_\,
            in3 => \N__31488\,
            lcout => n16547,
            ltout => \n16547_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i34_3_lut_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__46975\,
            in1 => \_gnd_net_\,
            in2 => \N__29638\,
            in3 => \N__37580\,
            lcout => OPEN,
            ltout => \n13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_state_i2_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110001100100"
        )
    port map (
            in0 => \N__39105\,
            in1 => \N__32160\,
            in2 => \N__29635\,
            in3 => \N__37528\,
            lcout => \eis_end_N_716\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVeis_state_i0C_net\,
            ce => \N__30406\,
            sr => \N__32099\
        );

    \mux_129_Mux_6_i26_3_lut_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__56887\,
            in1 => \N__31222\,
            in2 => \_gnd_net_\,
            in3 => \N__47413\,
            lcout => n26_adj_1495,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19345_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__57522\,
            in1 => \N__29632\,
            in2 => \N__29620\,
            in3 => \N__47699\,
            lcout => OPEN,
            ltout => \n21937_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n21937_bdd_4_lut_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__47700\,
            in1 => \N__36088\,
            in2 => \N__29590\,
            in3 => \N__29587\,
            lcout => OPEN,
            ltout => \n21940_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1542274_i1_3_lut_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56273\,
            in2 => \N__29686\,
            in3 => \N__29656\,
            lcout => OPEN,
            ltout => \n30_adj_1490_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i6_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__54051\,
            in1 => \N__35812\,
            in2 => \N__29683\,
            in3 => \_gnd_net_\,
            lcout => comm_buf_1_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55126\,
            ce => \N__38557\,
            sr => \N__36791\
        );

    \buf_dds1_i4_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101010000000"
        )
    port map (
            in0 => \N__46006\,
            in1 => \N__46666\,
            in2 => \N__45913\,
            in3 => \N__36144\,
            lcout => buf_dds1_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55138\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i12_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__33857\,
            in1 => \N__42143\,
            in2 => \_gnd_net_\,
            in3 => \N__45657\,
            lcout => buf_dds0_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55138\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i10_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__30185\,
            in1 => \N__45896\,
            in2 => \N__38731\,
            in3 => \N__46005\,
            lcout => buf_dds1_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55138\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i8_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__39328\,
            in1 => \N__43520\,
            in2 => \N__52193\,
            in3 => \N__31533\,
            lcout => \acadc_skipCount_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55138\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19482_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__57521\,
            in1 => \N__29680\,
            in2 => \N__29674\,
            in3 => \N__47697\,
            lcout => OPEN,
            ltout => \n22111_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22111_bdd_4_lut_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__47698\,
            in1 => \N__31905\,
            in2 => \N__29659\,
            in3 => \N__41722\,
            lcout => n22114,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i6_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__31906\,
            in1 => \N__52177\,
            in2 => \N__51429\,
            in3 => \N__39327\,
            lcout => \acadc_skipCount_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55138\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_4_lut_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100011"
        )
    port map (
            in0 => \N__37593\,
            in1 => \N__32156\,
            in2 => \N__39151\,
            in3 => \N__32067\,
            lcout => n13443,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6372_3_lut_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__42596\,
            in1 => \N__42459\,
            in2 => \_gnd_net_\,
            in3 => \N__43295\,
            lcout => n8_adj_1536,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i5_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__44847\,
            in1 => \N__43871\,
            in2 => \_gnd_net_\,
            in3 => \N__30041\,
            lcout => \AMPV_POW\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55151\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19145_2_lut_3_lut_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__32068\,
            in1 => \N__39141\,
            in2 => \_gnd_net_\,
            in3 => \N__32180\,
            lcout => n20757,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.DTRIG_39_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000001000"
        )
    port map (
            in0 => \N__30022\,
            in1 => \N__29949\,
            in2 => \N__50952\,
            in3 => \N__31861\,
            lcout => acadc_dtrig_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55151\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_rst_327_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__32069\,
            in1 => \_gnd_net_\,
            in2 => \N__38730\,
            in3 => \N__29886\,
            lcout => acadc_rst,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55151\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.DTRIG_39_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000001000"
        )
    port map (
            in0 => \N__29863\,
            in1 => \N__29794\,
            in2 => \N__48335\,
            in3 => \N__31885\,
            lcout => acadc_dtrig_v,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55151\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_device_acadc_i6_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__44848\,
            in1 => \N__39205\,
            in2 => \_gnd_net_\,
            in3 => \N__29705\,
            lcout => \VAC_OSR1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55151\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_126_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__31884\,
            in1 => \N__31859\,
            in2 => \_gnd_net_\,
            in3 => \N__38898\,
            lcout => OPEN,
            ltout => \n4_adj_1473_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19069_4_lut_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001110111"
        )
    port map (
            in0 => \N__37595\,
            in1 => \N__39108\,
            in2 => \N__30208\,
            in3 => \N__32157\,
            lcout => n20529,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14975_2_lut_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31882\,
            in2 => \_gnd_net_\,
            in3 => \N__31858\,
            lcout => n17357,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_269_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__37594\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39107\,
            lcout => n35,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i10_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__52176\,
            in1 => \N__32366\,
            in2 => \N__38732\,
            in3 => \N__45656\,
            lcout => buf_dds0_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55166\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_61_i14_2_lut_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33700\,
            in2 => \_gnd_net_\,
            in3 => \N__30203\,
            lcout => n14_adj_1498,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__33676\,
            in1 => \N__36948\,
            in2 => \N__33634\,
            in3 => \N__36563\,
            lcout => n18_adj_1587,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22147_bdd_4_lut_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__30186\,
            in1 => \N__30163\,
            in2 => \N__32370\,
            in3 => \N__57531\,
            lcout => n22150,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18095_4_lut_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010101110"
        )
    port map (
            in0 => \N__32094\,
            in1 => \N__32161\,
            in2 => \N__39157\,
            in3 => \N__37603\,
            lcout => OPEN,
            ltout => \n20690_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_trig_300_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010000000100"
        )
    port map (
            in0 => \N__32163\,
            in1 => \N__39156\,
            in2 => \N__30145\,
            in3 => \N__30133\,
            lcout => acadc_trig,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVacadc_trig_300C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_end_299_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001011110000"
        )
    port map (
            in0 => \N__32164\,
            in1 => \N__32095\,
            in2 => \N__30099\,
            in3 => \N__30106\,
            lcout => eis_end,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVacadc_trig_300C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i24_4_lut_adj_234_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010101100"
        )
    port map (
            in0 => \N__30461\,
            in1 => \N__30415\,
            in2 => \N__37605\,
            in3 => \N__38941\,
            lcout => OPEN,
            ltout => \n11_adj_1620_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19112_3_lut_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111111111111"
        )
    port map (
            in0 => \N__32162\,
            in1 => \_gnd_net_\,
            in2 => \N__30409\,
            in3 => \N__39152\,
            lcout => n11730,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_187_i9_2_lut_3_lut_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__57540\,
            in1 => \N__56965\,
            in2 => \_gnd_net_\,
            in3 => \N__47695\,
            lcout => n9_adj_1407,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i19095_2_lut_LC_12_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34962\,
            in2 => \_gnd_net_\,
            in3 => \N__34930\,
            lcout => \ADC_VDC.genclk.n14695\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i19040_4_lut_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__30390\,
            in1 => \N__30378\,
            in2 => \N__30366\,
            in3 => \N__30348\,
            lcout => OPEN,
            ltout => \ADC_VDC.genclk.n21169_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i18722_4_lut_LC_12_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30538\,
            in1 => \N__30220\,
            in2 => \N__30337\,
            in3 => \N__30280\,
            lcout => \ADC_VDC.genclk.n21167\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i11_4_lut_LC_12_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30333\,
            in1 => \N__30318\,
            in2 => \N__30307\,
            in3 => \N__30291\,
            lcout => \ADC_VDC.genclk.n27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i10_4_lut_LC_12_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30270\,
            in1 => \N__30258\,
            in2 => \N__30247\,
            in3 => \N__30231\,
            lcout => \ADC_VDC.genclk.n26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i12_4_lut_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30594\,
            in1 => \N__30579\,
            in2 => \N__30568\,
            in3 => \N__30549\,
            lcout => \ADC_VDC.genclk.n28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i19072_2_lut_LC_12_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__34935\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34963\,
            lcout => \ADC_VDC.genclk.n11721\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i19088_4_lut_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010101010"
        )
    port map (
            in0 => \N__34294\,
            in1 => \N__34485\,
            in2 => \N__34877\,
            in3 => \N__30637\,
            lcout => \ADC_VDC.n4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i19137_4_lut_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110011011111"
        )
    port map (
            in0 => \N__30624\,
            in1 => \N__34487\,
            in2 => \N__34356\,
            in3 => \N__30754\,
            lcout => \ADC_VDC.n17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i7713_3_lut_4_lut_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001011011010"
        )
    port map (
            in0 => \N__34743\,
            in1 => \N__34158\,
            in2 => \N__34878\,
            in3 => \N__30772\,
            lcout => OPEN,
            ltout => \ADC_VDC.n10112_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_4_lut_4_lut_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101011111110"
        )
    port map (
            in0 => \N__34486\,
            in1 => \N__34295\,
            in2 => \N__30511\,
            in3 => \N__30625\,
            lcout => \ADC_VDC.n12793\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.adc_state_i2_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__34744\,
            in1 => \N__34488\,
            in2 => \_gnd_net_\,
            in3 => \N__34159\,
            lcout => adc_state_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32778\,
            ce => \N__30499\,
            sr => \N__30493\
        );

    \ADC_VDC.i1_4_lut_adj_37_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011111110"
        )
    port map (
            in0 => \N__30481\,
            in1 => \N__34293\,
            in2 => \N__34561\,
            in3 => \N__30623\,
            lcout => \ADC_VDC.n72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i18115_2_lut_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34741\,
            in2 => \_gnd_net_\,
            in3 => \N__30770\,
            lcout => \ADC_VDC.n20710\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i2_3_lut_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__32435\,
            in1 => \N__32930\,
            in2 => \_gnd_net_\,
            in3 => \N__32951\,
            lcout => \ADC_VDC.n20490\,
            ltout => \ADC_VDC.n20490_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_2_lut_adj_32_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__32509\,
            in1 => \_gnd_net_\,
            in2 => \N__30688\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \ADC_VDC.n11251_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i4_4_lut_adj_34_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__32463\,
            in1 => \N__32566\,
            in2 => \N__30685\,
            in3 => \N__32546\,
            lcout => \ADC_VDC.n15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i5_3_lut_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__32952\,
            in1 => \N__32931\,
            in2 => \_gnd_net_\,
            in3 => \N__30778\,
            lcout => OPEN,
            ltout => \ADC_VDC.n20523_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i18909_4_lut_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__32464\,
            in1 => \N__34307\,
            in2 => \N__30682\,
            in3 => \N__32632\,
            lcout => \ADC_VDC.n21178\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i18807_4_lut_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010000000"
        )
    port map (
            in0 => \N__30601\,
            in1 => \N__32465\,
            in2 => \N__34768\,
            in3 => \N__30663\,
            lcout => \ADC_VDC.n21025\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i18117_2_lut_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34865\,
            in2 => \_gnd_net_\,
            in3 => \N__30636\,
            lcout => \ADC_VDC.n20712\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i19071_4_lut_4_lut_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011101101"
        )
    port map (
            in0 => \N__34740\,
            in1 => \N__34368\,
            in2 => \N__34620\,
            in3 => \N__34157\,
            lcout => \ADC_VDC.n11662\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i18962_4_lut_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__32590\,
            in1 => \N__32542\,
            in2 => \N__32640\,
            in3 => \N__32505\,
            lcout => \ADC_VDC.n21028\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_137_Mux_7_i1_3_lut_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__30810\,
            in1 => \N__42624\,
            in2 => \_gnd_net_\,
            in3 => \N__51632\,
            lcout => n1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i4_4_lut_adj_35_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__32541\,
            in1 => \N__32589\,
            in2 => \N__32511\,
            in3 => \N__32436\,
            lcout => \ADC_VDC.n10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i40_3_lut_4_lut_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100100101"
        )
    port map (
            in0 => \N__34739\,
            in1 => \N__34156\,
            in2 => \N__34864\,
            in3 => \N__30771\,
            lcout => \ADC_VDC.n19_adj_1405\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \wdtick_cnt_3763_3764__i1_LC_12_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100010001"
        )
    port map (
            in0 => \N__30701\,
            in1 => \N__30740\,
            in2 => \_gnd_net_\,
            in3 => \N__30721\,
            lcout => wdtick_cnt_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40928\,
            ce => \N__33040\,
            sr => \N__40683\
        );

    \wdtick_cnt_3763_3764__i3_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101010100000"
        )
    port map (
            in0 => \N__30723\,
            in1 => \_gnd_net_\,
            in2 => \N__30745\,
            in3 => \N__30702\,
            lcout => wdtick_cnt_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40928\,
            ce => \N__33040\,
            sr => \N__40683\
        );

    \wdtick_cnt_3763_3764__i2_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30739\,
            in2 => \_gnd_net_\,
            in3 => \N__30722\,
            lcout => wdtick_cnt_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40928\,
            ce => \N__33040\,
            sr => \N__40683\
        );

    \wdtick_flag_289_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100010000"
        )
    port map (
            in0 => \N__30744\,
            in1 => \N__30724\,
            in2 => \N__30706\,
            in3 => \N__50256\,
            lcout => wdtick_flag,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__40938\,
            ce => 'H',
            sr => \N__40684\
        );

    \i1_2_lut_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__51209\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__54563\,
            lcout => n12205,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18699_2_lut_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__38202\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53462\,
            lcout => n20931,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i7_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__30932\,
            in1 => \N__30992\,
            in2 => \N__36897\,
            in3 => \N__49288\,
            lcout => comm_cmd_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55081\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_i3_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__56146\,
            in1 => \N__30991\,
            in2 => \N__35567\,
            in3 => \N__30931\,
            lcout => comm_cmd_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55081\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_278_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__53461\,
            in1 => \N__56144\,
            in2 => \_gnd_net_\,
            in3 => \N__38201\,
            lcout => n20622,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_0_i30_3_lut_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__30898\,
            in1 => \N__30883\,
            in2 => \_gnd_net_\,
            in3 => \N__56145\,
            lcout => n30_adj_1475,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_adj_120_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__54562\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51208\,
            lcout => n20627,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_4__i0_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__30871\,
            in1 => \N__53979\,
            in2 => \_gnd_net_\,
            in3 => \N__36252\,
            lcout => comm_buf_4_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55086\,
            ce => \N__49825\,
            sr => \N__33106\
        );

    \comm_buf_4__i7_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__53978\,
            in1 => \N__36881\,
            in2 => \_gnd_net_\,
            in3 => \N__30850\,
            lcout => comm_buf_4_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55086\,
            ce => \N__49825\,
            sr => \N__33106\
        );

    \comm_buf_4__i6_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35802\,
            in1 => \N__30832\,
            in2 => \_gnd_net_\,
            in3 => \N__53982\,
            lcout => comm_buf_4_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55086\,
            ce => \N__49825\,
            sr => \N__33106\
        );

    \comm_buf_4__i5_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__53977\,
            in1 => \N__38017\,
            in2 => \_gnd_net_\,
            in3 => \N__31123\,
            lcout => comm_buf_4_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55086\,
            ce => \N__49825\,
            sr => \N__33106\
        );

    \comm_buf_4__i4_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35664\,
            in1 => \N__31105\,
            in2 => \_gnd_net_\,
            in3 => \N__53981\,
            lcout => comm_buf_4_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55086\,
            ce => \N__49825\,
            sr => \N__33106\
        );

    \comm_buf_4__i3_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__53976\,
            in1 => \N__35559\,
            in2 => \_gnd_net_\,
            in3 => \N__31087\,
            lcout => comm_buf_4_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55086\,
            ce => \N__49825\,
            sr => \N__33106\
        );

    \comm_buf_4__i2_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35451\,
            in1 => \N__31069\,
            in2 => \_gnd_net_\,
            in3 => \N__53980\,
            lcout => comm_buf_4_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55086\,
            ce => \N__49825\,
            sr => \N__33106\
        );

    \comm_buf_4__i1_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__53975\,
            in1 => \N__35967\,
            in2 => \_gnd_net_\,
            in3 => \N__31048\,
            lcout => comm_buf_4_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55086\,
            ce => \N__49825\,
            sr => \N__33106\
        );

    \data_idxvec_i0_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__31027\,
            in1 => \N__35895\,
            in2 => \N__54711\,
            in3 => \N__31012\,
            lcout => data_idxvec_0,
            ltout => OPEN,
            carryin => \bfn_12_12_0_\,
            carryout => n19335,
            clk => \N__55094\,
            ce => \N__38581\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i1_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__38443\,
            in1 => \N__36039\,
            in2 => \N__54713\,
            in3 => \N__31009\,
            lcout => data_idxvec_1,
            ltout => OPEN,
            carryin => n19335,
            carryout => n19336,
            clk => \N__55094\,
            ce => \N__38581\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i2_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__41283\,
            in1 => \N__54645\,
            in2 => \N__33340\,
            in3 => \N__31006\,
            lcout => data_idxvec_2,
            ltout => OPEN,
            carryin => n19336,
            carryout => n19337,
            clk => \N__55094\,
            ce => \N__38581\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i3_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__38855\,
            in1 => \N__33390\,
            in2 => \N__54714\,
            in3 => \N__31003\,
            lcout => data_idxvec_3,
            ltout => OPEN,
            carryin => n19337,
            carryout => n19338,
            clk => \N__55094\,
            ce => \N__38581\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i4_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__38470\,
            in1 => \N__54649\,
            in2 => \N__33439\,
            in3 => \N__31228\,
            lcout => data_idxvec_4,
            ltout => OPEN,
            carryin => n19338,
            carryout => n19339,
            clk => \N__55094\,
            ce => \N__38581\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i5_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__50132\,
            in1 => \N__31287\,
            in2 => \N__54715\,
            in3 => \N__31225\,
            lcout => data_idxvec_5,
            ltout => OPEN,
            carryin => n19339,
            carryout => n19340,
            clk => \N__55094\,
            ce => \N__38581\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i6_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__51375\,
            in1 => \N__31221\,
            in2 => \N__54712\,
            in3 => \N__31207\,
            lcout => data_idxvec_6,
            ltout => OPEN,
            carryin => n19340,
            carryout => n19341,
            clk => \N__55094\,
            ce => \N__38581\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i7_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__41259\,
            in1 => \N__36678\,
            in2 => \N__54716\,
            in3 => \N__31204\,
            lcout => data_idxvec_7,
            ltout => OPEN,
            carryin => n19341,
            carryout => n19342,
            clk => \N__55094\,
            ce => \N__38581\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i8_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__41781\,
            in1 => \N__54576\,
            in2 => \N__41470\,
            in3 => \N__31201\,
            lcout => data_idxvec_8,
            ltout => OPEN,
            carryin => \bfn_12_13_0_\,
            carryout => n19343,
            clk => \N__55103\,
            ce => \N__38580\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i9_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__38143\,
            in1 => \N__31194\,
            in2 => \N__54693\,
            in3 => \N__31180\,
            lcout => data_idxvec_9,
            ltout => OPEN,
            carryin => n19343,
            carryout => n19344,
            clk => \N__55103\,
            ce => \N__38580\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i10_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__41943\,
            in1 => \N__54580\,
            in2 => \N__31177\,
            in3 => \N__31156\,
            lcout => data_idxvec_10,
            ltout => OPEN,
            carryin => n19344,
            carryout => n19345,
            clk => \N__55103\,
            ce => \N__38580\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i11_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__38590\,
            in1 => \N__44988\,
            in2 => \N__54694\,
            in3 => \N__31153\,
            lcout => data_idxvec_11,
            ltout => OPEN,
            carryin => n19345,
            carryout => n19346,
            clk => \N__55103\,
            ce => \N__38580\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i12_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__42126\,
            in1 => \N__54584\,
            in2 => \N__31146\,
            in3 => \N__31126\,
            lcout => data_idxvec_12,
            ltout => OPEN,
            carryin => n19346,
            carryout => n19347,
            clk => \N__55103\,
            ce => \N__38580\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i13_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__44849\,
            in1 => \N__31356\,
            in2 => \N__54695\,
            in3 => \N__31342\,
            lcout => data_idxvec_13,
            ltout => OPEN,
            carryin => n19347,
            carryout => n19348,
            clk => \N__55103\,
            ce => \N__38580\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i14_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__41526\,
            in1 => \N__54588\,
            in2 => \N__31332\,
            in3 => \N__31312\,
            lcout => data_idxvec_14,
            ltout => OPEN,
            carryin => n19348,
            carryout => n19349,
            clk => \N__55103\,
            ce => \N__38580\,
            sr => \_gnd_net_\
        );

    \data_idxvec_i15_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011000111100100"
        )
    port map (
            in0 => \N__54589\,
            in1 => \N__31302\,
            in2 => \N__45772\,
            in3 => \N__31309\,
            lcout => data_idxvec_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55103\,
            ce => \N__38580\,
            sr => \_gnd_net_\
        );

    \mux_129_Mux_5_i26_3_lut_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__56890\,
            in1 => \N__31288\,
            in2 => \_gnd_net_\,
            in3 => \N__46783\,
            lcout => OPEN,
            ltout => \n26_adj_1486_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19546_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010101010"
        )
    port map (
            in0 => \N__57523\,
            in1 => \N__31234\,
            in2 => \N__31273\,
            in3 => \N__47786\,
            lcout => OPEN,
            ltout => \n22177_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22177_bdd_4_lut_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__47787\,
            in1 => \N__38422\,
            in2 => \N__31270\,
            in3 => \N__31376\,
            lcout => OPEN,
            ltout => \n22180_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1542877_i1_3_lut_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31267\,
            in2 => \N__31255\,
            in3 => \N__56257\,
            lcout => OPEN,
            ltout => \n30_adj_1485_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i5_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__54095\,
            in1 => \N__38018\,
            in2 => \N__31252\,
            in3 => \_gnd_net_\,
            lcout => comm_buf_1_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55112\,
            ce => \N__38546\,
            sr => \N__36808\
        );

    \i18810_2_lut_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31249\,
            in2 => \_gnd_net_\,
            in3 => \N__56889\,
            lcout => n21036,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i3_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111000100010"
        )
    port map (
            in0 => \N__41797\,
            in1 => \N__54591\,
            in2 => \N__52194\,
            in3 => \N__36346\,
            lcout => data_index_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55123\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_354_Mux_0_i15_4_lut_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__54590\,
            in1 => \N__42874\,
            in2 => \N__52091\,
            in3 => \N__42859\,
            lcout => \data_index_9_N_212_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4_4_lut_adj_316_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__33610\,
            in1 => \N__33655\,
            in2 => \N__31381\,
            in3 => \N__33353\,
            lcout => OPEN,
            ltout => \n20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10_4_lut_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110110"
        )
    port map (
            in0 => \N__33733\,
            in1 => \N__31529\,
            in2 => \N__31513\,
            in3 => \N__31510\,
            lcout => OPEN,
            ltout => \n26_adj_1604_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15_4_lut_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31501\,
            in1 => \N__31891\,
            in2 => \N__31492\,
            in3 => \N__36271\,
            lcout => n31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_354_Mux_3_i15_4_lut_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__36345\,
            in1 => \N__54592\,
            in2 => \N__52092\,
            in3 => \N__41796\,
            lcout => \data_index_9_N_212_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i3_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__52181\,
            in1 => \N__39323\,
            in2 => \N__36396\,
            in3 => \N__33354\,
            lcout => \acadc_skipCount_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55123\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i5_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__31377\,
            in1 => \N__50181\,
            in2 => \N__39331\,
            in3 => \N__52185\,
            lcout => \acadc_skipCount_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55123\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19091_2_lut_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__33914\,
            in1 => \_gnd_net_\,
            in2 => \N__32185\,
            in3 => \_gnd_net_\,
            lcout => n14639,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_2_i16_3_lut_LC_12_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__32012\,
            in1 => \N__42753\,
            in2 => \_gnd_net_\,
            in3 => \N__56897\,
            lcout => n16_adj_1504,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i1_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100000000000"
        )
    port map (
            in0 => \N__45839\,
            in1 => \N__43382\,
            in2 => \N__31931\,
            in3 => \N__46013\,
            lcout => buf_dds1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55133\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_53_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__33492\,
            in1 => \N__31904\,
            in2 => \N__33754\,
            in3 => \N__35855\,
            lcout => n17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.i1_2_lut_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31883\,
            in2 => \_gnd_net_\,
            in3 => \N__31860\,
            lcout => \iac_raw_buf_N_728\,
            ltout => \iac_raw_buf_N_728_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \eis_state_1__bdd_4_lut_4_lut_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111010101010"
        )
    port map (
            in0 => \N__39137\,
            in1 => \N__32181\,
            in2 => \N__31840\,
            in3 => \N__37604\,
            lcout => n21997,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i3_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010011101110"
        )
    port map (
            in0 => \N__45838\,
            in1 => \N__31820\,
            in2 => \N__38869\,
            in3 => \N__54710\,
            lcout => buf_dds1_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55133\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_274_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__31804\,
            in1 => \N__52173\,
            in2 => \_gnd_net_\,
            in3 => \N__54596\,
            lcout => n12353,
            ltout => \n12353_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i1_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111101000000"
        )
    port map (
            in0 => \N__52175\,
            in1 => \N__43390\,
            in2 => \N__31792\,
            in3 => \N__32231\,
            lcout => buf_dds0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55145\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3787_3_lut_4_lut_4_lut_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__32070\,
            in1 => \N__32179\,
            in2 => \N__31789\,
            in3 => \N__46968\,
            lcout => \iac_raw_buf_N_726\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19122_4_lut_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000111"
        )
    port map (
            in0 => \N__32178\,
            in1 => \N__37602\,
            in2 => \N__32087\,
            in3 => \N__39142\,
            lcout => n11538,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18710_2_lut_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__56888\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32032\,
            lcout => n20949,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i0_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__52174\,
            in1 => \N__41355\,
            in2 => \N__40373\,
            in3 => \N__45655\,
            lcout => buf_dds0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55145\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i2_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__46014\,
            in1 => \N__32016\,
            in2 => \N__42823\,
            in3 => \N__45895\,
            lcout => buf_dds1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55145\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i7_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__39064\,
            in1 => \N__37138\,
            in2 => \N__55888\,
            in3 => \N__55622\,
            lcout => \SIG_DDS.tmp_buf_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55160\,
            ce => \N__40330\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.i12468_3_lut_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__55711\,
            in1 => \N__55873\,
            in2 => \_gnd_net_\,
            in3 => \N__55620\,
            lcout => n14869,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.i19105_4_lut_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011110"
        )
    port map (
            in0 => \N__55712\,
            in1 => \N__55874\,
            in2 => \N__53018\,
            in3 => \N__55621\,
            lcout => \SIG_DDS.n9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_7_i16_3_lut_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__42543\,
            in1 => \N__39063\,
            in2 => \_gnd_net_\,
            in3 => \N__56964\,
            lcout => OPEN,
            ltout => \n16_adj_1621_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n21961_bdd_4_lut_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__31986\,
            in1 => \N__31960\,
            in2 => \N__31948\,
            in3 => \N__47834\,
            lcout => n21964,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i10_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__55880\,
            in1 => \N__32371\,
            in2 => \N__32320\,
            in3 => \N__55662\,
            lcout => \SIG_DDS.tmp_buf_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55175\,
            ce => \N__40329\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i11_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__55663\,
            in1 => \N__55881\,
            in2 => \N__43108\,
            in3 => \N__32350\,
            lcout => \SIG_DDS.tmp_buf_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55175\,
            ce => \N__40329\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i9_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__55886\,
            in1 => \N__55668\,
            in2 => \N__32203\,
            in3 => \N__32344\,
            lcout => \SIG_DDS.tmp_buf_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55175\,
            ce => \N__40329\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i13_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__55664\,
            in1 => \N__55882\,
            in2 => \N__33838\,
            in3 => \N__32311\,
            lcout => \SIG_DDS.tmp_buf_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55175\,
            ce => \N__40329\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i14_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__55883\,
            in1 => \N__55665\,
            in2 => \N__32281\,
            in3 => \N__32271\,
            lcout => \SIG_DDS.tmp_buf_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55175\,
            ce => \N__40329\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i1_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__55666\,
            in1 => \N__55884\,
            in2 => \N__40342\,
            in3 => \N__32238\,
            lcout => \SIG_DDS.tmp_buf_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55175\,
            ce => \N__40329\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i8_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__55667\,
            in1 => \N__55885\,
            in2 => \N__32212\,
            in3 => \N__43417\,
            lcout => \SIG_DDS.tmp_buf_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55175\,
            ce => \N__40329\,
            sr => \_gnd_net_\
        );

    \comm_spi.i19174_4_lut_3_lut_LC_13_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__32194\,
            in1 => \N__32409\,
            in2 => \_gnd_net_\,
            in3 => \N__55464\,
            lcout => \comm_spi.n22629\,
            ltout => \comm_spi.n22629_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i12199_3_lut_LC_13_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__32401\,
            in1 => \_gnd_net_\,
            in2 => \N__32188\,
            in3 => \N__33802\,
            lcout => comm_rx_buf_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.t_clk_24_LC_13_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34931\,
            lcout => \VDC_CLK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADC_VDC.genclk.t_clk_24C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.div_state_i0_LC_13_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011111110110011"
        )
    port map (
            in0 => \N__32383\,
            in1 => \N__34970\,
            in2 => \N__34936\,
            in3 => \N__33781\,
            lcout => \ADC_VDC.genclk.div_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADC_VDC.genclk.t_clk_24C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i19159_4_lut_3_lut_LC_13_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__37346\,
            in1 => \N__33818\,
            in2 => \_gnd_net_\,
            in3 => \N__55463\,
            lcout => \comm_spi.n22632\,
            ltout => \comm_spi.n22632_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i12185_3_lut_LC_13_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__34995\,
            in1 => \_gnd_net_\,
            in2 => \N__32416\,
            in3 => \N__37424\,
            lcout => \comm_spi.imosi\,
            ltout => \comm_spi.imosi_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_86_2_lut_LC_13_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32413\,
            in3 => \N__55465\,
            lcout => \comm_spi.DOUT_7__N_738\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_87_2_lut_LC_13_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__32410\,
            in1 => \_gnd_net_\,
            in2 => \N__55473\,
            in3 => \_gnd_net_\,
            lcout => \comm_spi.DOUT_7__N_739\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_rx_i0_12197_12198_set_LC_13_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__37426\,
            in1 => \N__34994\,
            in2 => \_gnd_net_\,
            in3 => \N__33820\,
            lcout => \comm_spi.n14599\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52364\,
            ce => 'H',
            sr => \N__32395\
        );

    \ADC_VDC.genclk.div_state_1__I_0_1_lut_LC_13_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__34913\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \ADC_VDC.genclk.div_state_1__N_1266\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i19148_2_lut_4_lut_LC_13_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111110111111"
        )
    port map (
            in0 => \N__34914\,
            in1 => \N__33780\,
            in2 => \N__34975\,
            in3 => \N__32382\,
            lcout => \ADC_VDC.genclk.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i19194_4_lut_3_lut_LC_13_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__55458\,
            in1 => \N__48737\,
            in2 => \_gnd_net_\,
            in3 => \N__43562\,
            lcout => \comm_spi.n22635\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i24_4_lut_LC_13_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100001010"
        )
    port map (
            in0 => \N__34648\,
            in1 => \N__34154\,
            in2 => \N__34384\,
            in3 => \N__34466\,
            lcout => OPEN,
            ltout => \ADC_VDC.n11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_4_lut_LC_13_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011110000"
        )
    port map (
            in0 => \N__34360\,
            in1 => \N__32557\,
            in2 => \N__32560\,
            in3 => \N__34769\,
            lcout => \ADC_VDC.n18381\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i14977_2_lut_LC_13_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34465\,
            in2 => \_gnd_net_\,
            in3 => \N__34153\,
            lcout => \ADC_VDC.n17359\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.bit_cnt_3769__i0_LC_13_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32547\,
            in2 => \_gnd_net_\,
            in3 => \N__32518\,
            lcout => \ADC_VDC.bit_cnt_0\,
            ltout => OPEN,
            carryin => \bfn_13_6_0_\,
            carryout => \ADC_VDC.n19469\,
            clk => \N__32727\,
            ce => \N__34012\,
            sr => \N__32671\
        );

    \ADC_VDC.bit_cnt_3769__i1_LC_13_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32510\,
            in2 => \_gnd_net_\,
            in3 => \N__32479\,
            lcout => \ADC_VDC.bit_cnt_1\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19469\,
            carryout => \ADC_VDC.n19470\,
            clk => \N__32727\,
            ce => \N__34012\,
            sr => \N__32671\
        );

    \ADC_VDC.bit_cnt_3769__i2_LC_13_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32595\,
            in2 => \_gnd_net_\,
            in3 => \N__32476\,
            lcout => \ADC_VDC.bit_cnt_2\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19470\,
            carryout => \ADC_VDC.n19471\,
            clk => \N__32727\,
            ce => \N__34012\,
            sr => \N__32671\
        );

    \ADC_VDC.bit_cnt_3769__i3_LC_13_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32633\,
            in2 => \_gnd_net_\,
            in3 => \N__32473\,
            lcout => \ADC_VDC.bit_cnt_3\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19471\,
            carryout => \ADC_VDC.n19472\,
            clk => \N__32727\,
            ce => \N__34012\,
            sr => \N__32671\
        );

    \ADC_VDC.bit_cnt_3769__i4_LC_13_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32466\,
            in2 => \_gnd_net_\,
            in3 => \N__32440\,
            lcout => \ADC_VDC.bit_cnt_4\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19472\,
            carryout => \ADC_VDC.n19473\,
            clk => \N__32727\,
            ce => \N__34012\,
            sr => \N__32671\
        );

    \ADC_VDC.bit_cnt_3769__i5_LC_13_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32437\,
            in2 => \_gnd_net_\,
            in3 => \N__32419\,
            lcout => \ADC_VDC.bit_cnt_5\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19473\,
            carryout => \ADC_VDC.n19474\,
            clk => \N__32727\,
            ce => \N__34012\,
            sr => \N__32671\
        );

    \ADC_VDC.bit_cnt_3769__i6_LC_13_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32953\,
            in2 => \_gnd_net_\,
            in3 => \N__32938\,
            lcout => \ADC_VDC.bit_cnt_6\,
            ltout => OPEN,
            carryin => \ADC_VDC.n19474\,
            carryout => \ADC_VDC.n19475\,
            clk => \N__32727\,
            ce => \N__34012\,
            sr => \N__32671\
        );

    \ADC_VDC.bit_cnt_3769__i7_LC_13_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32932\,
            in2 => \_gnd_net_\,
            in3 => \N__32935\,
            lcout => \ADC_VDC.bit_cnt_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32727\,
            ce => \N__34012\,
            sr => \N__32671\
        );

    \comm_spi.imiso_83_12193_12194_set_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__40213\,
            in1 => \N__44272\,
            in2 => \_gnd_net_\,
            in3 => \N__40192\,
            lcout => \comm_spi.n14595\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.imiso_83_12193_12194_setC_net\,
            ce => 'H',
            sr => \N__40261\
        );

    \mux_130_Mux_6_i30_3_lut_LC_13_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__32659\,
            in1 => \N__41215\,
            in2 => \_gnd_net_\,
            in3 => \N__56256\,
            lcout => n30_adj_1595,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_2_lut_adj_33_LC_13_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32625\,
            in2 => \_gnd_net_\,
            in3 => \N__32591\,
            lcout => \ADC_VDC.n6_adj_1404\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_104_2_lut_LC_13_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__55461\,
            in1 => \N__37628\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \comm_spi.data_tx_7__N_778\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_96_2_lut_LC_13_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__37629\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55462\,
            lcout => \comm_spi.data_tx_7__N_762\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i3_12209_12210_set_LC_13_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__37666\,
            in1 => \N__37726\,
            in2 => \_gnd_net_\,
            in3 => \N__37693\,
            lcout => \comm_spi.n14611\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52425\,
            ce => 'H',
            sr => \N__33049\
        );

    \i9327_1_lut_LC_13_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50255\,
            lcout => n11727,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.bit_cnt_3767__i1_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__33010\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33032\,
            lcout => \comm_spi.bit_cnt_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.bit_cnt_3767__i1C_net\,
            ce => 'H',
            sr => \N__55437\
        );

    \comm_spi.bit_cnt_3767__i0_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33009\,
            lcout => \comm_spi.bit_cnt_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.bit_cnt_3767__i1C_net\,
            ce => 'H',
            sr => \N__55437\
        );

    \comm_spi.bit_cnt_3767__i3_LC_13_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__32988\,
            in1 => \N__46377\,
            in2 => \N__33016\,
            in3 => \N__33034\,
            lcout => \comm_spi.bit_cnt_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.bit_cnt_3767__i1C_net\,
            ce => 'H',
            sr => \N__55437\
        );

    \comm_spi.bit_cnt_3767__i2_LC_13_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111011110001000"
        )
    port map (
            in0 => \N__33033\,
            in1 => \N__33011\,
            in2 => \_gnd_net_\,
            in3 => \N__32987\,
            lcout => \comm_spi.bit_cnt_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.bit_cnt_3767__i1C_net\,
            ce => 'H',
            sr => \N__55437\
        );

    \i1_2_lut_3_lut_adj_275_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__54387\,
            in1 => \N__51210\,
            in2 => \_gnd_net_\,
            in3 => \N__53901\,
            lcout => n20653,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15208_2_lut_3_lut_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000100"
        )
    port map (
            in0 => \N__53903\,
            in1 => \N__42804\,
            in2 => \N__51261\,
            in3 => \_gnd_net_\,
            lcout => n14_adj_1528,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i2_3_lut_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__33031\,
            in1 => \N__33015\,
            in2 => \_gnd_net_\,
            in3 => \N__32989\,
            lcout => \comm_spi.n16858\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_0__bdd_4_lut_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__35149\,
            in1 => \N__49520\,
            in2 => \N__32971\,
            in3 => \N__51623\,
            lcout => OPEN,
            ltout => \n21991_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n21991_bdd_4_lut_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__49521\,
            in1 => \N__43383\,
            in2 => \N__32956\,
            in3 => \N__44112\,
            lcout => n21994,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12366_2_lut_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54388\,
            in2 => \_gnd_net_\,
            in3 => \N__49821\,
            lcout => n14763,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15190_2_lut_3_lut_LC_13_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__36394\,
            in1 => \N__51217\,
            in2 => \_gnd_net_\,
            in3 => \N__53904\,
            lcout => n14_adj_1558,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15207_2_lut_3_lut_LC_13_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000100"
        )
    port map (
            in0 => \N__53902\,
            in1 => \N__46646\,
            in2 => \N__51260\,
            in3 => \_gnd_net_\,
            lcout => n14_adj_1527,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_0__bdd_4_lut_19374_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__35191\,
            in1 => \N__49530\,
            in2 => \N__33100\,
            in3 => \N__51624\,
            lcout => OPEN,
            ltout => \n21979_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n21979_bdd_4_lut_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__49531\,
            in1 => \N__43768\,
            in2 => \N__33085\,
            in3 => \N__36395\,
            lcout => n21982,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_137_Mux_3_i4_3_lut_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35461\,
            in1 => \N__33082\,
            in2 => \_gnd_net_\,
            in3 => \N__51625\,
            lcout => OPEN,
            ltout => \n4_adj_1567_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18188_4_lut_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__51626\,
            in1 => \N__33076\,
            in2 => \N__33061\,
            in3 => \N__49534\,
            lcout => OPEN,
            ltout => \n20783_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i3_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__50069\,
            in1 => \_gnd_net_\,
            in2 => \N__33058\,
            in3 => \N__33055\,
            lcout => comm_tx_buf_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55098\,
            ce => \N__47128\,
            sr => \N__47061\
        );

    \i14948_3_lut_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35674\,
            in1 => \N__50182\,
            in2 => \_gnd_net_\,
            in3 => \N__50067\,
            lcout => OPEN,
            ltout => \n17331_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18308_4_lut_LC_13_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__50068\,
            in1 => \N__33190\,
            in2 => \N__33175\,
            in3 => \N__49532\,
            lcout => OPEN,
            ltout => \n20903_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i5_LC_13_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__51627\,
            in1 => \_gnd_net_\,
            in2 => \N__33172\,
            in3 => \N__38221\,
            lcout => comm_tx_buf_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55098\,
            ce => \N__47128\,
            sr => \N__47061\
        );

    \mux_137_Mux_6_i1_3_lut_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__40785\,
            in1 => \N__51428\,
            in2 => \_gnd_net_\,
            in3 => \N__51631\,
            lcout => OPEN,
            ltout => \n1_adj_1561_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i6_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011011000"
        )
    port map (
            in0 => \N__33112\,
            in1 => \N__33133\,
            in2 => \N__33169\,
            in3 => \N__50099\,
            lcout => comm_tx_buf_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55107\,
            ce => \N__47140\,
            sr => \N__47065\
        );

    \i18895_2_lut_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33162\,
            in2 => \_gnd_net_\,
            in3 => \N__51628\,
            lcout => n21051,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_137_Mux_6_i2_3_lut_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__51630\,
            in1 => \_gnd_net_\,
            in2 => \N__33148\,
            in3 => \N__35212\,
            lcout => n2_adj_1562,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_137_Mux_6_i4_3_lut_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35701\,
            in1 => \N__33127\,
            in2 => \_gnd_net_\,
            in3 => \N__51629\,
            lcout => OPEN,
            ltout => \n4_adj_1563_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_1__bdd_4_lut_19472_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010101010"
        )
    port map (
            in0 => \N__49533\,
            in1 => \N__33121\,
            in2 => \N__33115\,
            in3 => \N__50098\,
            lcout => n22093,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_101_2_lut_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__55459\,
            in1 => \N__40274\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \comm_spi.data_tx_7__N_769\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_93_2_lut_LC_13_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__40275\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55460\,
            lcout => \comm_spi.data_tx_7__N_759\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_2_i26_3_lut_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__33336\,
            in1 => \N__56832\,
            in2 => \_gnd_net_\,
            in3 => \N__46882\,
            lcout => OPEN,
            ltout => \n26_adj_1506_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18221_4_lut_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__56833\,
            in1 => \N__57482\,
            in2 => \N__33325\,
            in3 => \N__33322\,
            lcout => OPEN,
            ltout => \n20816_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_2__bdd_4_lut_19561_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__47788\,
            in1 => \N__33238\,
            in2 => \N__33304\,
            in3 => \N__56289\,
            lcout => OPEN,
            ltout => \n22087_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22087_bdd_4_lut_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__56290\,
            in1 => \N__33301\,
            in2 => \N__33286\,
            in3 => \N__33244\,
            lcout => OPEN,
            ltout => \n22090_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i2_LC_13_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35452\,
            in2 => \N__33283\,
            in3 => \N__53908\,
            lcout => comm_buf_1_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55118\,
            ce => \N__38544\,
            sr => \N__36807\
        );

    \i18251_3_lut_LC_13_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__33280\,
            in1 => \N__33271\,
            in2 => \_gnd_net_\,
            in3 => \N__57481\,
            lcout => n20846,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18220_3_lut_LC_13_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__57480\,
            in1 => \N__41596\,
            in2 => \_gnd_net_\,
            in3 => \N__36304\,
            lcout => n20815,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19477_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__33232\,
            in1 => \N__57532\,
            in2 => \N__33217\,
            in3 => \N__47782\,
            lcout => OPEN,
            ltout => \n22081_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22081_bdd_4_lut_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__47783\,
            in1 => \N__33469\,
            in2 => \N__33442\,
            in3 => \N__36124\,
            lcout => n22084,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_4_i26_3_lut_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__33438\,
            in1 => \N__56840\,
            in2 => \_gnd_net_\,
            in3 => \N__46813\,
            lcout => OPEN,
            ltout => \n26_adj_1484_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19531_LC_13_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110100000"
        )
    port map (
            in0 => \N__47784\,
            in1 => \N__33421\,
            in2 => \N__33409\,
            in3 => \N__57483\,
            lcout => OPEN,
            ltout => \n22159_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22159_bdd_4_lut_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011000010"
        )
    port map (
            in0 => \N__36949\,
            in1 => \N__47785\,
            in2 => \N__33406\,
            in3 => \N__38395\,
            lcout => OPEN,
            ltout => \n22162_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1541671_i1_3_lut_LC_13_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33403\,
            in2 => \N__33397\,
            in3 => \N__56287\,
            lcout => OPEN,
            ltout => \n30_adj_1493_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i4_LC_13_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35661\,
            in2 => \N__33394\,
            in3 => \N__54000\,
            lcout => comm_buf_1_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55127\,
            ce => \N__38550\,
            sr => \N__36790\
        );

    \mux_129_Mux_3_i26_3_lut_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__56841\,
            in1 => \N__33391\,
            in2 => \_gnd_net_\,
            in3 => \N__46851\,
            lcout => OPEN,
            ltout => \n26_adj_1502_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111000000"
        )
    port map (
            in0 => \N__33376\,
            in1 => \N__47780\,
            in2 => \N__33361\,
            in3 => \N__57550\,
            lcout => OPEN,
            ltout => \n22195_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22195_bdd_4_lut_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__47781\,
            in1 => \N__38833\,
            in2 => \N__33358\,
            in3 => \N__33355\,
            lcout => OPEN,
            ltout => \n22198_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1540465_i1_3_lut_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33502\,
            in2 => \N__33589\,
            in3 => \N__56288\,
            lcout => OPEN,
            ltout => \n30_adj_1503_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i3_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35569\,
            in2 => \N__33586\,
            in3 => \N__53909\,
            lcout => comm_buf_1_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55139\,
            ce => \N__38545\,
            sr => \N__36796\
        );

    \comm_cmd_1__bdd_4_lut_19403_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110001000"
        )
    port map (
            in0 => \N__33583\,
            in1 => \N__47778\,
            in2 => \N__33571\,
            in3 => \N__57549\,
            lcout => OPEN,
            ltout => \n22009_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22009_bdd_4_lut_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__47779\,
            in1 => \N__33541\,
            in2 => \N__33514\,
            in3 => \N__33511\,
            lcout => n22012,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipcnt_i0_i0_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46956\,
            in2 => \N__33496\,
            in3 => \_gnd_net_\,
            lcout => acadc_skipcnt_0,
            ltout => OPEN,
            carryin => \bfn_13_16_0_\,
            carryout => n19311,
            clk => \INVacadc_skipcnt_i0_i0C_net\,
            ce => \N__33936\,
            sr => \N__33481\
        );

    \add_73_2_THRU_CRY_0_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52799\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => n19311,
            carryout => \n19311_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_73_2_THRU_CRY_1_LC_13_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52803\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \n19311_THRU_CRY_0_THRU_CO\,
            carryout => \n19311_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_73_2_THRU_CRY_2_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52800\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \n19311_THRU_CRY_1_THRU_CO\,
            carryout => \n19311_THRU_CRY_2_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_73_2_THRU_CRY_3_LC_13_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52804\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \n19311_THRU_CRY_2_THRU_CO\,
            carryout => \n19311_THRU_CRY_3_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_73_2_THRU_CRY_4_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52801\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \n19311_THRU_CRY_3_THRU_CO\,
            carryout => \n19311_THRU_CRY_4_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_73_2_THRU_CRY_5_LC_13_16_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52805\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \n19311_THRU_CRY_4_THRU_CO\,
            carryout => \n19311_THRU_CRY_5_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_73_2_THRU_CRY_6_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52802\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \n19311_THRU_CRY_5_THRU_CO\,
            carryout => \n19311_THRU_CRY_6_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipcnt_i0_i1_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33675\,
            in2 => \_gnd_net_\,
            in3 => \N__33661\,
            lcout => acadc_skipcnt_1,
            ltout => OPEN,
            carryin => \bfn_13_17_0_\,
            carryout => n19312,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__33923\,
            sr => \N__33894\
        );

    \acadc_skipcnt_i0_i2_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36333\,
            in2 => \_gnd_net_\,
            in3 => \N__33658\,
            lcout => acadc_skipcnt_2,
            ltout => OPEN,
            carryin => n19312,
            carryout => n19313,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__33923\,
            sr => \N__33894\
        );

    \acadc_skipcnt_i0_i3_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33654\,
            in2 => \_gnd_net_\,
            in3 => \N__33637\,
            lcout => acadc_skipcnt_3,
            ltout => OPEN,
            carryin => n19313,
            carryout => n19314,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__33923\,
            sr => \N__33894\
        );

    \acadc_skipcnt_i0_i4_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33630\,
            in2 => \_gnd_net_\,
            in3 => \N__33613\,
            lcout => acadc_skipcnt_4,
            ltout => OPEN,
            carryin => n19314,
            carryout => n19315,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__33923\,
            sr => \N__33894\
        );

    \acadc_skipcnt_i0_i5_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33606\,
            in2 => \_gnd_net_\,
            in3 => \N__33592\,
            lcout => acadc_skipcnt_5,
            ltout => OPEN,
            carryin => n19315,
            carryout => n19316,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__33923\,
            sr => \N__33894\
        );

    \acadc_skipcnt_i0_i6_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33753\,
            in2 => \_gnd_net_\,
            in3 => \N__33739\,
            lcout => acadc_skipcnt_6,
            ltout => OPEN,
            carryin => n19316,
            carryout => n19317,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__33923\,
            sr => \N__33894\
        );

    \acadc_skipcnt_i0_i7_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36318\,
            in2 => \_gnd_net_\,
            in3 => \N__33736\,
            lcout => acadc_skipcnt_7,
            ltout => OPEN,
            carryin => n19317,
            carryout => n19318,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__33923\,
            sr => \N__33894\
        );

    \acadc_skipcnt_i0_i8_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33729\,
            in2 => \_gnd_net_\,
            in3 => \N__33715\,
            lcout => acadc_skipcnt_8,
            ltout => OPEN,
            carryin => n19318,
            carryout => n19319,
            clk => \INVacadc_skipcnt_i0_i1C_net\,
            ce => \N__33923\,
            sr => \N__33894\
        );

    \acadc_skipcnt_i0_i9_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36627\,
            in2 => \_gnd_net_\,
            in3 => \N__33712\,
            lcout => acadc_skipcnt_9,
            ltout => OPEN,
            carryin => \bfn_13_18_0_\,
            carryout => n19320,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__33937\,
            sr => \N__33898\
        );

    \acadc_skipcnt_i0_i10_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38790\,
            in2 => \_gnd_net_\,
            in3 => \N__33709\,
            lcout => acadc_skipcnt_10,
            ltout => OPEN,
            carryin => n19320,
            carryout => n19321,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__33937\,
            sr => \N__33898\
        );

    \acadc_skipcnt_i0_i11_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36411\,
            in2 => \_gnd_net_\,
            in3 => \N__33706\,
            lcout => acadc_skipcnt_11,
            ltout => OPEN,
            carryin => n19321,
            carryout => n19322,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__33937\,
            sr => \N__33898\
        );

    \acadc_skipcnt_i0_i12_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38808\,
            in2 => \_gnd_net_\,
            in3 => \N__33703\,
            lcout => acadc_skipcnt_12,
            ltout => OPEN,
            carryin => n19322,
            carryout => n19323,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__33937\,
            sr => \N__33898\
        );

    \acadc_skipcnt_i0_i13_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33696\,
            in2 => \_gnd_net_\,
            in3 => \N__33682\,
            lcout => acadc_skipcnt_13,
            ltout => OPEN,
            carryin => n19323,
            carryout => n19324,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__33937\,
            sr => \N__33898\
        );

    \acadc_skipcnt_i0_i14_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36426\,
            in2 => \_gnd_net_\,
            in3 => \N__33679\,
            lcout => acadc_skipcnt_14,
            ltout => OPEN,
            carryin => n19324,
            carryout => n19325,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__33937\,
            sr => \N__33898\
        );

    \acadc_skipcnt_i0_i15_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36612\,
            in2 => \_gnd_net_\,
            in3 => \N__33940\,
            lcout => acadc_skipcnt_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVacadc_skipcnt_i0_i9C_net\,
            ce => \N__33937\,
            sr => \N__33898\
        );

    \SIG_DDS.tmp_buf_i12_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__55878\,
            in1 => \N__55660\,
            in2 => \N__33877\,
            in3 => \N__33868\,
            lcout => \SIG_DDS.tmp_buf_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55196\,
            ce => \N__40315\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i2_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__55879\,
            in1 => \N__55661\,
            in2 => \N__33829\,
            in3 => \N__42754\,
            lcout => \SIG_DDS.tmp_buf_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55196\,
            ce => \N__40315\,
            sr => \_gnd_net_\
        );

    \comm_spi.data_rx_i0_12197_12198_reset_LC_14_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__37425\,
            in1 => \N__34996\,
            in2 => \_gnd_net_\,
            in3 => \N__33819\,
            lcout => \comm_spi.n14600\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52441\,
            ce => 'H',
            sr => \N__33796\
        );

    \ADC_VDC.genclk.i18725_4_lut_LC_14_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__37017\,
            in1 => \N__37110\,
            in2 => \N__37063\,
            in3 => \N__37125\,
            lcout => OPEN,
            ltout => \ADC_VDC.genclk.n21172_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i18906_4_lut_LC_14_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__33769\,
            in1 => \N__33760\,
            in2 => \N__33784\,
            in3 => \N__35002\,
            lcout => \ADC_VDC.genclk.n21166\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i12_4_lut_adj_27_LC_14_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37170\,
            in1 => \N__37251\,
            in2 => \N__37498\,
            in3 => \N__37218\,
            lcout => \ADC_VDC.genclk.n28_adj_1400\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i10_4_lut_adj_28_LC_14_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37077\,
            in1 => \N__37185\,
            in2 => \N__37039\,
            in3 => \N__37269\,
            lcout => \ADC_VDC.genclk.n26_adj_1401\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.i11_4_lut_adj_29_LC_14_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__37203\,
            in1 => \N__37092\,
            in2 => \N__37288\,
            in3 => \N__37236\,
            lcout => \ADC_VDC.genclk.n27_adj_1402\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.imosi_44_12183_12184_reset_LC_14_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37342\,
            lcout => \comm_spi.n14586\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55074\,
            ce => 'H',
            sr => \N__37300\
        );

    \ADC_VDC.genclk.div_state_i1_LC_14_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34974\,
            in2 => \_gnd_net_\,
            in3 => \N__34918\,
            lcout => \ADC_VDC.genclk.div_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADC_VDC.genclk.div_state_i1C_net\,
            ce => \N__34885\,
            sr => \_gnd_net_\
        );

    \ADC_VDC.i1_2_lut_LC_14_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__34872\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34747\,
            lcout => \ADC_VDC.n62\,
            ltout => \ADC_VDC.n62_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VDC.i16006_4_lut_LC_14_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100010111010"
        )
    port map (
            in0 => \N__34566\,
            in1 => \N__34375\,
            in2 => \N__34162\,
            in3 => \N__34155\,
            lcout => \ADC_VDC.n11736\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_137_Mux_7_i2_3_lut_LC_14_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__34003\,
            in1 => \N__35230\,
            in2 => \_gnd_net_\,
            in3 => \N__51622\,
            lcout => OPEN,
            ltout => \n2_adj_1559_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i7_LC_14_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001000100"
        )
    port map (
            in0 => \N__50101\,
            in1 => \N__33988\,
            in2 => \N__33979\,
            in3 => \N__35044\,
            lcout => comm_tx_buf_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55077\,
            ce => \N__47124\,
            sr => \N__47056\
        );

    \mux_137_Mux_7_i4_3_lut_LC_14_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35110\,
            in1 => \N__33976\,
            in2 => \_gnd_net_\,
            in3 => \N__51620\,
            lcout => n4_adj_1560,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19043_2_lut_LC_14_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__51621\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33964\,
            lcout => OPEN,
            ltout => \n21276_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_1__bdd_4_lut_LC_14_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__35053\,
            in1 => \N__49529\,
            in2 => \N__35047\,
            in3 => \N__50100\,
            lcout => n22105,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i19164_4_lut_3_lut_LC_14_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44271\,
            in1 => \N__37391\,
            in2 => \_gnd_net_\,
            in3 => \N__55409\,
            lcout => \comm_spi.n14588\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_100_2_lut_LC_14_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__55408\,
            in1 => \_gnd_net_\,
            in2 => \N__37396\,
            in3 => \_gnd_net_\,
            lcout => \comm_spi.data_tx_7__N_766\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_0__bdd_4_lut_19379_LC_14_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001001010"
        )
    port map (
            in0 => \N__51638\,
            in1 => \N__35173\,
            in2 => \N__49543\,
            in3 => \N__35038\,
            lcout => OPEN,
            ltout => \n21985_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n21985_bdd_4_lut_LC_14_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__49536\,
            in1 => \N__38712\,
            in2 => \N__35026\,
            in3 => \N__42815\,
            lcout => OPEN,
            ltout => \n21988_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i2_LC_14_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__50077\,
            in1 => \_gnd_net_\,
            in2 => \N__35023\,
            in3 => \N__35059\,
            lcout => comm_tx_buf_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55085\,
            ce => \N__47136\,
            sr => \N__47057\
        );

    \i14920_3_lut_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35131\,
            in1 => \N__41354\,
            in2 => \_gnd_net_\,
            in3 => \N__50075\,
            lcout => OPEN,
            ltout => \n17304_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18311_4_lut_LC_14_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__50076\,
            in1 => \N__35020\,
            in2 => \N__35008\,
            in3 => \N__49537\,
            lcout => OPEN,
            ltout => \n20906_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i0_LC_14_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38113\,
            in2 => \N__35005\,
            in3 => \N__51641\,
            lcout => comm_tx_buf_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55085\,
            ce => \N__47136\,
            sr => \N__47057\
        );

    \mux_137_Mux_2_i4_3_lut_LC_14_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__51639\,
            in1 => \N__35356\,
            in2 => \_gnd_net_\,
            in3 => \N__35098\,
            lcout => OPEN,
            ltout => \n4_adj_1568_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18191_4_lut_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__49535\,
            in1 => \N__35086\,
            in2 => \N__35062\,
            in3 => \N__51640\,
            lcout => n20786,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_rx_i7_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__46376\,
            in1 => \N__35757\,
            in2 => \_gnd_net_\,
            in3 => \N__46332\,
            lcout => comm_rx_buf_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52443\,
            ce => 'H',
            sr => \N__55431\
        );

    \comm_spi.data_rx_i6_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__46331\,
            in1 => \N__37953\,
            in2 => \_gnd_net_\,
            in3 => \N__46375\,
            lcout => comm_rx_buf_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52443\,
            ce => 'H',
            sr => \N__55431\
        );

    \comm_spi.data_rx_i5_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__46374\,
            in1 => \N__35617\,
            in2 => \_gnd_net_\,
            in3 => \N__46330\,
            lcout => comm_rx_buf_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52443\,
            ce => 'H',
            sr => \N__55431\
        );

    \comm_spi.data_rx_i4_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__46329\,
            in1 => \N__35509\,
            in2 => \_gnd_net_\,
            in3 => \N__46373\,
            lcout => comm_rx_buf_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52443\,
            ce => 'H',
            sr => \N__55431\
        );

    \comm_spi.data_rx_i3_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__46372\,
            in1 => \N__35401\,
            in2 => \_gnd_net_\,
            in3 => \N__46328\,
            lcout => comm_rx_buf_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52443\,
            ce => 'H',
            sr => \N__55431\
        );

    \comm_spi.data_rx_i2_LC_14_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__46327\,
            in1 => \N__35933\,
            in2 => \_gnd_net_\,
            in3 => \N__46371\,
            lcout => comm_rx_buf_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52443\,
            ce => 'H',
            sr => \N__55431\
        );

    \comm_spi.data_rx_i1_LC_14_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000000000"
        )
    port map (
            in0 => \N__46370\,
            in1 => \N__46326\,
            in2 => \_gnd_net_\,
            in3 => \N__36241\,
            lcout => comm_rx_buf_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52443\,
            ce => 'H',
            sr => \N__55431\
        );

    \comm_buf_2__i0_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__35239\,
            in1 => \N__53938\,
            in2 => \_gnd_net_\,
            in3 => \N__36233\,
            lcout => comm_buf_2_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55099\,
            ce => \N__37921\,
            sr => \N__38350\
        );

    \comm_buf_2__i7_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__53937\,
            in1 => \_gnd_net_\,
            in2 => \N__36858\,
            in3 => \N__47428\,
            lcout => comm_buf_2_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55099\,
            ce => \N__37921\,
            sr => \N__38350\
        );

    \comm_buf_2__i6_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35758\,
            in1 => \N__35221\,
            in2 => \_gnd_net_\,
            in3 => \N__53941\,
            lcout => comm_buf_2_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55099\,
            ce => \N__37921\,
            sr => \N__38350\
        );

    \comm_buf_2__i4_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__53936\,
            in1 => \N__35618\,
            in2 => \_gnd_net_\,
            in3 => \N__56053\,
            lcout => comm_buf_2_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55099\,
            ce => \N__37921\,
            sr => \N__38350\
        );

    \comm_buf_2__i3_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35510\,
            in1 => \N__35203\,
            in2 => \_gnd_net_\,
            in3 => \N__53940\,
            lcout => comm_buf_2_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55099\,
            ce => \N__37921\,
            sr => \N__38350\
        );

    \comm_buf_2__i2_LC_14_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__53935\,
            in1 => \_gnd_net_\,
            in2 => \N__35420\,
            in3 => \N__35185\,
            lcout => comm_buf_2_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55099\,
            ce => \N__37921\,
            sr => \N__38350\
        );

    \comm_buf_2__i1_LC_14_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35934\,
            in1 => \N__35164\,
            in2 => \_gnd_net_\,
            in3 => \N__53939\,
            lcout => comm_buf_2_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55099\,
            ce => \N__37921\,
            sr => \N__38350\
        );

    \comm_buf_5__i0_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__35143\,
            in1 => \N__53946\,
            in2 => \_gnd_net_\,
            in3 => \N__36237\,
            lcout => comm_buf_5_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55108\,
            ce => \N__38104\,
            sr => \N__38092\
        );

    \comm_buf_5__i7_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__53945\,
            in1 => \_gnd_net_\,
            in2 => \N__36880\,
            in3 => \N__35119\,
            lcout => comm_buf_5_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55108\,
            ce => \N__38104\,
            sr => \N__38092\
        );

    \comm_buf_5__i6_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35779\,
            in1 => \N__35716\,
            in2 => \_gnd_net_\,
            in3 => \N__53949\,
            lcout => comm_buf_5_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55108\,
            ce => \N__38104\,
            sr => \N__38092\
        );

    \comm_buf_5__i5_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__53944\,
            in1 => \_gnd_net_\,
            in2 => \N__37994\,
            in3 => \N__35689\,
            lcout => comm_buf_5_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55108\,
            ce => \N__38104\,
            sr => \N__38092\
        );

    \comm_buf_5__i4_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35636\,
            in1 => \N__35584\,
            in2 => \_gnd_net_\,
            in3 => \N__53948\,
            lcout => comm_buf_5_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55108\,
            ce => \N__38104\,
            sr => \N__38092\
        );

    \comm_buf_5__i3_LC_14_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__53943\,
            in1 => \N__35530\,
            in2 => \_gnd_net_\,
            in3 => \N__35482\,
            lcout => comm_buf_5_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55108\,
            ce => \N__38104\,
            sr => \N__38092\
        );

    \comm_buf_5__i2_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35421\,
            in1 => \N__35368\,
            in2 => \_gnd_net_\,
            in3 => \N__53947\,
            lcout => comm_buf_5_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55108\,
            ce => \N__38104\,
            sr => \N__38092\
        );

    \comm_buf_5__i1_LC_14_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__53942\,
            in1 => \N__35951\,
            in2 => \_gnd_net_\,
            in3 => \N__35347\,
            lcout => comm_buf_5_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55108\,
            ce => \N__38104\,
            sr => \N__38092\
        );

    \i18242_3_lut_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__57552\,
            in1 => \N__35335\,
            in2 => \_gnd_net_\,
            in3 => \N__35245\,
            lcout => n20837,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_1_i19_3_lut_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__56950\,
            in1 => \N__35308\,
            in2 => \_gnd_net_\,
            in3 => \N__35283\,
            lcout => n19_adj_1508,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_2__bdd_4_lut_19457_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101001100010"
        )
    port map (
            in0 => \N__47847\,
            in1 => \N__56264\,
            in2 => \N__36079\,
            in3 => \N__36001\,
            lcout => OPEN,
            ltout => \n22069_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22069_bdd_4_lut_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__56265\,
            in1 => \N__36067\,
            in2 => \N__36049\,
            in3 => \N__36046\,
            lcout => n22072,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_1_i26_3_lut_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__36040\,
            in1 => \N__56949\,
            in2 => \_gnd_net_\,
            in3 => \N__46908\,
            lcout => OPEN,
            ltout => \n26_adj_1509_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18230_4_lut_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__56951\,
            in1 => \N__57551\,
            in2 => \N__36025\,
            in3 => \N__36022\,
            lcout => n20825,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i1_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__35971\,
            in1 => \N__54031\,
            in2 => \_gnd_net_\,
            in3 => \N__35905\,
            lcout => comm_buf_1_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55119\,
            ce => \N__38523\,
            sr => \N__36780\
        );

    \mux_129_Mux_0_i26_3_lut_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__35899\,
            in1 => \N__56831\,
            in2 => \_gnd_net_\,
            in3 => \N__46935\,
            lcout => OPEN,
            ltout => \n26_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19452_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011001100"
        )
    port map (
            in0 => \N__35881\,
            in1 => \N__57479\,
            in2 => \N__35863\,
            in3 => \N__47726\,
            lcout => OPEN,
            ltout => \n22021_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22021_bdd_4_lut_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__47727\,
            in1 => \N__35860\,
            in2 => \N__35833\,
            in3 => \N__41752\,
            lcout => n22024,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1541068_i1_3_lut_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__35830\,
            in1 => \N__35824\,
            in2 => \_gnd_net_\,
            in3 => \N__56269\,
            lcout => OPEN,
            ltout => \n30_adj_1478_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i0_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54032\,
            in2 => \N__36262\,
            in3 => \N__36253\,
            lcout => comm_buf_1_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55128\,
            ce => \N__38533\,
            sr => \N__36795\
        );

    \ADC_VAC.ADC_DATA_i5_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__48526\,
            in1 => \N__48350\,
            in2 => \N__38304\,
            in3 => \N__36165\,
            lcout => buf_adcdata_vac_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55140\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i13_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100000110000"
        )
    port map (
            in0 => \N__48349\,
            in1 => \N__37884\,
            in2 => \N__36166\,
            in3 => \N__47967\,
            lcout => cmd_rdadctmp_13_adj_1430,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55140\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i14_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__37885\,
            in1 => \N__36164\,
            in2 => \N__38759\,
            in3 => \N__48351\,
            lcout => cmd_rdadctmp_14_adj_1429,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55140\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12345_2_lut_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54600\,
            in2 => \_gnd_net_\,
            in3 => \N__38497\,
            lcout => n14742,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i6_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__36108\,
            in1 => \N__45876\,
            in2 => \N__51430\,
            in3 => \N__45987\,
            lcout => buf_dds1_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55140\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_4_i16_3_lut_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__36151\,
            in1 => \N__42711\,
            in2 => \_gnd_net_\,
            in3 => \N__56983\,
            lcout => n16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_6_i16_3_lut_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__56984\,
            in1 => \N__36104\,
            in2 => \_gnd_net_\,
            in3 => \N__42654\,
            lcout => n16_adj_1488,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18229_3_lut_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__57525\,
            in1 => \N__36564\,
            in2 => \_gnd_net_\,
            in3 => \N__38374\,
            lcout => n20824,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_354_Mux_2_i15_4_lut_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__36636\,
            in1 => \N__54670\,
            in2 => \N__51984\,
            in3 => \N__41841\,
            lcout => \data_index_9_N_212_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7_4_lut_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__36430\,
            in1 => \N__36412\,
            in2 => \N__45477\,
            in3 => \N__36653\,
            lcout => n23_adj_1586,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6412_3_lut_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__41827\,
            in1 => \N__36378\,
            in2 => \_gnd_net_\,
            in3 => \N__43273\,
            lcout => n8_adj_1543,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i2_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__51893\,
            in1 => \N__39313\,
            in2 => \N__42808\,
            in3 => \N__36302\,
            lcout => \acadc_skipCount_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55153\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i2_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011101100001000"
        )
    port map (
            in0 => \N__36637\,
            in1 => \N__54671\,
            in2 => \N__51985\,
            in3 => \N__41842\,
            lcout => data_index_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55153\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6_4_lut_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__36334\,
            in1 => \N__36319\,
            in2 => \N__36303\,
            in3 => \N__36977\,
            lcout => OPEN,
            ltout => \n22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14_4_lut_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__36280\,
            in1 => \N__38776\,
            in2 => \N__36274\,
            in3 => \N__36574\,
            lcout => n30_adj_1571,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i7_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__51894\,
            in1 => \N__39314\,
            in2 => \N__42619\,
            in3 => \N__36978\,
            lcout => \acadc_skipCount_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55153\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i4_LC_14_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__44744\,
            in1 => \N__43847\,
            in2 => \_gnd_net_\,
            in3 => \N__42135\,
            lcout => \VDC_RNG0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55168\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i15_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__45766\,
            in1 => \N__39273\,
            in2 => \_gnd_net_\,
            in3 => \N__36588\,
            lcout => \acadc_skipCount_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55168\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_129_Mux_7_i26_3_lut_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47376\,
            in1 => \N__36682\,
            in2 => \_gnd_net_\,
            in3 => \N__56954\,
            lcout => n26_adj_1623,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i14_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__41528\,
            in1 => \N__39272\,
            in2 => \_gnd_net_\,
            in3 => \N__36657\,
            lcout => \acadc_skipCount_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55168\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6422_3_lut_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__42788\,
            in1 => \N__41861\,
            in2 => \_gnd_net_\,
            in3 => \N__43277\,
            lcout => n8_adj_1545,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i6_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__55949\,
            in1 => \_gnd_net_\,
            in2 => \N__41535\,
            in3 => \N__43848\,
            lcout => buf_control_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55168\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_4_lut_adj_175_LC_14_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__57493\,
            in1 => \N__56955\,
            in2 => \N__45382\,
            in3 => \N__47836\,
            lcout => n20626,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i8_4_lut_LC_14_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__36628\,
            in1 => \N__36613\,
            in2 => \N__36921\,
            in3 => \N__36587\,
            lcout => n24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i1_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__43374\,
            in1 => \N__39285\,
            in2 => \N__36568\,
            in3 => \N__52087\,
            lcout => \acadc_skipCount_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55183\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_301_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011000100"
        )
    port map (
            in0 => \N__36538\,
            in1 => \N__54675\,
            in2 => \N__52159\,
            in3 => \N__41626\,
            lcout => n12391,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19350_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011010100010"
        )
    port map (
            in0 => \N__57539\,
            in1 => \N__47844\,
            in2 => \N__37003\,
            in3 => \N__36991\,
            lcout => OPEN,
            ltout => \n21949_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n21949_bdd_4_lut_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__47845\,
            in1 => \N__41569\,
            in2 => \N__36985\,
            in3 => \N__36982\,
            lcout => OPEN,
            ltout => \n21952_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1535641_i1_3_lut_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36964\,
            in2 => \N__36952\,
            in3 => \N__56317\,
            lcout => n30_adj_1624,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i4_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__39286\,
            in1 => \N__46647\,
            in2 => \N__52160\,
            in3 => \N__36947\,
            lcout => \acadc_skipCount_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55183\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i9_LC_14_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__39287\,
            in1 => \N__44127\,
            in2 => \N__52161\,
            in3 => \N__36920\,
            lcout => \acadc_skipCount_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55183\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_1__i7_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__36894\,
            in1 => \N__54090\,
            in2 => \_gnd_net_\,
            in3 => \N__36814\,
            lcout => comm_buf_1_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55197\,
            ce => \N__38540\,
            sr => \N__36803\
        );

    \SIG_DDS.i19068_4_lut_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000100110"
        )
    port map (
            in0 => \N__55866\,
            in1 => \N__55737\,
            in2 => \N__53025\,
            in3 => \N__55628\,
            lcout => \SIG_DDS.n12700\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i3_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__55629\,
            in1 => \N__55867\,
            in2 => \N__36724\,
            in3 => \N__36697\,
            lcout => \SIG_DDS.tmp_buf_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55210\,
            ce => \N__40314\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i4_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__55868\,
            in1 => \N__55630\,
            in2 => \N__36691\,
            in3 => \N__42712\,
            lcout => \SIG_DDS.tmp_buf_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55210\,
            ce => \N__40314\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i5_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__55631\,
            in1 => \N__55869\,
            in2 => \N__37156\,
            in3 => \N__43065\,
            lcout => \SIG_DDS.tmp_buf_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55210\,
            ce => \N__40314\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i6_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__55870\,
            in1 => \N__55632\,
            in2 => \N__37147\,
            in3 => \N__42658\,
            lcout => \SIG_DDS.tmp_buf_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55210\,
            ce => \N__40314\,
            sr => \_gnd_net_\
        );

    \ADC_VDC.genclk.t0on_i0_LC_15_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37126\,
            in2 => \_gnd_net_\,
            in3 => \N__37114\,
            lcout => \ADC_VDC.genclk.t0on_0\,
            ltout => OPEN,
            carryin => \bfn_15_3_0_\,
            carryout => \ADC_VDC.genclk.n19425\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__37483\,
            sr => \N__37452\
        );

    \ADC_VDC.genclk.t0on_i1_LC_15_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37111\,
            in2 => \N__52828\,
            in3 => \N__37099\,
            lcout => \ADC_VDC.genclk.t0on_1\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19425\,
            carryout => \ADC_VDC.genclk.n19426\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__37483\,
            sr => \N__37452\
        );

    \ADC_VDC.genclk.t0on_i2_LC_15_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52776\,
            in2 => \N__37096\,
            in3 => \N__37081\,
            lcout => \ADC_VDC.genclk.t0on_2\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19426\,
            carryout => \ADC_VDC.genclk.n19427\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__37483\,
            sr => \N__37452\
        );

    \ADC_VDC.genclk.t0on_i3_LC_15_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37078\,
            in2 => \N__52829\,
            in3 => \N__37066\,
            lcout => \ADC_VDC.genclk.t0on_3\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19427\,
            carryout => \ADC_VDC.genclk.n19428\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__37483\,
            sr => \N__37452\
        );

    \ADC_VDC.genclk.t0on_i4_LC_15_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52780\,
            in2 => \N__37062\,
            in3 => \N__37042\,
            lcout => \ADC_VDC.genclk.t0on_4\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19428\,
            carryout => \ADC_VDC.genclk.n19429\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__37483\,
            sr => \N__37452\
        );

    \ADC_VDC.genclk.t0on_i5_LC_15_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37038\,
            in2 => \N__52830\,
            in3 => \N__37024\,
            lcout => \ADC_VDC.genclk.t0on_5\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19429\,
            carryout => \ADC_VDC.genclk.n19430\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__37483\,
            sr => \N__37452\
        );

    \ADC_VDC.genclk.t0on_i6_LC_15_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52784\,
            in2 => \N__37021\,
            in3 => \N__37006\,
            lcout => \ADC_VDC.genclk.t0on_6\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19430\,
            carryout => \ADC_VDC.genclk.n19431\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__37483\,
            sr => \N__37452\
        );

    \ADC_VDC.genclk.t0on_i7_LC_15_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37287\,
            in2 => \N__52831\,
            in3 => \N__37273\,
            lcout => \ADC_VDC.genclk.t0on_7\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19431\,
            carryout => \ADC_VDC.genclk.n19432\,
            clk => \INVADC_VDC.genclk.t0on_i0C_net\,
            ce => \N__37483\,
            sr => \N__37452\
        );

    \ADC_VDC.genclk.t0on_i8_LC_15_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37270\,
            in2 => \N__52794\,
            in3 => \N__37258\,
            lcout => \ADC_VDC.genclk.t0on_8\,
            ltout => OPEN,
            carryin => \bfn_15_4_0_\,
            carryout => \ADC_VDC.genclk.n19433\,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__37482\,
            sr => \N__37456\
        );

    \ADC_VDC.genclk.t0on_i9_LC_15_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52719\,
            in2 => \N__37255\,
            in3 => \N__37240\,
            lcout => \ADC_VDC.genclk.t0on_9\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19433\,
            carryout => \ADC_VDC.genclk.n19434\,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__37482\,
            sr => \N__37456\
        );

    \ADC_VDC.genclk.t0on_i10_LC_15_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37237\,
            in2 => \N__52791\,
            in3 => \N__37225\,
            lcout => \ADC_VDC.genclk.t0on_10\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19434\,
            carryout => \ADC_VDC.genclk.n19435\,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__37482\,
            sr => \N__37456\
        );

    \ADC_VDC.genclk.t0on_i11_LC_15_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52707\,
            in2 => \N__37222\,
            in3 => \N__37207\,
            lcout => \ADC_VDC.genclk.t0on_11\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19435\,
            carryout => \ADC_VDC.genclk.n19436\,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__37482\,
            sr => \N__37456\
        );

    \ADC_VDC.genclk.t0on_i12_LC_15_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37204\,
            in2 => \N__52792\,
            in3 => \N__37192\,
            lcout => \ADC_VDC.genclk.t0on_12\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19436\,
            carryout => \ADC_VDC.genclk.n19437\,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__37482\,
            sr => \N__37456\
        );

    \ADC_VDC.genclk.t0on_i13_LC_15_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52711\,
            in2 => \N__37189\,
            in3 => \N__37174\,
            lcout => \ADC_VDC.genclk.t0on_13\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19437\,
            carryout => \ADC_VDC.genclk.n19438\,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__37482\,
            sr => \N__37456\
        );

    \ADC_VDC.genclk.t0on_i14_LC_15_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37171\,
            in2 => \N__52793\,
            in3 => \N__37159\,
            lcout => \ADC_VDC.genclk.t0on_14\,
            ltout => OPEN,
            carryin => \ADC_VDC.genclk.n19438\,
            carryout => \ADC_VDC.genclk.n19439\,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__37482\,
            sr => \N__37456\
        );

    \ADC_VDC.genclk.t0on_i15_LC_15_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__37497\,
            in1 => \N__52715\,
            in2 => \_gnd_net_\,
            in3 => \N__37501\,
            lcout => \ADC_VDC.genclk.t0on_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVADC_VDC.genclk.t0on_i8C_net\,
            ce => \N__37482\,
            sr => \N__37456\
        );

    \comm_spi.imosi_44_12183_12184_set_LC_15_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__37355\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \comm_spi.n14585\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55075\,
            ce => 'H',
            sr => \N__37363\
        );

    \comm_spi.MISO_48_12187_12188_set_LC_15_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44323\,
            in1 => \N__44310\,
            in2 => \_gnd_net_\,
            in3 => \N__44270\,
            lcout => \comm_spi.n14589\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.MISO_48_12187_12188_setC_net\,
            ce => 'H',
            sr => \N__40256\
        );

    \comm_spi.RESET_I_0_105_2_lut_LC_15_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__55424\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37376\,
            lcout => \comm_spi.data_tx_7__N_781\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_92_2_lut_LC_15_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37395\,
            in2 => \_gnd_net_\,
            in3 => \N__55421\,
            lcout => \comm_spi.data_tx_7__N_758\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_97_2_lut_LC_15_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__55426\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37377\,
            lcout => \comm_spi.data_tx_7__N_763\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i19179_4_lut_3_lut_LC_15_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__37378\,
            in1 => \N__37718\,
            in2 => \_gnd_net_\,
            in3 => \N__55427\,
            lcout => \comm_spi.n22644\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_88_2_lut_LC_15_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__55423\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37356\,
            lcout => \comm_spi.imosi_N_744\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_89_2_lut_LC_15_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__37357\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55422\,
            lcout => \comm_spi.imosi_N_745\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_95_2_lut_LC_15_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__55425\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53164\,
            lcout => \comm_spi.data_tx_7__N_761\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i3_12209_12210_reset_LC_15_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__37719\,
            in1 => \N__37662\,
            in2 => \_gnd_net_\,
            in3 => \N__37689\,
            lcout => \comm_spi.n14612\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52407\,
            ce => 'H',
            sr => \N__37702\
        );

    \comm_spi.data_tx_i2_12205_12206_reset_LC_15_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50220\,
            in1 => \N__52468\,
            in2 => \_gnd_net_\,
            in3 => \N__52518\,
            lcout => \comm_spi.n14608\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52424\,
            ce => 'H',
            sr => \N__37678\
        );

    \comm_spi.data_tx_i2_12205_12206_set_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__50221\,
            in1 => \N__52461\,
            in2 => \_gnd_net_\,
            in3 => \N__52522\,
            lcout => \comm_spi.n14607\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52442\,
            ce => 'H',
            sr => \N__37645\
        );

    \comm_spi.i19184_4_lut_3_lut_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__55429\,
            in1 => \N__37633\,
            in2 => \_gnd_net_\,
            in3 => \N__46191\,
            lcout => \comm_spi.n22641\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i19189_4_lut_3_lut_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__46257\,
            in1 => \N__53160\,
            in2 => \_gnd_net_\,
            in3 => \N__55430\,
            lcout => \comm_spi.n22638\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15011_2_lut_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__41169\,
            in1 => \_gnd_net_\,
            in2 => \N__41197\,
            in3 => \_gnd_net_\,
            lcout => n17393,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18832_2_lut_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37606\,
            in2 => \_gnd_net_\,
            in3 => \N__38897\,
            lcout => n21067,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_4_lut_adj_229_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111011101"
        )
    port map (
            in0 => \N__51239\,
            in1 => \N__54486\,
            in2 => \N__54001\,
            in3 => \N__37516\,
            lcout => OPEN,
            ltout => \n11839_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_152_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010000000"
        )
    port map (
            in0 => \N__46500\,
            in1 => \N__49216\,
            in2 => \N__37909\,
            in3 => \N__37905\,
            lcout => n11846,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_284_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000001000000"
        )
    port map (
            in0 => \N__51240\,
            in1 => \N__37906\,
            in2 => \N__49235\,
            in3 => \N__54487\,
            lcout => n14722,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6817_2_lut_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__53838\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53487\,
            lcout => n9222,
            ltout => \n9222_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_303_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010001000"
        )
    port map (
            in0 => \N__49215\,
            in1 => \N__54485\,
            in2 => \N__37894\,
            in3 => \N__51238\,
            lcout => n12322,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i41_4_lut_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000101100"
        )
    port map (
            in0 => \N__56945\,
            in1 => \N__47851\,
            in2 => \N__57447\,
            in3 => \N__56270\,
            lcout => OPEN,
            ltout => \n24_adj_1579_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18910_2_lut_LC_15_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__37891\,
            in3 => \N__44401\,
            lcout => OPEN,
            ltout => \n21079_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i42_4_lut_LC_15_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__53839\,
            in1 => \N__50078\,
            in2 => \N__37888\,
            in3 => \N__46581\,
            lcout => n16_adj_1570,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15209_2_lut_3_lut_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__53874\,
            in1 => \N__43347\,
            in2 => \_gnd_net_\,
            in3 => \N__51207\,
            lcout => n14_adj_1529,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.cmd_rdadctmp_i15_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110001000100010"
        )
    port map (
            in0 => \N__45179\,
            in1 => \N__37871\,
            in2 => \N__48358\,
            in3 => \N__38767\,
            lcout => cmd_rdadctmp_15_adj_1428,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55120\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_291_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010001000"
        )
    port map (
            in0 => \N__49910\,
            in1 => \N__49860\,
            in2 => \N__53521\,
            in3 => \N__38131\,
            lcout => n12080,
            ltout => \n12080_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12352_2_lut_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__38125\,
            in3 => \N__54488\,
            lcout => n14749,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22129_bdd_4_lut_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010000"
        )
    port map (
            in0 => \N__49523\,
            in1 => \N__38122\,
            in2 => \N__43525\,
            in3 => \N__38047\,
            lcout => n22132,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_299_LC_15_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__49859\,
            in1 => \N__49909\,
            in2 => \_gnd_net_\,
            in3 => \N__51454\,
            lcout => n12206,
            ltout => \n12206_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12373_2_lut_LC_15_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__54489\,
            in1 => \_gnd_net_\,
            in2 => \N__38095\,
            in3 => \_gnd_net_\,
            lcout => n14770,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_2__bdd_4_lut_LC_15_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010101010"
        )
    port map (
            in0 => \N__50087\,
            in1 => \N__38083\,
            in2 => \N__38056\,
            in3 => \N__49522\,
            lcout => n22129,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_5_i22_3_lut_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__49077\,
            in1 => \N__38275\,
            in2 => \_gnd_net_\,
            in3 => \N__47848\,
            lcout => OPEN,
            ltout => \n22_adj_1599_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_5_i30_3_lut_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__38041\,
            in1 => \_gnd_net_\,
            in2 => \N__38029\,
            in3 => \N__56259\,
            lcout => OPEN,
            ltout => \n30_adj_1600_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_buf_2__i5_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54033\,
            in2 => \N__38026\,
            in3 => \N__37981\,
            lcout => comm_buf_2_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55129\,
            ce => \N__37920\,
            sr => \N__38346\
        );

    \mux_130_Mux_5_i19_3_lut_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__56953\,
            in1 => \N__38329\,
            in2 => \_gnd_net_\,
            in3 => \N__38303\,
            lcout => n19_adj_1598,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_2__bdd_4_lut_19491_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__38269\,
            in1 => \N__50088\,
            in2 => \N__38263\,
            in3 => \N__49524\,
            lcout => OPEN,
            ltout => \n22123_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n22123_bdd_4_lut_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010111100000"
        )
    port map (
            in0 => \N__49525\,
            in1 => \N__38242\,
            in2 => \N__38224\,
            in3 => \N__44871\,
            lcout => n22126,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_283_LC_15_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__38209\,
            in1 => \N__56952\,
            in2 => \_gnd_net_\,
            in3 => \N__56260\,
            lcout => n11324,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_272_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__53499\,
            in1 => \N__56258\,
            in2 => \_gnd_net_\,
            in3 => \N__38208\,
            lcout => n20613,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i2_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__43864\,
            in1 => \N__38719\,
            in2 => \N__52147\,
            in3 => \N__38162\,
            lcout => \SELIRNG0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55141\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i5_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__50136\,
            in1 => \N__42005\,
            in2 => \_gnd_net_\,
            in3 => \N__38417\,
            lcout => req_data_cnt_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55141\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15204_2_lut_3_lut_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__54027\,
            in1 => \N__51282\,
            in2 => \_gnd_net_\,
            in3 => \N__44108\,
            lcout => n14_adj_1552,
            ltout => \n14_adj_1552_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i9_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__42006\,
            in2 => \N__38134\,
            in3 => \N__41646\,
            lcout => req_data_cnt_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55141\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15202_2_lut_3_lut_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__43796\,
            in1 => \N__51283\,
            in2 => \_gnd_net_\,
            in3 => \N__53957\,
            lcout => n14_adj_1550,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15_4_lut_adj_315_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111101000111"
        )
    port map (
            in0 => \N__43299\,
            in1 => \N__54668\,
            in2 => \N__42353\,
            in3 => \N__52065\,
            lcout => n12254,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i15_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__42004\,
            in1 => \_gnd_net_\,
            in2 => \N__45768\,
            in3 => \N__41684\,
            lcout => req_data_cnt_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55141\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_290_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101010001000"
        )
    port map (
            in0 => \N__49858\,
            in1 => \N__49908\,
            in2 => \N__53532\,
            in3 => \N__40813\,
            lcout => n12007,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i4_LC_15_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38390\,
            in2 => \N__42025\,
            in3 => \N__38469\,
            lcout => req_data_cnt_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55154\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i1_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__38442\,
            in1 => \N__42019\,
            in2 => \_gnd_net_\,
            in3 => \N__38373\,
            lcout => req_data_cnt_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55154\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i4_4_lut_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__46852\,
            in1 => \N__46782\,
            in2 => \N__38418\,
            in3 => \N__38825\,
            lcout => n20_adj_1496,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_adj_69_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__46812\,
            in1 => \N__46912\,
            in2 => \N__38394\,
            in3 => \N__38372\,
            lcout => OPEN,
            ltout => \n18_adj_1553_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13_4_lut_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__38359\,
            in1 => \N__41875\,
            in2 => \N__38353\,
            in3 => \N__41698\,
            lcout => OPEN,
            ltout => \n29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_80_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38937\,
            in2 => \N__38902\,
            in3 => \N__42151\,
            lcout => n16_adj_1609,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i3_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__42020\,
            in1 => \N__38865\,
            in2 => \_gnd_net_\,
            in3 => \N__38826\,
            lcout => req_data_cnt_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55154\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5_4_lut_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__38812\,
            in1 => \N__38794\,
            in2 => \N__38613\,
            in3 => \N__44717\,
            lcout => n21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_6__I_0_363_i9_2_lut_3_lut_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__57548\,
            in1 => \N__56966\,
            in2 => \_gnd_net_\,
            in3 => \N__47843\,
            lcout => OPEN,
            ltout => \n9_adj_1408_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_271_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110100000000"
        )
    port map (
            in0 => \N__41622\,
            in1 => \N__51914\,
            in2 => \N__38770\,
            in3 => \N__54625\,
            lcout => n11901,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i12_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44718\,
            in1 => \N__42139\,
            in2 => \_gnd_net_\,
            in3 => \N__39315\,
            lcout => \acadc_skipCount_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55169\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i6_LC_15_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__48314\,
            in1 => \N__48504\,
            in2 => \N__38763\,
            in3 => \N__40853\,
            lcout => buf_adcdata_vac_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55169\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i10_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__38612\,
            in1 => \N__51978\,
            in2 => \N__38734\,
            in3 => \N__39316\,
            lcout => \acadc_skipCount_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55169\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i12_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__42024\,
            in1 => \_gnd_net_\,
            in2 => \N__42145\,
            in3 => \N__56397\,
            lcout => req_data_cnt_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55169\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acadc_skipCount_i11_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__51915\,
            in1 => \N__39317\,
            in2 => \N__43816\,
            in3 => \N__45470\,
            lcout => \acadc_skipCount_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55169\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_276_LC_15_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100010"
        )
    port map (
            in0 => \N__54624\,
            in1 => \N__45561\,
            in2 => \N__52062\,
            in3 => \N__45380\,
            lcout => n12367,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i4_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__54709\,
            in1 => \N__39043\,
            in2 => \N__52061\,
            in3 => \N__42490\,
            lcout => data_index_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55184\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_adj_84_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__53522\,
            in1 => \N__47835\,
            in2 => \N__39183\,
            in3 => \N__57395\,
            lcout => n8780,
            ltout => \n8780_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14930_3_lut_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41347\,
            in2 => \N__39160\,
            in3 => \N__42840\,
            lcout => n17314,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12226_2_lut_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__39150\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48631\,
            lcout => n14632,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i7_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__51951\,
            in1 => \N__39057\,
            in2 => \N__42615\,
            in3 => \N__45693\,
            lcout => buf_dds0_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55184\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6402_3_lut_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__46654\,
            in1 => \N__42508\,
            in2 => \_gnd_net_\,
            in3 => \N__43284\,
            lcout => n8_adj_1541,
            ltout => \n8_adj_1541_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_354_Mux_4_i15_4_lut_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__51950\,
            in1 => \N__54623\,
            in2 => \N__39037\,
            in3 => \N__42489\,
            lcout => \data_index_9_N_212_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_count_i0_i0_LC_15_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46986\,
            in2 => \N__40097\,
            in3 => \_gnd_net_\,
            lcout => data_count_0,
            ltout => OPEN,
            carryin => \bfn_15_17_0_\,
            carryout => n19287,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__48655\,
            sr => \N__48586\
        );

    \data_count_i0_i1_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39986\,
            in2 => \_gnd_net_\,
            in3 => \N__39967\,
            lcout => data_count_1,
            ltout => OPEN,
            carryin => n19287,
            carryout => n19288,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__48655\,
            sr => \N__48586\
        );

    \data_count_i0_i2_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39881\,
            in2 => \_gnd_net_\,
            in3 => \N__39859\,
            lcout => data_count_2,
            ltout => OPEN,
            carryin => n19288,
            carryout => n19289,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__48655\,
            sr => \N__48586\
        );

    \data_count_i0_i3_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39779\,
            in2 => \_gnd_net_\,
            in3 => \N__39757\,
            lcout => data_count_3,
            ltout => OPEN,
            carryin => n19289,
            carryout => n19290,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__48655\,
            sr => \N__48586\
        );

    \data_count_i0_i4_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39671\,
            in2 => \_gnd_net_\,
            in3 => \N__39649\,
            lcout => data_count_4,
            ltout => OPEN,
            carryin => n19290,
            carryout => n19291,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__48655\,
            sr => \N__48586\
        );

    \data_count_i0_i5_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39563\,
            in2 => \_gnd_net_\,
            in3 => \N__39541\,
            lcout => data_count_5,
            ltout => OPEN,
            carryin => n19291,
            carryout => n19292,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__48655\,
            sr => \N__48586\
        );

    \data_count_i0_i6_LC_15_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39458\,
            in2 => \_gnd_net_\,
            in3 => \N__39436\,
            lcout => data_count_6,
            ltout => OPEN,
            carryin => n19292,
            carryout => n19293,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__48655\,
            sr => \N__48586\
        );

    \data_count_i0_i7_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39356\,
            in2 => \_gnd_net_\,
            in3 => \N__39334\,
            lcout => data_count_7,
            ltout => OPEN,
            carryin => n19293,
            carryout => n19294,
            clk => \INVdata_count_i0_i0C_net\,
            ce => \N__48655\,
            sr => \N__48586\
        );

    \data_count_i0_i8_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40523\,
            in2 => \_gnd_net_\,
            in3 => \N__40501\,
            lcout => data_count_8,
            ltout => OPEN,
            carryin => \bfn_15_18_0_\,
            carryout => n19295,
            clk => \INVdata_count_i0_i8C_net\,
            ce => \N__48663\,
            sr => \N__48596\
        );

    \data_count_i0_i9_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40412\,
            in2 => \_gnd_net_\,
            in3 => \N__40498\,
            lcout => data_count_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVdata_count_i0_i8C_net\,
            ce => \N__48663\,
            sr => \N__48596\
        );

    \SIG_DDS.tmp_buf_i15_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__55872\,
            in1 => \N__55634\,
            in2 => \N__40390\,
            in3 => \N__45591\,
            lcout => tmp_buf_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55221\,
            ce => \N__40316\,
            sr => \_gnd_net_\
        );

    \SIG_DDS.tmp_buf_i0_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__55871\,
            in1 => \N__55633\,
            in2 => \N__42916\,
            in3 => \N__40375\,
            lcout => \SIG_DDS.tmp_buf_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55221\,
            ce => \N__40316\,
            sr => \_gnd_net_\
        );

    \comm_spi.i19199_4_lut_3_lut_LC_16_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__40229\,
            in1 => \N__40288\,
            in2 => \_gnd_net_\,
            in3 => \N__55472\,
            lcout => \comm_spi.n22623\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i7_12190_12191_set_LC_16_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__40230\,
            in1 => \N__43546\,
            in2 => \_gnd_net_\,
            in3 => \N__43641\,
            lcout => \comm_spi.n14592\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52319\,
            ce => 'H',
            sr => \N__40260\
        );

    \comm_spi.data_tx_i7_12190_12191_reset_LC_16_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__43645\,
            in1 => \N__40234\,
            in2 => \_gnd_net_\,
            in3 => \N__43545\,
            lcout => \comm_spi.n14593\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52391\,
            ce => 'H',
            sr => \N__44233\
        );

    \comm_spi.imiso_83_12193_12194_reset_LC_16_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40209\,
            in1 => \N__40185\,
            in2 => \_gnd_net_\,
            in3 => \N__44283\,
            lcout => \comm_spi.n14596\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.imiso_83_12193_12194_resetC_net\,
            ce => 'H',
            sr => \N__44232\
        );

    \clk_cnt_3761_3762__i2_LC_16_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__41165\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41189\,
            lcout => clk_cnt_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56024\,
            ce => 'H',
            sr => \N__40723\
        );

    \clk_cnt_3761_3762__i1_LC_16_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41164\,
            lcout => clk_cnt_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56024\,
            ce => 'H',
            sr => \N__40723\
        );

    \i1_4_lut_adj_162_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100010"
        )
    port map (
            in0 => \N__44418\,
            in1 => \N__57547\,
            in2 => \N__40711\,
            in3 => \N__47833\,
            lcout => \comm_state_3_N_412_3\,
            ltout => \comm_state_3_N_412_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18743_2_lut_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__53491\,
            in1 => \_gnd_net_\,
            in2 => \N__40690\,
            in3 => \_gnd_net_\,
            lcout => n21162,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15273_2_lut_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__53686\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53489\,
            lcout => n17656,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18105_2_lut_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__53490\,
            in1 => \N__53685\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \n20700_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_273_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000010"
        )
    port map (
            in0 => \N__49210\,
            in1 => \N__51197\,
            in2 => \N__40687\,
            in3 => \N__54367\,
            lcout => n11411,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \flagcntwd_303_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110111011101"
        )
    port map (
            in0 => \N__53492\,
            in1 => \N__53687\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => flagcntwd,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55100\,
            ce => \N__40660\,
            sr => \N__40648\
        );

    \i1_2_lut_adj_249_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51196\,
            in2 => \_gnd_net_\,
            in3 => \N__53488\,
            lcout => n11333,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i11_4_lut_adj_223_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__44487\,
            in1 => \N__44631\,
            in2 => \N__44689\,
            in3 => \N__44539\,
            lcout => n27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15200_2_lut_3_lut_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__53871\,
            in1 => \N__40784\,
            in2 => \_gnd_net_\,
            in3 => \N__51106\,
            lcout => n14_adj_1548,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15201_2_lut_3_lut_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__46700\,
            in1 => \N__51074\,
            in2 => \_gnd_net_\,
            in3 => \N__53872\,
            lcout => n14_adj_1549,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i9_4_lut_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__44616\,
            in1 => \N__44454\,
            in2 => \N__44572\,
            in3 => \N__44506\,
            lcout => n25_adj_1616,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18268_3_lut_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001010101"
        )
    port map (
            in0 => \N__53494\,
            in1 => \N__49790\,
            in2 => \_gnd_net_\,
            in3 => \N__53873\,
            lcout => n20863,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_LC_16_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__49791\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53493\,
            lcout => n14514,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_73_LC_16_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001000"
        )
    port map (
            in0 => \N__49211\,
            in1 => \N__54372\,
            in2 => \_gnd_net_\,
            in3 => \N__51073\,
            lcout => n20556,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12_4_lut_adj_221_LC_16_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__44586\,
            in1 => \N__44953\,
            in2 => \N__44671\,
            in3 => \N__44520\,
            lcout => n28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10_4_lut_adj_222_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__44553\,
            in1 => \N__44601\,
            in2 => \N__44650\,
            in3 => \N__44473\,
            lcout => OPEN,
            ltout => \n26_adj_1625_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15_4_lut_adj_227_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__40747\,
            in1 => \N__40741\,
            in2 => \N__40735\,
            in3 => \N__40732\,
            lcout => OPEN,
            ltout => \n19553_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7_4_lut_adj_228_LC_16_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__44931\,
            in1 => \N__53038\,
            in2 => \N__40726\,
            in3 => \N__41203\,
            lcout => n14700,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12387_3_lut_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010101010"
        )
    port map (
            in0 => \N__47081\,
            in1 => \N__54537\,
            in2 => \_gnd_net_\,
            in3 => \N__49302\,
            lcout => n14784,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_6_i22_3_lut_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__48564\,
            in1 => \N__40831\,
            in2 => \_gnd_net_\,
            in3 => \N__47832\,
            lcout => n22_adj_1594,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_adj_225_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__44703\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44967\,
            lcout => n10_adj_1582,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_RTD_287_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__40961\,
            in1 => \N__41196\,
            in2 => \_gnd_net_\,
            in3 => \N__41170\,
            lcout => \clk_RTD\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56026\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SecClk_292_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40906\,
            in2 => \_gnd_net_\,
            in3 => \N__44902\,
            lcout => \TEST_LED\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56026\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_6_i19_3_lut_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__40888\,
            in1 => \N__40860\,
            in2 => \_gnd_net_\,
            in3 => \N__56939\,
            lcout => n19_adj_1593,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i45_4_lut_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000100000"
        )
    port map (
            in0 => \N__44411\,
            in1 => \N__53837\,
            in2 => \N__40825\,
            in3 => \N__46996\,
            lcout => n20_adj_1607,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_2_lut_3_lut_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__56940\,
            in1 => \N__57543\,
            in2 => \_gnd_net_\,
            in3 => \N__47754\,
            lcout => n10553,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_137_Mux_4_i4_3_lut_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__40804\,
            in1 => \N__51579\,
            in2 => \_gnd_net_\,
            in3 => \N__40795\,
            lcout => n4_adj_1566,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18184_3_lut_LC_16_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__56938\,
            in1 => \N__41469\,
            in2 => \_gnd_net_\,
            in3 => \N__47343\,
            lcout => n20779,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_57_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011010000"
        )
    port map (
            in0 => \N__45562\,
            in1 => \N__52063\,
            in2 => \N__54669\,
            in3 => \N__41615\,
            lcout => n12415,
            ltout => \n12415_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i6_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__51376\,
            in1 => \_gnd_net_\,
            in2 => \N__41440\,
            in3 => \N__41718\,
            lcout => req_data_cnt_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55142\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i5_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__45292\,
            in1 => \N__44800\,
            in2 => \_gnd_net_\,
            in3 => \N__41386\,
            lcout => \buf_cfgRTD_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55142\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i13_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__44799\,
            in1 => \N__41987\,
            in2 => \_gnd_net_\,
            in3 => \N__45087\,
            lcout => req_data_cnt_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55142\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i0_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__41990\,
            in1 => \N__52064\,
            in2 => \N__41363\,
            in3 => \N__41744\,
            lcout => req_data_cnt_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55142\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i2_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__41284\,
            in1 => \N__41988\,
            in2 => \_gnd_net_\,
            in3 => \N__41591\,
            lcout => req_data_cnt_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55142\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i7_LC_16_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__41989\,
            in1 => \N__41263\,
            in2 => \_gnd_net_\,
            in3 => \N__41565\,
            lcout => req_data_cnt_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55142\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1536244_i1_3_lut_LC_16_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__45028\,
            in1 => \N__41242\,
            in2 => \_gnd_net_\,
            in3 => \N__56315\,
            lcout => n30_adj_1520,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i11_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__41992\,
            in1 => \N__43802\,
            in2 => \N__52158\,
            in3 => \N__45255\,
            lcout => req_data_cnt_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55155\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i8_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__41782\,
            in1 => \N__41991\,
            in2 => \_gnd_net_\,
            in3 => \N__41895\,
            lcout => req_data_cnt_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55155\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_74_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__46936\,
            in1 => \N__47412\,
            in2 => \N__41751\,
            in3 => \N__41714\,
            lcout => n17_adj_1554,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i8_4_lut_adj_55_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__48682\,
            in1 => \N__47307\,
            in2 => \N__41691\,
            in3 => \N__41642\,
            lcout => n24_adj_1530,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_4_lut_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__56803\,
            in1 => \N__47790\,
            in2 => \N__57533\,
            in3 => \N__41614\,
            lcout => n10540,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6_4_lut_adj_56_LC_16_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__46881\,
            in1 => \N__47377\,
            in2 => \N__41592\,
            in3 => \N__41561\,
            lcout => n22_adj_1492,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_adj_313_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111011"
        )
    port map (
            in0 => \N__51659\,
            in1 => \N__51200\,
            in2 => \_gnd_net_\,
            in3 => \N__53956\,
            lcout => n10579,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i14_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__41506\,
            in1 => \N__42008\,
            in2 => \_gnd_net_\,
            in3 => \N__45231\,
            lcout => req_data_cnt_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55170\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5_4_lut_adj_59_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__47221\,
            in1 => \N__41912\,
            in2 => \N__47278\,
            in3 => \N__56387\,
            lcout => OPEN,
            ltout => \n21_adj_1494_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14_4_lut_adj_79_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__42169\,
            in1 => \N__45211\,
            in2 => \N__42160\,
            in3 => \N__42157\,
            lcout => n30_adj_1597,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_cfgRTD_i4_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__42119\,
            in1 => \N__45279\,
            in2 => \_gnd_net_\,
            in3 => \N__42044\,
            lcout => \buf_cfgRTD_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55170\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \req_data_cnt_i10_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__41913\,
            in1 => \N__42007\,
            in2 => \_gnd_net_\,
            in3 => \N__41950\,
            lcout => req_data_cnt_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55170\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__47200\,
            in1 => \N__47344\,
            in2 => \N__45091\,
            in3 => \N__41891\,
            lcout => n19_adj_1499,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_125_2_lut_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__42841\,
            in1 => \N__42839\,
            in2 => \N__42339\,
            in3 => \N__41869\,
            lcout => n7_adj_1515,
            ltout => OPEN,
            carryin => \bfn_16_15_0_\,
            carryout => n19326,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_125_3_lut_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__43321\,
            in1 => \N__43320\,
            in2 => \N__42343\,
            in3 => \N__41866\,
            lcout => n7_adj_1546,
            ltout => OPEN,
            carryin => n19326,
            carryout => n19327,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_125_4_lut_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__41863\,
            in1 => \N__41862\,
            in2 => \N__42340\,
            in3 => \N__41830\,
            lcout => n7_adj_1544,
            ltout => OPEN,
            carryin => n19327,
            carryout => n19328,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_125_5_lut_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__41826\,
            in1 => \N__41825\,
            in2 => \N__42344\,
            in3 => \N__41785\,
            lcout => n7_adj_1542,
            ltout => OPEN,
            carryin => n19328,
            carryout => n19329,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_125_6_lut_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__42507\,
            in1 => \N__42506\,
            in2 => \N__42341\,
            in3 => \N__42481\,
            lcout => n7_adj_1540,
            ltout => OPEN,
            carryin => n19329,
            carryout => n19330,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_125_7_lut_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__46038\,
            in1 => \N__46037\,
            in2 => \N__42345\,
            in3 => \N__42478\,
            lcout => n17336,
            ltout => OPEN,
            carryin => n19330,
            carryout => n19331,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_125_8_lut_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__42679\,
            in1 => \N__42678\,
            in2 => \N__42342\,
            in3 => \N__42475\,
            lcout => n7_adj_1537,
            ltout => OPEN,
            carryin => n19331,
            carryout => n19332,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_125_9_lut_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__42472\,
            in1 => \N__42471\,
            in2 => \N__42346\,
            in3 => \N__42412\,
            lcout => n7_adj_1535,
            ltout => OPEN,
            carryin => n19332,
            carryout => n19333,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_125_10_lut_LC_16_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__42409\,
            in1 => \N__42408\,
            in2 => \N__42358\,
            in3 => \N__42361\,
            lcout => n7_adj_1533,
            ltout => OPEN,
            carryin => \bfn_16_16_0_\,
            carryout => n19334,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_125_11_lut_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001110101100"
        )
    port map (
            in0 => \N__42725\,
            in1 => \N__42726\,
            in2 => \N__42357\,
            in3 => \N__42268\,
            lcout => n7_adj_1531,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i9_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__54635\,
            in1 => \N__43038\,
            in2 => \N__52033\,
            in3 => \N__43023\,
            lcout => data_index_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55199\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14955_3_lut_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__50183\,
            in1 => \N__46042\,
            in2 => \_gnd_net_\,
            in3 => \N__43275\,
            lcout => n17338,
            ltout => \n17338_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14957_4_lut_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__51920\,
            in1 => \N__54610\,
            in2 => \N__42265\,
            in3 => \N__46053\,
            lcout => \data_index_9_N_212_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i0_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__54611\,
            in1 => \N__42873\,
            in2 => \N__52077\,
            in3 => \N__42855\,
            lcout => data_index_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55199\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i2_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__45697\,
            in1 => \N__51979\,
            in2 => \N__42822\,
            in3 => \N__42746\,
            lcout => buf_dds0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55199\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6352_3_lut_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44107\,
            in1 => \N__42727\,
            in2 => \_gnd_net_\,
            in3 => \N__43274\,
            lcout => n8_adj_1532,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i4_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__51975\,
            in1 => \N__42701\,
            in2 => \N__46665\,
            in3 => \N__45675\,
            lcout => buf_dds0_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55212\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6382_3_lut_LC_16_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__51431\,
            in1 => \N__42677\,
            in2 => \_gnd_net_\,
            in3 => \N__43276\,
            lcout => n8_adj_1538,
            ltout => \n8_adj_1538_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i6_LC_16_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__51976\,
            in1 => \N__54705\,
            in2 => \N__42682\,
            in3 => \N__43981\,
            lcout => data_index_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55212\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i6_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__45676\,
            in1 => \N__51977\,
            in2 => \N__51438\,
            in3 => \N__42644\,
            lcout => buf_dds0_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55212\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds1_i7_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010001000"
        )
    port map (
            in0 => \N__45965\,
            in1 => \N__42530\,
            in2 => \N__42625\,
            in3 => \N__45829\,
            lcout => buf_dds1_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55212\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i0_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__51974\,
            in1 => \N__43865\,
            in2 => \N__43532\,
            in3 => \N__50285\,
            lcout => buf_control_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55212\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i1_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__54704\,
            in1 => \N__43228\,
            in2 => \N__52043\,
            in3 => \N__43219\,
            lcout => data_index_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55222\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i8_LC_16_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__45696\,
            in1 => \N__43524\,
            in2 => \N__52042\,
            in3 => \N__43409\,
            lcout => buf_dds0_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55222\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6432_3_lut_LC_16_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__43375\,
            in1 => \N__43319\,
            in2 => \_gnd_net_\,
            in3 => \N__43291\,
            lcout => n8_adj_1547,
            ltout => \n8_adj_1547_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_354_Mux_1_i15_4_lut_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__51929\,
            in1 => \N__54597\,
            in2 => \N__43222\,
            in3 => \N__43218\,
            lcout => \data_index_9_N_212_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i11_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__43821\,
            in1 => \N__45694\,
            in2 => \N__43097\,
            in3 => \N__51930\,
            lcout => buf_dds0_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55222\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i5_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111010100100000"
        )
    port map (
            in0 => \N__45695\,
            in1 => \N__51983\,
            in2 => \N__50190\,
            in3 => \N__43055\,
            lcout => buf_dds0_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55222\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_354_Mux_9_i15_4_lut_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__54703\,
            in1 => \N__43039\,
            in2 => \N__52124\,
            in3 => \N__43024\,
            lcout => \data_index_9_N_212_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.MOSI_31_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__42915\,
            in1 => \N__42885\,
            in2 => \_gnd_net_\,
            in3 => \N__55566\,
            lcout => \DDS_MOSI\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55231\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i1_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__52059\,
            in1 => \N__43872\,
            in2 => \N__44147\,
            in3 => \N__44009\,
            lcout => \DDS_RNG_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55231\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_354_Mux_6_i15_4_lut_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__54702\,
            in1 => \N__43990\,
            in2 => \N__52123\,
            in3 => \N__43980\,
            lcout => \data_index_9_N_212_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_control_i3_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111001101000000"
        )
    port map (
            in0 => \N__52060\,
            in1 => \N__43873\,
            in2 => \N__43822\,
            in3 => \N__45497\,
            lcout => \SELIRNG1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55231\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.bit_cnt_i0_LC_16_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001011010"
        )
    port map (
            in0 => \N__55567\,
            in1 => \_gnd_net_\,
            in2 => \N__43673\,
            in3 => \N__43710\,
            lcout => bit_cnt_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55231\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i6_12221_12222_reset_LC_17_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43573\,
            in1 => \N__46246\,
            in2 => \_gnd_net_\,
            in3 => \N__46293\,
            lcout => \comm_spi.n14624\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52416\,
            ce => 'H',
            sr => \N__43630\
        );

    \comm_spi.i19154_4_lut_3_lut_LC_17_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__52960\,
            in1 => \N__43612\,
            in2 => \_gnd_net_\,
            in3 => \N__55428\,
            lcout => \comm_spi.n22626\,
            ltout => \comm_spi.n22626_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i12181_3_lut_LC_17_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52969\,
            in2 => \N__43606\,
            in3 => \N__48769\,
            lcout => \comm_spi.iclk\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.i12189_3_lut_LC_17_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__44287\,
            in1 => \N__44242\,
            in2 => \_gnd_net_\,
            in3 => \N__43603\,
            lcout => \ICE_SPI_MISO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i6_12221_12222_set_LC_17_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__43569\,
            in1 => \N__46242\,
            in2 => \_gnd_net_\,
            in3 => \N__46294\,
            lcout => \comm_spi.n14623\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52379\,
            ce => 'H',
            sr => \N__44341\
        );

    \comm_spi.MISO_48_12187_12188_reset_LC_17_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__44322\,
            in1 => \N__44311\,
            in2 => \_gnd_net_\,
            in3 => \N__44282\,
            lcout => \comm_spi.n14590\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.MISO_48_12187_12188_resetC_net\,
            ce => 'H',
            sr => \N__44231\
        );

    \comm_state_i1_LC_17_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__54249\,
            in1 => \N__44428\,
            in2 => \N__52113\,
            in3 => \N__44179\,
            lcout => comm_state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55101\,
            ce => \N__44161\,
            sr => \_gnd_net_\
        );

    \comm_state_1__bdd_4_lut_LC_17_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010010101010"
        )
    port map (
            in0 => \N__53681\,
            in1 => \N__44197\,
            in2 => \N__52232\,
            in3 => \N__51110\,
            lcout => OPEN,
            ltout => \n21913_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n21913_bdd_4_lut_LC_17_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__51111\,
            in1 => \N__53498\,
            in2 => \N__44182\,
            in3 => \N__44170\,
            lcout => n21916,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i227_2_lut_LC_17_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49800\,
            in2 => \_gnd_net_\,
            in3 => \N__49641\,
            lcout => n1252,
            ltout => \n1252_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_342_Mux_1_i2_3_lut_4_lut_LC_17_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__49798\,
            in1 => \N__53680\,
            in2 => \N__44173\,
            in3 => \N__53495\,
            lcout => n2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19013_4_lut_LC_17_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010101000000"
        )
    port map (
            in0 => \N__53679\,
            in1 => \N__49113\,
            in2 => \N__51199\,
            in3 => \N__49799\,
            lcout => OPEN,
            ltout => \n21088_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19124_4_lut_LC_17_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111011101"
        )
    port map (
            in0 => \N__46303\,
            in1 => \N__54245\,
            in2 => \N__44164\,
            in3 => \N__53496\,
            lcout => n14_adj_1497,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_3__I_0_342_Mux_1_i8_3_lut_4_lut_LC_17_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000110110001"
        )
    port map (
            in0 => \N__53497\,
            in1 => \N__44440\,
            in2 => \N__53830\,
            in3 => \N__44434\,
            lcout => n8_adj_1555,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i458_2_lut_LC_17_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__49755\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__49632\,
            lcout => n2342,
            ltout => \n2342_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i32_4_lut_LC_17_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011000000"
        )
    port map (
            in0 => \N__51198\,
            in1 => \N__53658\,
            in2 => \N__44422\,
            in3 => \N__44419\,
            lcout => OPEN,
            ltout => \n15_adj_1602_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_i2_LC_17_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011111000"
        )
    port map (
            in0 => \N__44371\,
            in1 => \N__44362\,
            in2 => \N__44374\,
            in3 => \N__53512\,
            lcout => comm_state_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55109\,
            ce => \N__49555\,
            sr => \N__54609\
        );

    \i1_2_lut_adj_277_LC_17_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49751\,
            in2 => \_gnd_net_\,
            in3 => \N__51105\,
            lcout => n20571,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_4_lut_adj_254_LC_17_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111101"
        )
    port map (
            in0 => \N__53656\,
            in1 => \N__49492\,
            in2 => \N__49348\,
            in3 => \N__49324\,
            lcout => n20641,
            ltout => \n20641_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i33_3_lut_LC_17_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__53511\,
            in1 => \N__53657\,
            in2 => \N__44365\,
            in3 => \_gnd_net_\,
            lcout => n12_adj_1603,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i22_4_lut_4_lut_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011001000100"
        )
    port map (
            in0 => \N__53655\,
            in1 => \N__53510\,
            in2 => \N__49782\,
            in3 => \N__49633\,
            lcout => n7_adj_1588,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_312_LC_17_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__54238\,
            in1 => \N__53654\,
            in2 => \_gnd_net_\,
            in3 => \N__51104\,
            lcout => n20650,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \secclk_cnt_3765_3766__i1_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44587\,
            in2 => \_gnd_net_\,
            in3 => \N__44575\,
            lcout => secclk_cnt_0,
            ltout => OPEN,
            carryin => \bfn_17_9_0_\,
            carryout => n19447,
            clk => \N__56025\,
            ce => 'H',
            sr => \N__44910\
        );

    \secclk_cnt_3765_3766__i2_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44571\,
            in2 => \_gnd_net_\,
            in3 => \N__44557\,
            lcout => secclk_cnt_1,
            ltout => OPEN,
            carryin => n19447,
            carryout => n19448,
            clk => \N__56025\,
            ce => 'H',
            sr => \N__44910\
        );

    \secclk_cnt_3765_3766__i3_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44554\,
            in2 => \_gnd_net_\,
            in3 => \N__44542\,
            lcout => secclk_cnt_2,
            ltout => OPEN,
            carryin => n19448,
            carryout => n19449,
            clk => \N__56025\,
            ce => 'H',
            sr => \N__44910\
        );

    \secclk_cnt_3765_3766__i4_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44535\,
            in2 => \_gnd_net_\,
            in3 => \N__44524\,
            lcout => secclk_cnt_3,
            ltout => OPEN,
            carryin => n19449,
            carryout => n19450,
            clk => \N__56025\,
            ce => 'H',
            sr => \N__44910\
        );

    \secclk_cnt_3765_3766__i5_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44521\,
            in2 => \_gnd_net_\,
            in3 => \N__44509\,
            lcout => secclk_cnt_4,
            ltout => OPEN,
            carryin => n19450,
            carryout => n19451,
            clk => \N__56025\,
            ce => 'H',
            sr => \N__44910\
        );

    \secclk_cnt_3765_3766__i6_LC_17_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44505\,
            in2 => \_gnd_net_\,
            in3 => \N__44491\,
            lcout => secclk_cnt_5,
            ltout => OPEN,
            carryin => n19451,
            carryout => n19452,
            clk => \N__56025\,
            ce => 'H',
            sr => \N__44910\
        );

    \secclk_cnt_3765_3766__i7_LC_17_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44488\,
            in2 => \_gnd_net_\,
            in3 => \N__44476\,
            lcout => secclk_cnt_6,
            ltout => OPEN,
            carryin => n19452,
            carryout => n19453,
            clk => \N__56025\,
            ce => 'H',
            sr => \N__44910\
        );

    \secclk_cnt_3765_3766__i8_LC_17_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44472\,
            in2 => \_gnd_net_\,
            in3 => \N__44458\,
            lcout => secclk_cnt_7,
            ltout => OPEN,
            carryin => n19453,
            carryout => n19454,
            clk => \N__56025\,
            ce => 'H',
            sr => \N__44910\
        );

    \secclk_cnt_3765_3766__i9_LC_17_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44455\,
            in2 => \_gnd_net_\,
            in3 => \N__44443\,
            lcout => secclk_cnt_8,
            ltout => OPEN,
            carryin => \bfn_17_10_0_\,
            carryout => n19455,
            clk => \N__56027\,
            ce => 'H',
            sr => \N__44906\
        );

    \secclk_cnt_3765_3766__i10_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44704\,
            in2 => \_gnd_net_\,
            in3 => \N__44692\,
            lcout => secclk_cnt_9,
            ltout => OPEN,
            carryin => n19455,
            carryout => n19456,
            clk => \N__56027\,
            ce => 'H',
            sr => \N__44906\
        );

    \secclk_cnt_3765_3766__i11_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44688\,
            in2 => \_gnd_net_\,
            in3 => \N__44674\,
            lcout => secclk_cnt_10,
            ltout => OPEN,
            carryin => n19456,
            carryout => n19457,
            clk => \N__56027\,
            ce => 'H',
            sr => \N__44906\
        );

    \secclk_cnt_3765_3766__i12_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44670\,
            in2 => \_gnd_net_\,
            in3 => \N__44656\,
            lcout => secclk_cnt_11,
            ltout => OPEN,
            carryin => n19457,
            carryout => n19458,
            clk => \N__56027\,
            ce => 'H',
            sr => \N__44906\
        );

    \secclk_cnt_3765_3766__i13_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53067\,
            in2 => \_gnd_net_\,
            in3 => \N__44653\,
            lcout => secclk_cnt_12,
            ltout => OPEN,
            carryin => n19458,
            carryout => n19459,
            clk => \N__56027\,
            ce => 'H',
            sr => \N__44906\
        );

    \secclk_cnt_3765_3766__i14_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44649\,
            in2 => \_gnd_net_\,
            in3 => \N__44635\,
            lcout => secclk_cnt_13,
            ltout => OPEN,
            carryin => n19459,
            carryout => n19460,
            clk => \N__56027\,
            ce => 'H',
            sr => \N__44906\
        );

    \secclk_cnt_3765_3766__i15_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44632\,
            in2 => \_gnd_net_\,
            in3 => \N__44620\,
            lcout => secclk_cnt_14,
            ltout => OPEN,
            carryin => n19460,
            carryout => n19461,
            clk => \N__56027\,
            ce => 'H',
            sr => \N__44906\
        );

    \secclk_cnt_3765_3766__i16_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44617\,
            in2 => \_gnd_net_\,
            in3 => \N__44605\,
            lcout => secclk_cnt_15,
            ltout => OPEN,
            carryin => n19461,
            carryout => n19462,
            clk => \N__56027\,
            ce => 'H',
            sr => \N__44906\
        );

    \secclk_cnt_3765_3766__i17_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44602\,
            in2 => \_gnd_net_\,
            in3 => \N__44590\,
            lcout => secclk_cnt_16,
            ltout => OPEN,
            carryin => \bfn_17_11_0_\,
            carryout => n19463,
            clk => \N__56028\,
            ce => 'H',
            sr => \N__44911\
        );

    \secclk_cnt_3765_3766__i18_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44968\,
            in2 => \_gnd_net_\,
            in3 => \N__44956\,
            lcout => secclk_cnt_17,
            ltout => OPEN,
            carryin => n19463,
            carryout => n19464,
            clk => \N__56028\,
            ce => 'H',
            sr => \N__44911\
        );

    \secclk_cnt_3765_3766__i19_LC_17_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44952\,
            in2 => \_gnd_net_\,
            in3 => \N__44938\,
            lcout => secclk_cnt_18,
            ltout => OPEN,
            carryin => n19464,
            carryout => n19465,
            clk => \N__56028\,
            ce => 'H',
            sr => \N__44911\
        );

    \secclk_cnt_3765_3766__i20_LC_17_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53103\,
            in2 => \_gnd_net_\,
            in3 => \N__44935\,
            lcout => secclk_cnt_19,
            ltout => OPEN,
            carryin => n19465,
            carryout => n19466,
            clk => \N__56028\,
            ce => 'H',
            sr => \N__44911\
        );

    \secclk_cnt_3765_3766__i21_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44932\,
            in2 => \_gnd_net_\,
            in3 => \N__44920\,
            lcout => secclk_cnt_20,
            ltout => OPEN,
            carryin => n19466,
            carryout => n19467,
            clk => \N__56028\,
            ce => 'H',
            sr => \N__44911\
        );

    \secclk_cnt_3765_3766__i22_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53088\,
            in2 => \_gnd_net_\,
            in3 => \N__44917\,
            lcout => secclk_cnt_21,
            ltout => OPEN,
            carryin => n19467,
            carryout => n19468,
            clk => \N__56028\,
            ce => 'H',
            sr => \N__44911\
        );

    \secclk_cnt_3765_3766__i23_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53052\,
            in2 => \_gnd_net_\,
            in3 => \N__44914\,
            lcout => secclk_cnt_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__56028\,
            ce => 'H',
            sr => \N__44911\
        );

    \i1_2_lut_3_lut_adj_307_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__44872\,
            in1 => \N__51204\,
            in2 => \_gnd_net_\,
            in3 => \N__53828\,
            lcout => n14_adj_1556,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_4_i23_3_lut_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__44754\,
            in1 => \N__56927\,
            in2 => \_gnd_net_\,
            in3 => \N__44725\,
            lcout => n23_adj_1517,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_4_i22_3_lut_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__48828\,
            in1 => \N__51310\,
            in2 => \_gnd_net_\,
            in3 => \N__47825\,
            lcout => n22_adj_1606,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12250_3_lut_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__51205\,
            in1 => \N__54451\,
            in2 => \_gnd_net_\,
            in3 => \N__45431\,
            lcout => n14652,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18804_2_lut_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__56928\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45086\,
            lcout => n21022,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_317_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111011110"
        )
    port map (
            in0 => \N__45039\,
            in1 => \N__51578\,
            in2 => \N__50094\,
            in3 => \N__45445\,
            lcout => n4_adj_1576,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_length_i2_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__56929\,
            in1 => \N__45040\,
            in2 => \N__45058\,
            in3 => \N__45432\,
            lcout => comm_length_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55156\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_cmd_1__bdd_4_lut_19355_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101010001010"
        )
    port map (
            in0 => \N__57535\,
            in1 => \N__44998\,
            in2 => \N__47849\,
            in3 => \N__44974\,
            lcout => OPEN,
            ltout => \n21955_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \n21955_bdd_4_lut_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001011000010"
        )
    port map (
            in0 => \N__45451\,
            in1 => \N__47829\,
            in2 => \N__45031\,
            in3 => \N__45022\,
            lcout => n21958,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18787_2_lut_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__56932\,
            in1 => \N__45254\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n21024,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19055_2_lut_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45016\,
            in2 => \_gnd_net_\,
            in3 => \N__56931\,
            lcout => n20950,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_3_i26_3_lut_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__56930\,
            in1 => \N__44992\,
            in2 => \_gnd_net_\,
            in3 => \N__47240\,
            lcout => n26_adj_1519,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_128_Mux_3_i23_3_lut_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__45510\,
            in1 => \N__56933\,
            in2 => \_gnd_net_\,
            in3 => \N__45478\,
            lcout => n23_adj_1518,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_length_i0_LC_17_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001110100110"
        )
    port map (
            in0 => \N__57536\,
            in1 => \N__56311\,
            in2 => \N__56977\,
            in3 => \N__47831\,
            lcout => comm_length_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55171\,
            ce => \N__45439\,
            sr => \N__45403\
        );

    \comm_length_i1_LC_17_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011110011101111"
        )
    port map (
            in0 => \N__47830\,
            in1 => \N__56934\,
            in2 => \N__56341\,
            in3 => \N__57537\,
            lcout => comm_length_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55171\,
            ce => \N__45439\,
            sr => \N__45403\
        );

    \ADC_IAC.ADC_DATA_i7_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__49008\,
            in1 => \N__50962\,
            in2 => \N__47880\,
            in3 => \N__45155\,
            lcout => buf_adcdata_iac_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55185\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_280_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001010"
        )
    port map (
            in0 => \N__54441\,
            in1 => \N__51782\,
            in2 => \N__45394\,
            in3 => \N__45376\,
            lcout => n12381,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i7_4_lut_adj_58_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111110110111110"
        )
    port map (
            in0 => \N__48699\,
            in1 => \N__47241\,
            in2 => \N__45256\,
            in3 => \N__45227\,
            lcout => n23_adj_1491,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i7_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__48535\,
            in1 => \N__48347\,
            in2 => \N__45201\,
            in3 => \N__47928\,
            lcout => buf_adcdata_vac_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55185\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i15_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__50961\,
            in1 => \N__48798\,
            in2 => \N__45159\,
            in3 => \N__50519\,
            lcout => cmd_rdadctmp_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55185\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i16_LC_17_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110010001000100"
        )
    port map (
            in0 => \N__50518\,
            in1 => \N__45113\,
            in2 => \N__45163\,
            in3 => \N__50963\,
            lcout => cmd_rdadctmp_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55185\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i46_2_lut_LC_17_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49767\,
            in2 => \_gnd_net_\,
            in3 => \N__53987\,
            lcout => n23_adj_1574,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_index_i5_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010111100100000"
        )
    port map (
            in0 => \N__46060\,
            in1 => \N__51786\,
            in2 => \N__54599\,
            in3 => \N__46054\,
            lcout => data_index_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55200\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_4_lut_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000011111111"
        )
    port map (
            in0 => \N__51206\,
            in1 => \N__53829\,
            in2 => \N__54598\,
            in3 => \N__45810\,
            lcout => n16708,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15037_2_lut_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__53986\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53466\,
            lcout => n3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_4_lut_adj_243_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111111111111"
        )
    port map (
            in0 => \N__49801\,
            in1 => \N__54433\,
            in2 => \N__51259\,
            in3 => \N__49645\,
            lcout => n4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_251_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__49240\,
            in1 => \N__54440\,
            in2 => \N__50980\,
            in3 => \N__45933\,
            lcout => n11805,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf_dds0_i15_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__45767\,
            in1 => \N__45581\,
            in2 => \_gnd_net_\,
            in3 => \N__45674\,
            lcout => buf_dds0_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55223\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \equal_188_i9_2_lut_3_lut_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__57534\,
            in1 => \N__56989\,
            in2 => \_gnd_net_\,
            in3 => \N__47850\,
            lcout => n9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.dds_state_i1_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55862\,
            in2 => \_gnd_net_\,
            in3 => \N__55739\,
            lcout => dds_state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55232\,
            ce => \N__45534\,
            sr => \N__55659\
        );

    \comm_spi.data_tx_i5_12217_12218_reset_LC_18_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46273\,
            in1 => \N__46231\,
            in2 => \_gnd_net_\,
            in3 => \N__46138\,
            lcout => \comm_spi.n14620\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52417\,
            ce => 'H',
            sr => \N__46282\
        );

    \comm_spi.data_tx_i5_12217_12218_set_LC_18_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46269\,
            in1 => \N__46227\,
            in2 => \_gnd_net_\,
            in3 => \N__46137\,
            lcout => \comm_spi.n14619\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52426\,
            ce => 'H',
            sr => \N__48709\
        );

    \comm_spi.data_tx_i4_12213_12214_set_LC_18_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46207\,
            in1 => \N__46180\,
            in2 => \_gnd_net_\,
            in3 => \N__46159\,
            lcout => \comm_spi.n14615\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52360\,
            ce => 'H',
            sr => \N__46216\
        );

    \comm_spi.data_tx_i4_12213_12214_reset_LC_18_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__46206\,
            in1 => \N__46179\,
            in2 => \_gnd_net_\,
            in3 => \N__46155\,
            lcout => \comm_spi.n14616\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52430\,
            ce => 'H',
            sr => \N__53131\
        );

    \comm_state_3__I_0_342_Mux_3_i7_4_lut_LC_18_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011110000"
        )
    port map (
            in0 => \N__46120\,
            in1 => \N__52233\,
            in2 => \N__46111\,
            in3 => \N__51062\,
            lcout => OPEN,
            ltout => \n17658_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_i3_LC_18_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000001111"
        )
    port map (
            in0 => \N__51919\,
            in1 => \N__46096\,
            in2 => \N__46087\,
            in3 => \N__54176\,
            lcout => comm_state_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55121\,
            ce => \N__46453\,
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_260_LC_18_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__54175\,
            in1 => \N__51061\,
            in2 => \_gnd_net_\,
            in3 => \N__53637\,
            lcout => n12220,
            ltout => \n12220_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_LC_18_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011100000"
        )
    port map (
            in0 => \N__46084\,
            in1 => \N__46438\,
            in2 => \N__46063\,
            in3 => \N__46398\,
            lcout => OPEN,
            ltout => \n4_adj_1483_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_adj_52_LC_18_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010110000"
        )
    port map (
            in0 => \N__46467\,
            in1 => \N__49750\,
            in2 => \N__46510\,
            in3 => \N__46507\,
            lcout => n20510,
            ltout => \n20510_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_146_LC_18_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__46387\,
            in1 => \N__46483\,
            in2 => \N__46471\,
            in3 => \N__46468\,
            lcout => n20534,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_2_lut_3_lut_LC_18_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53474\,
            in2 => \N__49796\,
            in3 => \N__49626\,
            lcout => n11810,
            ltout => \n11810_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_LC_18_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010101010"
        )
    port map (
            in0 => \N__49140\,
            in1 => \_gnd_net_\,
            in2 => \N__46432\,
            in3 => \N__46399\,
            lcout => OPEN,
            ltout => \n20672_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_71_LC_18_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000000000000"
        )
    port map (
            in0 => \N__46422\,
            in1 => \N__49126\,
            in2 => \N__46408\,
            in3 => \N__46405\,
            lcout => n20536,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_306_LC_18_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53475\,
            in2 => \N__49795\,
            in3 => \N__49625\,
            lcout => n20585,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_4_lut_adj_241_LC_18_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011111110"
        )
    port map (
            in0 => \N__49627\,
            in1 => \N__49774\,
            in2 => \N__49144\,
            in3 => \N__53438\,
            lcout => n11824,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_valid_85_LC_18_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46381\,
            in2 => \_gnd_net_\,
            in3 => \N__46342\,
            lcout => comm_data_vld,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcomm_spi.data_valid_85C_net\,
            ce => 'H',
            sr => \N__55383\
        );

    \i18843_2_lut_3_lut_LC_18_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__49628\,
            in1 => \N__49770\,
            in2 => \_gnd_net_\,
            in3 => \N__53900\,
            lcout => n21087,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_1__bdd_4_lut_19462_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011001100"
        )
    port map (
            in0 => \N__46753\,
            in1 => \N__49396\,
            in2 => \N__46717\,
            in3 => \N__50006\,
            lcout => OPEN,
            ltout => \n22063_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i4_LC_18_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010010100100"
        )
    port map (
            in0 => \N__50007\,
            in1 => \N__46597\,
            in2 => \N__46741\,
            in3 => \N__46537\,
            lcout => comm_tx_buf_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55143\,
            ce => \N__47104\,
            sr => \N__47048\
        );

    \i19042_2_lut_LC_18_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51516\,
            in2 => \_gnd_net_\,
            in3 => \N__46738\,
            lcout => n21081,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_137_Mux_4_i1_3_lut_LC_18_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__51518\,
            in1 => \N__46707\,
            in2 => \_gnd_net_\,
            in3 => \N__46664\,
            lcout => n1_adj_1564,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_181_LC_18_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__49781\,
            in1 => \N__49298\,
            in2 => \_gnd_net_\,
            in3 => \N__49624\,
            lcout => n18824,
            ltout => \n18824_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_LC_18_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51515\,
            in2 => \N__46591\,
            in3 => \N__49395\,
            lcout => n20507,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_137_Mux_4_i2_3_lut_LC_18_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__51517\,
            in1 => \_gnd_net_\,
            in2 => \N__46567\,
            in3 => \N__46552\,
            lcout => n2_adj_1565,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_137_Mux_1_i4_3_lut_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__46531\,
            in1 => \N__46522\,
            in2 => \_gnd_net_\,
            in3 => \N__51605\,
            lcout => OPEN,
            ltout => \n4_adj_1569_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18197_4_lut_LC_18_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__51606\,
            in1 => \N__49467\,
            in2 => \N__47179\,
            in3 => \N__47176\,
            lcout => OPEN,
            ltout => \n20792_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_tx_buf_i1_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__50010\,
            in1 => \_gnd_net_\,
            in2 => \N__47158\,
            in3 => \N__47155\,
            lcout => comm_tx_buf_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55157\,
            ce => \N__47135\,
            sr => \N__47052\
        );

    \i19037_3_lut_4_lut_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__51604\,
            in1 => \N__50009\,
            in2 => \N__49514\,
            in3 => \N__49939\,
            lcout => n21069,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \data_cntvec_i0_i0_LC_18_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46928\,
            in2 => \N__46987\,
            in3 => \_gnd_net_\,
            lcout => data_cntvec_0,
            ltout => OPEN,
            carryin => \bfn_18_12_0_\,
            carryout => n19296,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__48662\,
            sr => \N__48604\
        );

    \data_cntvec_i0_i1_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46907\,
            in2 => \_gnd_net_\,
            in3 => \N__46885\,
            lcout => data_cntvec_1,
            ltout => OPEN,
            carryin => n19296,
            carryout => n19297,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__48662\,
            sr => \N__48604\
        );

    \data_cntvec_i0_i2_LC_18_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46871\,
            in2 => \_gnd_net_\,
            in3 => \N__46855\,
            lcout => data_cntvec_2,
            ltout => OPEN,
            carryin => n19297,
            carryout => n19298,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__48662\,
            sr => \N__48604\
        );

    \data_cntvec_i0_i3_LC_18_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46838\,
            in2 => \_gnd_net_\,
            in3 => \N__46816\,
            lcout => data_cntvec_3,
            ltout => OPEN,
            carryin => n19298,
            carryout => n19299,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__48662\,
            sr => \N__48604\
        );

    \data_cntvec_i0_i4_LC_18_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46802\,
            in2 => \_gnd_net_\,
            in3 => \N__46786\,
            lcout => data_cntvec_4,
            ltout => OPEN,
            carryin => n19299,
            carryout => n19300,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__48662\,
            sr => \N__48604\
        );

    \data_cntvec_i0_i5_LC_18_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46772\,
            in2 => \_gnd_net_\,
            in3 => \N__46756\,
            lcout => data_cntvec_5,
            ltout => OPEN,
            carryin => n19300,
            carryout => n19301,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__48662\,
            sr => \N__48604\
        );

    \data_cntvec_i0_i6_LC_18_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47402\,
            in2 => \_gnd_net_\,
            in3 => \N__47380\,
            lcout => data_cntvec_6,
            ltout => OPEN,
            carryin => n19301,
            carryout => n19302,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__48662\,
            sr => \N__48604\
        );

    \data_cntvec_i0_i7_LC_18_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47369\,
            in2 => \_gnd_net_\,
            in3 => \N__47347\,
            lcout => data_cntvec_7,
            ltout => OPEN,
            carryin => n19302,
            carryout => n19303,
            clk => \INVdata_cntvec_i0_i0C_net\,
            ce => \N__48662\,
            sr => \N__48604\
        );

    \data_cntvec_i0_i8_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47336\,
            in2 => \_gnd_net_\,
            in3 => \N__47314\,
            lcout => data_cntvec_8,
            ltout => OPEN,
            carryin => \bfn_18_13_0_\,
            carryout => n19304,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__48667\,
            sr => \N__48603\
        );

    \data_cntvec_i0_i9_LC_18_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47297\,
            in2 => \_gnd_net_\,
            in3 => \N__47281\,
            lcout => data_cntvec_9,
            ltout => OPEN,
            carryin => n19304,
            carryout => n19305,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__48667\,
            sr => \N__48603\
        );

    \data_cntvec_i0_i10_LC_18_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47267\,
            in2 => \_gnd_net_\,
            in3 => \N__47245\,
            lcout => data_cntvec_10,
            ltout => OPEN,
            carryin => n19305,
            carryout => n19306,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__48667\,
            sr => \N__48603\
        );

    \data_cntvec_i0_i11_LC_18_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47242\,
            in2 => \_gnd_net_\,
            in3 => \N__47224\,
            lcout => data_cntvec_11,
            ltout => OPEN,
            carryin => n19306,
            carryout => n19307,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__48667\,
            sr => \N__48603\
        );

    \data_cntvec_i0_i12_LC_18_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47217\,
            in2 => \_gnd_net_\,
            in3 => \N__47203\,
            lcout => data_cntvec_12,
            ltout => OPEN,
            carryin => n19307,
            carryout => n19308,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__48667\,
            sr => \N__48603\
        );

    \data_cntvec_i0_i13_LC_18_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47196\,
            in2 => \_gnd_net_\,
            in3 => \N__47182\,
            lcout => data_cntvec_13,
            ltout => OPEN,
            carryin => n19308,
            carryout => n19309,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__48667\,
            sr => \N__48603\
        );

    \data_cntvec_i0_i14_LC_18_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48700\,
            in2 => \_gnd_net_\,
            in3 => \N__48688\,
            lcout => data_cntvec_14,
            ltout => OPEN,
            carryin => n19309,
            carryout => n19310,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__48667\,
            sr => \N__48603\
        );

    \data_cntvec_i0_i15_LC_18_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48681\,
            in2 => \_gnd_net_\,
            in3 => \N__48685\,
            lcout => data_cntvec_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVdata_cntvec_i0_i8C_net\,
            ce => \N__48667\,
            sr => \N__48603\
        );

    \i6956_2_lut_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51221\,
            in2 => \_gnd_net_\,
            in3 => \N__53985\,
            lcout => n9273,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i6_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__49009\,
            in1 => \N__50964\,
            in2 => \N__48799\,
            in3 => \N__48557\,
            lcout => buf_adcdata_iac_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55201\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_VAC.ADC_DATA_i4_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__48534\,
            in1 => \N__48348\,
            in2 => \N__47968\,
            in3 => \N__51330\,
            lcout => buf_adcdata_vac_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55201\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_7_i19_3_lut_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47924\,
            in1 => \N__47908\,
            in2 => \_gnd_net_\,
            in3 => \N__56988\,
            lcout => OPEN,
            ltout => \n19_adj_1589_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_7_i22_3_lut_LC_18_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47873\,
            in2 => \N__47854\,
            in3 => \N__47846\,
            lcout => OPEN,
            ltout => \n22_adj_1590_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_7_i30_3_lut_LC_18_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47443\,
            in2 => \N__47431\,
            in3 => \N__56316\,
            lcout => n30_adj_1591,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i5_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__49000\,
            in1 => \N__50911\,
            in2 => \N__50323\,
            in3 => \N__49070\,
            lcout => buf_adcdata_iac_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55213\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i12_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000011001100"
        )
    port map (
            in0 => \N__50912\,
            in1 => \N__50540\,
            in2 => \N__49048\,
            in3 => \N__50527\,
            lcout => cmd_rdadctmp_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.ADC_DATA_i4_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__49004\,
            in1 => \N__50913\,
            in2 => \N__50547\,
            in3 => \N__48821\,
            lcout => buf_adcdata_iac_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.dds_state_i2_LC_18_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__55613\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55795\,
            lcout => dds_state_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55224\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i14_LC_18_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__48785\,
            in1 => \N__50914\,
            in2 => \N__50322\,
            in3 => \N__50526\,
            lcout => cmd_rdadctmp_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55233\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.iclk_40_12179_12180_set_LC_19_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52952\,
            lcout => \comm_spi.n14581\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55091\,
            ce => 'H',
            sr => \N__48760\
        );

    \comm_spi.RESET_I_0_90_2_lut_LC_19_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__52953\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55405\,
            lcout => \comm_spi.iclk_N_754\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_94_2_lut_LC_19_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48748\,
            in2 => \_gnd_net_\,
            in3 => \N__55406\,
            lcout => \comm_spi.data_tx_7__N_760\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i0_12175_12176_set_LC_19_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__52795\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \comm_spi.n14577\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52375\,
            ce => 'H',
            sr => \N__52897\
        );

    \comm_response_302_LC_19_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000100110"
        )
    port map (
            in0 => \N__53742\,
            in1 => \N__54244\,
            in2 => \N__51264\,
            in3 => \N__53450\,
            lcout => \ICE_GPMI_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55122\,
            ce => \N__49249\,
            sr => \_gnd_net_\
        );

    \i1_3_lut_4_lut_adj_258_LC_19_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001110100010"
        )
    port map (
            in0 => \N__53449\,
            in1 => \N__51234\,
            in2 => \N__54368\,
            in3 => \N__49186\,
            lcout => n11406,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i17_4_lut_3_lut_LC_19_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010110100000"
        )
    port map (
            in0 => \N__53741\,
            in1 => \_gnd_net_\,
            in2 => \N__51263\,
            in3 => \N__53448\,
            lcout => OPEN,
            ltout => \n10_adj_1572_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_285_LC_19_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011001000"
        )
    port map (
            in0 => \N__54240\,
            in1 => \N__49185\,
            in2 => \N__49147\,
            in3 => \_gnd_net_\,
            lcout => n11836,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_292_LC_19_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111111"
        )
    port map (
            in0 => \N__54239\,
            in1 => \N__51230\,
            in2 => \_gnd_net_\,
            in3 => \N__53740\,
            lcout => n20643,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_3_lut_adj_286_LC_19_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101111111111"
        )
    port map (
            in0 => \N__49699\,
            in1 => \N__53437\,
            in2 => \_gnd_net_\,
            in3 => \N__49635\,
            lcout => n4_adj_1596,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_index_i1_LC_19_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101111100100000"
        )
    port map (
            in0 => \N__49640\,
            in1 => \N__49769\,
            in2 => \N__51577\,
            in3 => \N__49462\,
            lcout => comm_index_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55144\,
            ce => \N__49102\,
            sr => \N__49093\
        );

    \comm_index_i0_LC_19_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100111001100"
        )
    port map (
            in0 => \N__49768\,
            in1 => \N__51533\,
            in2 => \_gnd_net_\,
            in3 => \N__49639\,
            lcout => comm_index_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55144\,
            ce => \N__49102\,
            sr => \N__49093\
        );

    \comm_index_i2_LC_19_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110110011001100"
        )
    port map (
            in0 => \N__51537\,
            in1 => \N__50008\,
            in2 => \N__49513\,
            in3 => \N__49120\,
            lcout => comm_index_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55144\,
            ce => \N__49102\,
            sr => \N__49093\
        );

    \comm_spi.i19169_4_lut_3_lut_LC_19_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__53193\,
            in1 => \N__50205\,
            in2 => \_gnd_net_\,
            in3 => \N__55382\,
            lcout => \comm_spi.n22647\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15191_2_lut_3_lut_LC_19_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__51225\,
            in1 => \N__50194\,
            in2 => \_gnd_net_\,
            in3 => \N__53884\,
            lcout => n14_adj_1557,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_adj_297_LC_19_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__50002\,
            in1 => \N__53361\,
            in2 => \N__49429\,
            in3 => \N__49940\,
            lcout => n20563,
            ltout => \n20563_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19_4_lut_adj_295_LC_19_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001110011"
        )
    port map (
            in0 => \N__51529\,
            in1 => \N__53883\,
            in2 => \N__49918\,
            in3 => \N__51684\,
            lcout => OPEN,
            ltout => \n12_adj_1539_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_3_lut_adj_296_LC_19_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49915\,
            in2 => \N__49873\,
            in3 => \N__49846\,
            lcout => n12164,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_4_lut_4_lut_LC_19_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011000000000"
        )
    port map (
            in0 => \N__51226\,
            in1 => \N__53885\,
            in2 => \N__49797\,
            in3 => \N__49634\,
            lcout => OPEN,
            ltout => \n21_adj_1573_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19127_4_lut_LC_19_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111100110111"
        )
    port map (
            in0 => \N__49573\,
            in1 => \N__56362\,
            in2 => \N__49558\,
            in3 => \N__51227\,
            lcout => n18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_adj_318_LC_19_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101100110"
        )
    port map (
            in0 => \N__49463\,
            in1 => \N__49344\,
            in2 => \_gnd_net_\,
            in3 => \N__49323\,
            lcout => OPEN,
            ltout => \n5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i19063_3_lut_LC_19_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000000000"
        )
    port map (
            in0 => \N__49303\,
            in1 => \_gnd_net_\,
            in2 => \N__49270\,
            in3 => \N__53882\,
            lcout => OPEN,
            ltout => \n21658_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18270_4_lut_LC_19_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010101010"
        )
    port map (
            in0 => \N__52246\,
            in1 => \N__52234\,
            in2 => \N__52198\,
            in3 => \N__51229\,
            lcout => OPEN,
            ltout => \n20865_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_state_i0_LC_19_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51881\,
            in2 => \N__51703\,
            in3 => \N__54536\,
            lcout => comm_state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55173\,
            ce => \N__51700\,
            sr => \_gnd_net_\
        );

    \i19_4_lut_adj_298_LC_19_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000100010001"
        )
    port map (
            in0 => \N__53881\,
            in1 => \N__51677\,
            in2 => \N__51619\,
            in3 => \N__51460\,
            lcout => n12_adj_1585,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15206_2_lut_3_lut_LC_19_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__51228\,
            in1 => \N__51442\,
            in2 => \_gnd_net_\,
            in3 => \N__53984\,
            lcout => n14_adj_1526,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_4_i19_3_lut_LC_19_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__51358\,
            in1 => \N__51326\,
            in2 => \_gnd_net_\,
            in3 => \N__56941\,
            lcout => n19_adj_1605,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18139_2_lut_3_lut_LC_19_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__51262\,
            in1 => \N__53983\,
            in2 => \_gnd_net_\,
            in3 => \N__53417\,
            lcout => n20734,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ADC_IAC.cmd_rdadctmp_i13_LC_19_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__50315\,
            in1 => \N__50915\,
            in2 => \N__50548\,
            in3 => \N__50517\,
            lcout => cmd_rdadctmp_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55234\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14972_2_lut_2_lut_LC_19_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__50292\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50266\,
            lcout => \CONT_SD\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.i23_4_lut_LC_19_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010011101"
        )
    port map (
            in0 => \N__55832\,
            in1 => \N__55738\,
            in2 => \N__53026\,
            in3 => \N__55585\,
            lcout => \SIG_DDS.n9_adj_1385\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.iclk_40_12179_12180_reset_LC_20_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52941\,
            lcout => \comm_spi.n14582\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55102\,
            ce => 'H',
            sr => \N__52906\
        );

    \comm_spi.RESET_I_0_91_2_lut_LC_20_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__52942\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55407\,
            lcout => \comm_spi.iclk_N_755\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_2_lut_LC_20_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__55377\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53258\,
            lcout => \comm_spi.data_tx_7__N_787\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_99_2_lut_LC_20_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__55378\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53259\,
            lcout => \comm_spi.data_tx_7__N_765\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.data_tx_i0_12175_12176_reset_LC_20_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__52724\,
            lcout => \comm_spi.n14578\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52437\,
            ce => 'H',
            sr => \N__52534\
        );

    \comm_spi.data_tx_i1_12201_12202_reset_LC_20_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__53233\,
            in1 => \N__52482\,
            in2 => \_gnd_net_\,
            in3 => \N__52497\,
            lcout => \comm_spi.n14604\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52415\,
            ce => 'H',
            sr => \N__53176\
        );

    \comm_spi.data_tx_i1_12201_12202_set_LC_20_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__53229\,
            in1 => \N__52501\,
            in2 => \_gnd_net_\,
            in3 => \N__52486\,
            lcout => \comm_spi.n14603\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__52444\,
            ce => 'H',
            sr => \N__53212\
        );

    \comm_spi.i19204_4_lut_3_lut_LC_20_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__53260\,
            in1 => \N__53228\,
            in2 => \_gnd_net_\,
            in3 => \N__55404\,
            lcout => \comm_spi.n22650\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_98_2_lut_LC_20_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__53200\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55403\,
            lcout => \comm_spi.data_tx_7__N_764\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_106_2_lut_LC_20_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__55402\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__53199\,
            lcout => \comm_spi.data_tx_7__N_784\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \comm_spi.RESET_I_0_103_2_lut_LC_20_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__53148\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__55401\,
            lcout => \comm_spi.data_tx_7__N_775\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6_4_lut_adj_231_LC_20_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__57715\,
            in1 => \N__57568\,
            in2 => \N__57673\,
            in3 => \N__53116\,
            lcout => n20502,
            ltout => \n20502_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15112_2_lut_LC_20_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__53119\,
            in3 => \N__57588\,
            lcout => n10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5_4_lut_adj_224_LC_20_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__57652\,
            in1 => \N__57616\,
            in2 => \N__57697\,
            in3 => \N__57634\,
            lcout => n12_adj_1583,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclk_294_LC_20_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101001100110"
        )
    port map (
            in0 => \N__55977\,
            in1 => \N__57589\,
            in2 => \_gnd_net_\,
            in3 => \N__53110\,
            lcout => dds0_mclk,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVdds0_mclk_294C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6_4_lut_adj_226_LC_20_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__53104\,
            in1 => \N__53089\,
            in2 => \N__53074\,
            in3 => \N__53053\,
            lcout => n14_adj_1578,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18214_4_lut_LC_20_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__57553\,
            in1 => \N__56978\,
            in2 => \N__56416\,
            in3 => \N__56401\,
            lcout => n20809,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15033_2_lut_LC_20_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54535\,
            in2 => \_gnd_net_\,
            in3 => \N__53371\,
            lcout => n17415,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mux_130_Mux_4_i30_3_lut_LC_20_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__56353\,
            in1 => \N__56310\,
            in2 => \_gnd_net_\,
            in3 => \N__56065\,
            lcout => n30_adj_1608,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \clk_16MHz_I_0_3_lut_LC_20_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__56041\,
            in1 => \N__55981\,
            in2 => \_gnd_net_\,
            in3 => \N__55966\,
            lcout => \DDS_MCLK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.SCLK_27_LC_20_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001010110001"
        )
    port map (
            in0 => \N__55744\,
            in1 => \N__55860\,
            in2 => \N__55905\,
            in3 => \N__55627\,
            lcout => \DDS_SCK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55241\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SIG_DDS.CS_28_LC_20_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000110111011"
        )
    port map (
            in0 => \N__55861\,
            in1 => \N__55740\,
            in2 => \_gnd_net_\,
            in3 => \N__55626\,
            lcout => \DDS_CS\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55244\,
            ce => \N__55483\,
            sr => \_gnd_net_\
        );

    \comm_clear_301_LC_22_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0111011100110011"
        )
    port map (
            in0 => \N__54561\,
            in1 => \N__54035\,
            in2 => \_gnd_net_\,
            in3 => \N__53486\,
            lcout => comm_clear,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__55187\,
            ce => \N__53266\,
            sr => \_gnd_net_\
        );

    \i2_2_lut_3_lut_adj_220_LC_22_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__54544\,
            in1 => \N__54034\,
            in2 => \_gnd_net_\,
            in3 => \N__53485\,
            lcout => n11347,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3772__i0_LC_22_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57714\,
            in2 => \_gnd_net_\,
            in3 => \N__57700\,
            lcout => dds0_mclkcnt_0,
            ltout => OPEN,
            carryin => \bfn_22_11_0_\,
            carryout => n19440,
            clk => \INVdds0_mclkcnt_i7_3772__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3772__i1_LC_22_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57693\,
            in2 => \_gnd_net_\,
            in3 => \N__57676\,
            lcout => dds0_mclkcnt_1,
            ltout => OPEN,
            carryin => n19440,
            carryout => n19441,
            clk => \INVdds0_mclkcnt_i7_3772__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3772__i2_LC_22_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57669\,
            in2 => \_gnd_net_\,
            in3 => \N__57655\,
            lcout => dds0_mclkcnt_2,
            ltout => OPEN,
            carryin => n19441,
            carryout => n19442,
            clk => \INVdds0_mclkcnt_i7_3772__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3772__i3_LC_22_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57651\,
            in2 => \_gnd_net_\,
            in3 => \N__57637\,
            lcout => dds0_mclkcnt_3,
            ltout => OPEN,
            carryin => n19442,
            carryout => n19443,
            clk => \INVdds0_mclkcnt_i7_3772__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3772__i4_LC_22_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57633\,
            in2 => \_gnd_net_\,
            in3 => \N__57619\,
            lcout => dds0_mclkcnt_4,
            ltout => OPEN,
            carryin => n19443,
            carryout => n19444,
            clk => \INVdds0_mclkcnt_i7_3772__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3772__i5_LC_22_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57615\,
            in2 => \_gnd_net_\,
            in3 => \N__57601\,
            lcout => dds0_mclkcnt_5,
            ltout => OPEN,
            carryin => n19444,
            carryout => n19445,
            clk => \INVdds0_mclkcnt_i7_3772__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3772__i6_LC_22_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57598\,
            in2 => \_gnd_net_\,
            in3 => \N__57574\,
            lcout => dds0_mclkcnt_6,
            ltout => OPEN,
            carryin => n19445,
            carryout => n19446,
            clk => \INVdds0_mclkcnt_i7_3772__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \dds0_mclkcnt_i7_3772__i7_LC_22_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57567\,
            in2 => \_gnd_net_\,
            in3 => \N__57571\,
            lcout => dds0_mclkcnt_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVdds0_mclkcnt_i7_3772__i0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
