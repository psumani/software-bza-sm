// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jan 27 2023 14:59:49

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "zim" view "INTERFACE"

module zim (
    VAC_DRDY,
    IAC_FLT1,
    DDS_SCK,
    ICE_IOR_166,
    ICE_IOR_119,
    DDS_MOSI,
    VAC_MISO,
    DDS_MOSI1,
    ICE_IOR_146,
    VDC_CLK,
    ICE_IOT_222,
    IAC_CS,
    ICE_IOL_18B,
    ICE_IOL_13A,
    ICE_IOB_81,
    VAC_OSR1,
    IAC_MOSI,
    DDS_CS1,
    ICE_IOL_4B,
    ICE_IOB_94,
    VAC_CS,
    VAC_CLK,
    ICE_SPI_CE0,
    ICE_IOR_167,
    ICE_IOR_118,
    RTD_SDO,
    IAC_OSR0,
    VDC_SCLK,
    VAC_FLT1,
    ICE_SPI_MOSI,
    ICE_IOR_165,
    ICE_IOR_147,
    ICE_IOL_14A,
    ICE_IOL_13B,
    ICE_IOB_91,
    ICE_GPMO_0,
    DDS_RNG_0,
    VDC_RNG0,
    ICE_SPI_SCLK,
    ICE_IOR_152,
    ICE_IOL_12A,
    RTD_DRDY,
    ICE_SPI_MISO,
    ICE_IOT_177,
    ICE_IOR_141,
    ICE_IOB_80,
    ICE_IOB_102,
    ICE_GPMO_2,
    ICE_GPMI_0,
    IAC_MISO,
    VAC_OSR0,
    VAC_MOSI,
    TEST_LED,
    ICE_IOR_148,
    STAT_COMM,
    ICE_SYSCLK,
    ICE_IOR_161,
    ICE_IOB_95,
    ICE_IOB_82,
    ICE_IOB_104,
    IAC_CLK,
    DDS_CS,
    SELIRNG0,
    RTD_SDI,
    ICE_IOT_221,
    ICE_IOT_197,
    DDS_MCLK,
    RTD_SCLK,
    RTD_CS,
    ICE_IOR_137,
    IAC_OSR1,
    VAC_FLT0,
    ICE_IOR_144,
    ICE_IOR_128,
    ICE_GPMO_1,
    IAC_SCLK,
    EIS_SYNCCLK,
    ICE_IOR_139,
    ICE_IOL_4A,
    VAC_SCLK,
    THERMOSTAT,
    ICE_IOR_164,
    ICE_IOB_103,
    AMPV_POW,
    VDC_SDO,
    ICE_IOT_174,
    ICE_IOR_140,
    ICE_IOB_96,
    CONT_SD,
    AC_ADC_SYNC,
    SELIRNG1,
    ICE_IOL_12B,
    ICE_IOR_160,
    ICE_IOR_136,
    DDS_MCLK1,
    ICE_IOT_198,
    ICE_IOT_173,
    IAC_DRDY,
    ICE_IOT_178,
    ICE_IOR_138,
    ICE_IOR_120,
    IAC_FLT0,
    DDS_SCK1);

    input VAC_DRDY;
    output IAC_FLT1;
    output DDS_SCK;
    input ICE_IOR_166;
    input ICE_IOR_119;
    output DDS_MOSI;
    input VAC_MISO;
    output DDS_MOSI1;
    input ICE_IOR_146;
    output VDC_CLK;
    input ICE_IOT_222;
    output IAC_CS;
    input ICE_IOL_18B;
    input ICE_IOL_13A;
    input ICE_IOB_81;
    output VAC_OSR1;
    output IAC_MOSI;
    output DDS_CS1;
    input ICE_IOL_4B;
    input ICE_IOB_94;
    output VAC_CS;
    output VAC_CLK;
    input ICE_SPI_CE0;
    input ICE_IOR_167;
    input ICE_IOR_118;
    input RTD_SDO;
    output IAC_OSR0;
    output VDC_SCLK;
    output VAC_FLT1;
    input ICE_SPI_MOSI;
    input ICE_IOR_165;
    input ICE_IOR_147;
    input ICE_IOL_14A;
    input ICE_IOL_13B;
    input ICE_IOB_91;
    input ICE_GPMO_0;
    output DDS_RNG_0;
    output VDC_RNG0;
    input ICE_SPI_SCLK;
    input ICE_IOR_152;
    input ICE_IOL_12A;
    input RTD_DRDY;
    output ICE_SPI_MISO;
    input ICE_IOT_177;
    input ICE_IOR_141;
    input ICE_IOB_80;
    input ICE_IOB_102;
    input ICE_GPMO_2;
    output ICE_GPMI_0;
    input IAC_MISO;
    output VAC_OSR0;
    output VAC_MOSI;
    output TEST_LED;
    input ICE_IOR_148;
    output STAT_COMM;
    input ICE_SYSCLK;
    input ICE_IOR_161;
    input ICE_IOB_95;
    input ICE_IOB_82;
    input ICE_IOB_104;
    output IAC_CLK;
    output DDS_CS;
    output SELIRNG0;
    output RTD_SDI;
    input ICE_IOT_221;
    input ICE_IOT_197;
    output DDS_MCLK;
    output RTD_SCLK;
    output RTD_CS;
    input ICE_IOR_137;
    output IAC_OSR1;
    output VAC_FLT0;
    input ICE_IOR_144;
    input ICE_IOR_128;
    input ICE_GPMO_1;
    output IAC_SCLK;
    input EIS_SYNCCLK;
    input ICE_IOR_139;
    input ICE_IOL_4A;
    output VAC_SCLK;
    input THERMOSTAT;
    input ICE_IOR_164;
    input ICE_IOB_103;
    output AMPV_POW;
    input VDC_SDO;
    input ICE_IOT_174;
    input ICE_IOR_140;
    input ICE_IOB_96;
    output CONT_SD;
    output AC_ADC_SYNC;
    output SELIRNG1;
    input ICE_IOL_12B;
    input ICE_IOR_160;
    input ICE_IOR_136;
    output DDS_MCLK1;
    input ICE_IOT_198;
    input ICE_IOT_173;
    input IAC_DRDY;
    input ICE_IOT_178;
    input ICE_IOR_138;
    input ICE_IOR_120;
    output IAC_FLT0;
    output DDS_SCK1;

    wire N__58652;
    wire N__58651;
    wire N__58650;
    wire N__58643;
    wire N__58642;
    wire N__58641;
    wire N__58634;
    wire N__58633;
    wire N__58632;
    wire N__58625;
    wire N__58624;
    wire N__58623;
    wire N__58616;
    wire N__58615;
    wire N__58614;
    wire N__58607;
    wire N__58606;
    wire N__58605;
    wire N__58598;
    wire N__58597;
    wire N__58596;
    wire N__58589;
    wire N__58588;
    wire N__58587;
    wire N__58580;
    wire N__58579;
    wire N__58578;
    wire N__58571;
    wire N__58570;
    wire N__58569;
    wire N__58562;
    wire N__58561;
    wire N__58560;
    wire N__58553;
    wire N__58552;
    wire N__58551;
    wire N__58544;
    wire N__58543;
    wire N__58542;
    wire N__58535;
    wire N__58534;
    wire N__58533;
    wire N__58526;
    wire N__58525;
    wire N__58524;
    wire N__58517;
    wire N__58516;
    wire N__58515;
    wire N__58508;
    wire N__58507;
    wire N__58506;
    wire N__58499;
    wire N__58498;
    wire N__58497;
    wire N__58490;
    wire N__58489;
    wire N__58488;
    wire N__58481;
    wire N__58480;
    wire N__58479;
    wire N__58472;
    wire N__58471;
    wire N__58470;
    wire N__58463;
    wire N__58462;
    wire N__58461;
    wire N__58454;
    wire N__58453;
    wire N__58452;
    wire N__58445;
    wire N__58444;
    wire N__58443;
    wire N__58436;
    wire N__58435;
    wire N__58434;
    wire N__58427;
    wire N__58426;
    wire N__58425;
    wire N__58418;
    wire N__58417;
    wire N__58416;
    wire N__58409;
    wire N__58408;
    wire N__58407;
    wire N__58400;
    wire N__58399;
    wire N__58398;
    wire N__58391;
    wire N__58390;
    wire N__58389;
    wire N__58382;
    wire N__58381;
    wire N__58380;
    wire N__58373;
    wire N__58372;
    wire N__58371;
    wire N__58364;
    wire N__58363;
    wire N__58362;
    wire N__58355;
    wire N__58354;
    wire N__58353;
    wire N__58346;
    wire N__58345;
    wire N__58344;
    wire N__58337;
    wire N__58336;
    wire N__58335;
    wire N__58328;
    wire N__58327;
    wire N__58326;
    wire N__58319;
    wire N__58318;
    wire N__58317;
    wire N__58310;
    wire N__58309;
    wire N__58308;
    wire N__58301;
    wire N__58300;
    wire N__58299;
    wire N__58292;
    wire N__58291;
    wire N__58290;
    wire N__58283;
    wire N__58282;
    wire N__58281;
    wire N__58274;
    wire N__58273;
    wire N__58272;
    wire N__58265;
    wire N__58264;
    wire N__58263;
    wire N__58256;
    wire N__58255;
    wire N__58254;
    wire N__58247;
    wire N__58246;
    wire N__58245;
    wire N__58238;
    wire N__58237;
    wire N__58236;
    wire N__58229;
    wire N__58228;
    wire N__58227;
    wire N__58220;
    wire N__58219;
    wire N__58218;
    wire N__58211;
    wire N__58210;
    wire N__58209;
    wire N__58202;
    wire N__58201;
    wire N__58200;
    wire N__58193;
    wire N__58192;
    wire N__58191;
    wire N__58184;
    wire N__58183;
    wire N__58182;
    wire N__58175;
    wire N__58174;
    wire N__58173;
    wire N__58166;
    wire N__58165;
    wire N__58164;
    wire N__58157;
    wire N__58156;
    wire N__58155;
    wire N__58148;
    wire N__58147;
    wire N__58146;
    wire N__58139;
    wire N__58138;
    wire N__58137;
    wire N__58130;
    wire N__58129;
    wire N__58128;
    wire N__58121;
    wire N__58120;
    wire N__58119;
    wire N__58112;
    wire N__58111;
    wire N__58110;
    wire N__58103;
    wire N__58102;
    wire N__58101;
    wire N__58094;
    wire N__58093;
    wire N__58092;
    wire N__58085;
    wire N__58084;
    wire N__58083;
    wire N__58076;
    wire N__58075;
    wire N__58074;
    wire N__58067;
    wire N__58066;
    wire N__58065;
    wire N__58058;
    wire N__58057;
    wire N__58056;
    wire N__58049;
    wire N__58048;
    wire N__58047;
    wire N__58040;
    wire N__58039;
    wire N__58038;
    wire N__58031;
    wire N__58030;
    wire N__58029;
    wire N__58022;
    wire N__58021;
    wire N__58020;
    wire N__58013;
    wire N__58012;
    wire N__58011;
    wire N__58004;
    wire N__58003;
    wire N__58002;
    wire N__57995;
    wire N__57994;
    wire N__57993;
    wire N__57986;
    wire N__57985;
    wire N__57984;
    wire N__57977;
    wire N__57976;
    wire N__57975;
    wire N__57968;
    wire N__57967;
    wire N__57966;
    wire N__57959;
    wire N__57958;
    wire N__57957;
    wire N__57950;
    wire N__57949;
    wire N__57948;
    wire N__57941;
    wire N__57940;
    wire N__57939;
    wire N__57932;
    wire N__57931;
    wire N__57930;
    wire N__57923;
    wire N__57922;
    wire N__57921;
    wire N__57914;
    wire N__57913;
    wire N__57912;
    wire N__57905;
    wire N__57904;
    wire N__57903;
    wire N__57896;
    wire N__57895;
    wire N__57894;
    wire N__57887;
    wire N__57886;
    wire N__57885;
    wire N__57878;
    wire N__57877;
    wire N__57876;
    wire N__57869;
    wire N__57868;
    wire N__57867;
    wire N__57860;
    wire N__57859;
    wire N__57858;
    wire N__57851;
    wire N__57850;
    wire N__57849;
    wire N__57842;
    wire N__57841;
    wire N__57840;
    wire N__57833;
    wire N__57832;
    wire N__57831;
    wire N__57824;
    wire N__57823;
    wire N__57822;
    wire N__57815;
    wire N__57814;
    wire N__57813;
    wire N__57806;
    wire N__57805;
    wire N__57804;
    wire N__57797;
    wire N__57796;
    wire N__57795;
    wire N__57788;
    wire N__57787;
    wire N__57786;
    wire N__57779;
    wire N__57778;
    wire N__57777;
    wire N__57770;
    wire N__57769;
    wire N__57768;
    wire N__57761;
    wire N__57760;
    wire N__57759;
    wire N__57752;
    wire N__57751;
    wire N__57750;
    wire N__57743;
    wire N__57742;
    wire N__57741;
    wire N__57734;
    wire N__57733;
    wire N__57732;
    wire N__57715;
    wire N__57714;
    wire N__57711;
    wire N__57708;
    wire N__57705;
    wire N__57700;
    wire N__57697;
    wire N__57694;
    wire N__57693;
    wire N__57690;
    wire N__57687;
    wire N__57684;
    wire N__57679;
    wire N__57676;
    wire N__57673;
    wire N__57670;
    wire N__57669;
    wire N__57666;
    wire N__57663;
    wire N__57660;
    wire N__57655;
    wire N__57652;
    wire N__57651;
    wire N__57648;
    wire N__57645;
    wire N__57642;
    wire N__57637;
    wire N__57634;
    wire N__57633;
    wire N__57630;
    wire N__57627;
    wire N__57624;
    wire N__57619;
    wire N__57616;
    wire N__57615;
    wire N__57612;
    wire N__57609;
    wire N__57606;
    wire N__57601;
    wire N__57598;
    wire N__57595;
    wire N__57592;
    wire N__57589;
    wire N__57588;
    wire N__57583;
    wire N__57580;
    wire N__57577;
    wire N__57574;
    wire N__57571;
    wire N__57568;
    wire N__57567;
    wire N__57564;
    wire N__57561;
    wire N__57558;
    wire N__57553;
    wire N__57552;
    wire N__57551;
    wire N__57550;
    wire N__57549;
    wire N__57548;
    wire N__57547;
    wire N__57544;
    wire N__57543;
    wire N__57542;
    wire N__57541;
    wire N__57540;
    wire N__57539;
    wire N__57538;
    wire N__57537;
    wire N__57536;
    wire N__57535;
    wire N__57534;
    wire N__57533;
    wire N__57532;
    wire N__57531;
    wire N__57526;
    wire N__57525;
    wire N__57524;
    wire N__57523;
    wire N__57522;
    wire N__57521;
    wire N__57516;
    wire N__57513;
    wire N__57510;
    wire N__57507;
    wire N__57504;
    wire N__57503;
    wire N__57502;
    wire N__57497;
    wire N__57494;
    wire N__57493;
    wire N__57490;
    wire N__57489;
    wire N__57486;
    wire N__57485;
    wire N__57484;
    wire N__57483;
    wire N__57482;
    wire N__57481;
    wire N__57480;
    wire N__57479;
    wire N__57472;
    wire N__57469;
    wire N__57466;
    wire N__57465;
    wire N__57464;
    wire N__57463;
    wire N__57462;
    wire N__57459;
    wire N__57456;
    wire N__57453;
    wire N__57450;
    wire N__57449;
    wire N__57448;
    wire N__57447;
    wire N__57446;
    wire N__57445;
    wire N__57444;
    wire N__57443;
    wire N__57442;
    wire N__57441;
    wire N__57440;
    wire N__57437;
    wire N__57436;
    wire N__57433;
    wire N__57430;
    wire N__57427;
    wire N__57422;
    wire N__57419;
    wire N__57414;
    wire N__57411;
    wire N__57410;
    wire N__57409;
    wire N__57408;
    wire N__57407;
    wire N__57404;
    wire N__57399;
    wire N__57396;
    wire N__57395;
    wire N__57394;
    wire N__57393;
    wire N__57392;
    wire N__57391;
    wire N__57390;
    wire N__57389;
    wire N__57388;
    wire N__57387;
    wire N__57386;
    wire N__57383;
    wire N__57380;
    wire N__57377;
    wire N__57374;
    wire N__57371;
    wire N__57370;
    wire N__57367;
    wire N__57364;
    wire N__57359;
    wire N__57356;
    wire N__57353;
    wire N__57350;
    wire N__57347;
    wire N__57346;
    wire N__57345;
    wire N__57342;
    wire N__57341;
    wire N__57334;
    wire N__57331;
    wire N__57328;
    wire N__57323;
    wire N__57318;
    wire N__57315;
    wire N__57312;
    wire N__57311;
    wire N__57310;
    wire N__57305;
    wire N__57300;
    wire N__57297;
    wire N__57294;
    wire N__57291;
    wire N__57288;
    wire N__57279;
    wire N__57274;
    wire N__57271;
    wire N__57262;
    wire N__57259;
    wire N__57254;
    wire N__57251;
    wire N__57250;
    wire N__57243;
    wire N__57242;
    wire N__57241;
    wire N__57238;
    wire N__57233;
    wire N__57230;
    wire N__57225;
    wire N__57220;
    wire N__57215;
    wire N__57212;
    wire N__57209;
    wire N__57206;
    wire N__57193;
    wire N__57192;
    wire N__57191;
    wire N__57190;
    wire N__57189;
    wire N__57188;
    wire N__57187;
    wire N__57186;
    wire N__57185;
    wire N__57184;
    wire N__57183;
    wire N__57182;
    wire N__57181;
    wire N__57172;
    wire N__57163;
    wire N__57160;
    wire N__57157;
    wire N__57154;
    wire N__57149;
    wire N__57142;
    wire N__57135;
    wire N__57126;
    wire N__57119;
    wire N__57116;
    wire N__57113;
    wire N__57108;
    wire N__57091;
    wire N__57086;
    wire N__57081;
    wire N__57074;
    wire N__57071;
    wire N__57064;
    wire N__57061;
    wire N__57058;
    wire N__57055;
    wire N__57050;
    wire N__57045;
    wire N__57040;
    wire N__57037;
    wire N__57032;
    wire N__57029;
    wire N__57018;
    wire N__56989;
    wire N__56988;
    wire N__56985;
    wire N__56984;
    wire N__56983;
    wire N__56982;
    wire N__56979;
    wire N__56978;
    wire N__56977;
    wire N__56974;
    wire N__56969;
    wire N__56968;
    wire N__56967;
    wire N__56966;
    wire N__56965;
    wire N__56964;
    wire N__56961;
    wire N__56960;
    wire N__56959;
    wire N__56958;
    wire N__56957;
    wire N__56956;
    wire N__56955;
    wire N__56954;
    wire N__56953;
    wire N__56952;
    wire N__56951;
    wire N__56950;
    wire N__56949;
    wire N__56946;
    wire N__56945;
    wire N__56942;
    wire N__56941;
    wire N__56940;
    wire N__56939;
    wire N__56938;
    wire N__56935;
    wire N__56934;
    wire N__56933;
    wire N__56932;
    wire N__56931;
    wire N__56930;
    wire N__56929;
    wire N__56928;
    wire N__56927;
    wire N__56922;
    wire N__56921;
    wire N__56918;
    wire N__56915;
    wire N__56914;
    wire N__56913;
    wire N__56912;
    wire N__56911;
    wire N__56910;
    wire N__56909;
    wire N__56908;
    wire N__56907;
    wire N__56906;
    wire N__56905;
    wire N__56904;
    wire N__56903;
    wire N__56902;
    wire N__56901;
    wire N__56898;
    wire N__56897;
    wire N__56894;
    wire N__56891;
    wire N__56890;
    wire N__56889;
    wire N__56888;
    wire N__56887;
    wire N__56886;
    wire N__56885;
    wire N__56884;
    wire N__56883;
    wire N__56880;
    wire N__56875;
    wire N__56868;
    wire N__56867;
    wire N__56866;
    wire N__56865;
    wire N__56860;
    wire N__56855;
    wire N__56848;
    wire N__56845;
    wire N__56842;
    wire N__56841;
    wire N__56840;
    wire N__56837;
    wire N__56834;
    wire N__56833;
    wire N__56832;
    wire N__56831;
    wire N__56824;
    wire N__56811;
    wire N__56804;
    wire N__56803;
    wire N__56802;
    wire N__56801;
    wire N__56800;
    wire N__56799;
    wire N__56798;
    wire N__56797;
    wire N__56794;
    wire N__56791;
    wire N__56786;
    wire N__56781;
    wire N__56778;
    wire N__56775;
    wire N__56772;
    wire N__56763;
    wire N__56760;
    wire N__56757;
    wire N__56754;
    wire N__56749;
    wire N__56746;
    wire N__56743;
    wire N__56738;
    wire N__56733;
    wire N__56730;
    wire N__56727;
    wire N__56726;
    wire N__56725;
    wire N__56722;
    wire N__56717;
    wire N__56714;
    wire N__56707;
    wire N__56700;
    wire N__56699;
    wire N__56698;
    wire N__56695;
    wire N__56694;
    wire N__56693;
    wire N__56690;
    wire N__56687;
    wire N__56686;
    wire N__56685;
    wire N__56684;
    wire N__56683;
    wire N__56678;
    wire N__56675;
    wire N__56672;
    wire N__56667;
    wire N__56662;
    wire N__56659;
    wire N__56652;
    wire N__56649;
    wire N__56646;
    wire N__56643;
    wire N__56642;
    wire N__56641;
    wire N__56640;
    wire N__56639;
    wire N__56638;
    wire N__56637;
    wire N__56636;
    wire N__56635;
    wire N__56634;
    wire N__56625;
    wire N__56616;
    wire N__56607;
    wire N__56598;
    wire N__56595;
    wire N__56584;
    wire N__56579;
    wire N__56568;
    wire N__56567;
    wire N__56564;
    wire N__56563;
    wire N__56562;
    wire N__56559;
    wire N__56556;
    wire N__56551;
    wire N__56546;
    wire N__56543;
    wire N__56536;
    wire N__56533;
    wire N__56528;
    wire N__56517;
    wire N__56512;
    wire N__56509;
    wire N__56502;
    wire N__56499;
    wire N__56490;
    wire N__56487;
    wire N__56480;
    wire N__56471;
    wire N__56462;
    wire N__56451;
    wire N__56446;
    wire N__56441;
    wire N__56416;
    wire N__56413;
    wire N__56410;
    wire N__56407;
    wire N__56404;
    wire N__56401;
    wire N__56398;
    wire N__56397;
    wire N__56394;
    wire N__56391;
    wire N__56388;
    wire N__56387;
    wire N__56382;
    wire N__56379;
    wire N__56374;
    wire N__56371;
    wire N__56368;
    wire N__56365;
    wire N__56362;
    wire N__56359;
    wire N__56356;
    wire N__56353;
    wire N__56350;
    wire N__56347;
    wire N__56346;
    wire N__56345;
    wire N__56344;
    wire N__56343;
    wire N__56342;
    wire N__56341;
    wire N__56340;
    wire N__56339;
    wire N__56338;
    wire N__56337;
    wire N__56336;
    wire N__56335;
    wire N__56334;
    wire N__56331;
    wire N__56326;
    wire N__56321;
    wire N__56318;
    wire N__56317;
    wire N__56316;
    wire N__56315;
    wire N__56312;
    wire N__56311;
    wire N__56310;
    wire N__56309;
    wire N__56308;
    wire N__56301;
    wire N__56296;
    wire N__56291;
    wire N__56290;
    wire N__56289;
    wire N__56288;
    wire N__56287;
    wire N__56284;
    wire N__56281;
    wire N__56278;
    wire N__56275;
    wire N__56274;
    wire N__56273;
    wire N__56272;
    wire N__56271;
    wire N__56270;
    wire N__56269;
    wire N__56266;
    wire N__56265;
    wire N__56264;
    wire N__56261;
    wire N__56260;
    wire N__56259;
    wire N__56258;
    wire N__56257;
    wire N__56256;
    wire N__56253;
    wire N__56248;
    wire N__56245;
    wire N__56240;
    wire N__56233;
    wire N__56228;
    wire N__56225;
    wire N__56222;
    wire N__56213;
    wire N__56210;
    wire N__56207;
    wire N__56204;
    wire N__56201;
    wire N__56198;
    wire N__56195;
    wire N__56192;
    wire N__56187;
    wire N__56184;
    wire N__56181;
    wire N__56176;
    wire N__56173;
    wire N__56170;
    wire N__56169;
    wire N__56166;
    wire N__56161;
    wire N__56156;
    wire N__56147;
    wire N__56146;
    wire N__56145;
    wire N__56144;
    wire N__56139;
    wire N__56134;
    wire N__56131;
    wire N__56118;
    wire N__56115;
    wire N__56112;
    wire N__56109;
    wire N__56106;
    wire N__56103;
    wire N__56098;
    wire N__56091;
    wire N__56082;
    wire N__56065;
    wire N__56062;
    wire N__56059;
    wire N__56056;
    wire N__56053;
    wire N__56050;
    wire N__56047;
    wire N__56044;
    wire N__56041;
    wire N__56040;
    wire N__56037;
    wire N__56034;
    wire N__56031;
    wire N__56030;
    wire N__56029;
    wire N__56028;
    wire N__56027;
    wire N__56026;
    wire N__56025;
    wire N__56024;
    wire N__56023;
    wire N__56022;
    wire N__56019;
    wire N__56018;
    wire N__56017;
    wire N__56016;
    wire N__56015;
    wire N__55984;
    wire N__55981;
    wire N__55978;
    wire N__55977;
    wire N__55974;
    wire N__55971;
    wire N__55966;
    wire N__55963;
    wire N__55962;
    wire N__55959;
    wire N__55956;
    wire N__55953;
    wire N__55950;
    wire N__55949;
    wire N__55944;
    wire N__55941;
    wire N__55938;
    wire N__55933;
    wire N__55930;
    wire N__55927;
    wire N__55924;
    wire N__55921;
    wire N__55918;
    wire N__55915;
    wire N__55912;
    wire N__55909;
    wire N__55906;
    wire N__55905;
    wire N__55902;
    wire N__55899;
    wire N__55896;
    wire N__55893;
    wire N__55888;
    wire N__55887;
    wire N__55886;
    wire N__55885;
    wire N__55884;
    wire N__55883;
    wire N__55882;
    wire N__55881;
    wire N__55880;
    wire N__55879;
    wire N__55878;
    wire N__55875;
    wire N__55874;
    wire N__55873;
    wire N__55872;
    wire N__55871;
    wire N__55870;
    wire N__55869;
    wire N__55868;
    wire N__55867;
    wire N__55866;
    wire N__55863;
    wire N__55862;
    wire N__55861;
    wire N__55860;
    wire N__55845;
    wire N__55840;
    wire N__55833;
    wire N__55832;
    wire N__55827;
    wire N__55816;
    wire N__55813;
    wire N__55810;
    wire N__55807;
    wire N__55804;
    wire N__55801;
    wire N__55796;
    wire N__55795;
    wire N__55792;
    wire N__55787;
    wire N__55784;
    wire N__55781;
    wire N__55776;
    wire N__55771;
    wire N__55768;
    wire N__55765;
    wire N__55760;
    wire N__55753;
    wire N__55744;
    wire N__55741;
    wire N__55740;
    wire N__55739;
    wire N__55738;
    wire N__55737;
    wire N__55734;
    wire N__55731;
    wire N__55728;
    wire N__55725;
    wire N__55722;
    wire N__55713;
    wire N__55712;
    wire N__55711;
    wire N__55708;
    wire N__55705;
    wire N__55700;
    wire N__55697;
    wire N__55696;
    wire N__55695;
    wire N__55690;
    wire N__55687;
    wire N__55682;
    wire N__55679;
    wire N__55672;
    wire N__55669;
    wire N__55668;
    wire N__55667;
    wire N__55666;
    wire N__55665;
    wire N__55664;
    wire N__55663;
    wire N__55662;
    wire N__55661;
    wire N__55660;
    wire N__55659;
    wire N__55656;
    wire N__55655;
    wire N__55640;
    wire N__55635;
    wire N__55634;
    wire N__55633;
    wire N__55632;
    wire N__55631;
    wire N__55630;
    wire N__55629;
    wire N__55628;
    wire N__55627;
    wire N__55626;
    wire N__55623;
    wire N__55622;
    wire N__55621;
    wire N__55620;
    wire N__55617;
    wire N__55614;
    wire N__55613;
    wire N__55608;
    wire N__55603;
    wire N__55592;
    wire N__55589;
    wire N__55586;
    wire N__55585;
    wire N__55582;
    wire N__55579;
    wire N__55574;
    wire N__55571;
    wire N__55568;
    wire N__55567;
    wire N__55566;
    wire N__55563;
    wire N__55556;
    wire N__55553;
    wire N__55550;
    wire N__55547;
    wire N__55540;
    wire N__55537;
    wire N__55534;
    wire N__55529;
    wire N__55524;
    wire N__55515;
    wire N__55504;
    wire N__55501;
    wire N__55498;
    wire N__55495;
    wire N__55492;
    wire N__55489;
    wire N__55486;
    wire N__55483;
    wire N__55480;
    wire N__55477;
    wire N__55474;
    wire N__55473;
    wire N__55472;
    wire N__55469;
    wire N__55466;
    wire N__55465;
    wire N__55464;
    wire N__55463;
    wire N__55462;
    wire N__55461;
    wire N__55460;
    wire N__55459;
    wire N__55458;
    wire N__55455;
    wire N__55452;
    wire N__55443;
    wire N__55438;
    wire N__55437;
    wire N__55432;
    wire N__55431;
    wire N__55430;
    wire N__55429;
    wire N__55428;
    wire N__55427;
    wire N__55426;
    wire N__55425;
    wire N__55424;
    wire N__55423;
    wire N__55422;
    wire N__55421;
    wire N__55418;
    wire N__55415;
    wire N__55410;
    wire N__55409;
    wire N__55408;
    wire N__55407;
    wire N__55406;
    wire N__55405;
    wire N__55404;
    wire N__55403;
    wire N__55402;
    wire N__55401;
    wire N__55398;
    wire N__55395;
    wire N__55392;
    wire N__55389;
    wire N__55384;
    wire N__55383;
    wire N__55382;
    wire N__55379;
    wire N__55378;
    wire N__55377;
    wire N__55362;
    wire N__55355;
    wire N__55350;
    wire N__55347;
    wire N__55342;
    wire N__55333;
    wire N__55328;
    wire N__55321;
    wire N__55318;
    wire N__55315;
    wire N__55312;
    wire N__55307;
    wire N__55304;
    wire N__55299;
    wire N__55294;
    wire N__55291;
    wire N__55284;
    wire N__55281;
    wire N__55274;
    wire N__55271;
    wire N__55268;
    wire N__55263;
    wire N__55258;
    wire N__55255;
    wire N__55246;
    wire N__55245;
    wire N__55244;
    wire N__55243;
    wire N__55242;
    wire N__55241;
    wire N__55240;
    wire N__55239;
    wire N__55238;
    wire N__55237;
    wire N__55236;
    wire N__55235;
    wire N__55234;
    wire N__55233;
    wire N__55232;
    wire N__55231;
    wire N__55230;
    wire N__55229;
    wire N__55228;
    wire N__55227;
    wire N__55226;
    wire N__55225;
    wire N__55224;
    wire N__55223;
    wire N__55222;
    wire N__55221;
    wire N__55220;
    wire N__55219;
    wire N__55218;
    wire N__55217;
    wire N__55216;
    wire N__55215;
    wire N__55214;
    wire N__55213;
    wire N__55212;
    wire N__55211;
    wire N__55210;
    wire N__55209;
    wire N__55208;
    wire N__55207;
    wire N__55206;
    wire N__55205;
    wire N__55204;
    wire N__55203;
    wire N__55202;
    wire N__55201;
    wire N__55200;
    wire N__55199;
    wire N__55198;
    wire N__55197;
    wire N__55196;
    wire N__55195;
    wire N__55194;
    wire N__55193;
    wire N__55192;
    wire N__55191;
    wire N__55190;
    wire N__55189;
    wire N__55188;
    wire N__55187;
    wire N__55186;
    wire N__55185;
    wire N__55184;
    wire N__55183;
    wire N__55182;
    wire N__55181;
    wire N__55180;
    wire N__55179;
    wire N__55178;
    wire N__55177;
    wire N__55176;
    wire N__55175;
    wire N__55174;
    wire N__55173;
    wire N__55172;
    wire N__55171;
    wire N__55170;
    wire N__55169;
    wire N__55168;
    wire N__55167;
    wire N__55166;
    wire N__55165;
    wire N__55164;
    wire N__55163;
    wire N__55162;
    wire N__55161;
    wire N__55160;
    wire N__55159;
    wire N__55158;
    wire N__55157;
    wire N__55156;
    wire N__55155;
    wire N__55154;
    wire N__55153;
    wire N__55152;
    wire N__55151;
    wire N__55150;
    wire N__55149;
    wire N__55148;
    wire N__55147;
    wire N__55146;
    wire N__55145;
    wire N__55144;
    wire N__55143;
    wire N__55142;
    wire N__55141;
    wire N__55140;
    wire N__55139;
    wire N__55138;
    wire N__55137;
    wire N__55136;
    wire N__55135;
    wire N__55134;
    wire N__55133;
    wire N__55132;
    wire N__55131;
    wire N__55130;
    wire N__55129;
    wire N__55128;
    wire N__55127;
    wire N__55126;
    wire N__55125;
    wire N__55124;
    wire N__55123;
    wire N__55122;
    wire N__55121;
    wire N__55120;
    wire N__55119;
    wire N__55118;
    wire N__55117;
    wire N__55116;
    wire N__55115;
    wire N__55114;
    wire N__55113;
    wire N__55112;
    wire N__55111;
    wire N__55110;
    wire N__55109;
    wire N__55108;
    wire N__55107;
    wire N__55106;
    wire N__55105;
    wire N__55104;
    wire N__55103;
    wire N__55102;
    wire N__55101;
    wire N__55100;
    wire N__55099;
    wire N__55098;
    wire N__55097;
    wire N__55096;
    wire N__55095;
    wire N__55094;
    wire N__55093;
    wire N__55092;
    wire N__55091;
    wire N__55090;
    wire N__55089;
    wire N__55088;
    wire N__55087;
    wire N__55086;
    wire N__55085;
    wire N__55084;
    wire N__55083;
    wire N__55082;
    wire N__55081;
    wire N__55080;
    wire N__55079;
    wire N__55078;
    wire N__55077;
    wire N__55076;
    wire N__55075;
    wire N__55074;
    wire N__54727;
    wire N__54724;
    wire N__54723;
    wire N__54722;
    wire N__54721;
    wire N__54720;
    wire N__54719;
    wire N__54718;
    wire N__54717;
    wire N__54716;
    wire N__54715;
    wire N__54714;
    wire N__54713;
    wire N__54712;
    wire N__54711;
    wire N__54710;
    wire N__54709;
    wire N__54706;
    wire N__54705;
    wire N__54704;
    wire N__54703;
    wire N__54702;
    wire N__54701;
    wire N__54700;
    wire N__54699;
    wire N__54696;
    wire N__54695;
    wire N__54694;
    wire N__54693;
    wire N__54690;
    wire N__54687;
    wire N__54684;
    wire N__54681;
    wire N__54676;
    wire N__54675;
    wire N__54674;
    wire N__54673;
    wire N__54672;
    wire N__54671;
    wire N__54670;
    wire N__54669;
    wire N__54668;
    wire N__54667;
    wire N__54666;
    wire N__54665;
    wire N__54664;
    wire N__54663;
    wire N__54662;
    wire N__54661;
    wire N__54660;
    wire N__54659;
    wire N__54658;
    wire N__54657;
    wire N__54656;
    wire N__54653;
    wire N__54650;
    wire N__54649;
    wire N__54646;
    wire N__54645;
    wire N__54642;
    wire N__54639;
    wire N__54636;
    wire N__54635;
    wire N__54632;
    wire N__54629;
    wire N__54626;
    wire N__54625;
    wire N__54624;
    wire N__54623;
    wire N__54620;
    wire N__54617;
    wire N__54612;
    wire N__54611;
    wire N__54610;
    wire N__54609;
    wire N__54604;
    wire N__54601;
    wire N__54600;
    wire N__54599;
    wire N__54598;
    wire N__54597;
    wire N__54596;
    wire N__54593;
    wire N__54592;
    wire N__54591;
    wire N__54590;
    wire N__54589;
    wire N__54588;
    wire N__54585;
    wire N__54584;
    wire N__54581;
    wire N__54580;
    wire N__54577;
    wire N__54576;
    wire N__54571;
    wire N__54564;
    wire N__54563;
    wire N__54562;
    wire N__54561;
    wire N__54558;
    wire N__54555;
    wire N__54550;
    wire N__54545;
    wire N__54544;
    wire N__54541;
    wire N__54538;
    wire N__54537;
    wire N__54536;
    wire N__54535;
    wire N__54522;
    wire N__54511;
    wire N__54508;
    wire N__54495;
    wire N__54490;
    wire N__54489;
    wire N__54488;
    wire N__54487;
    wire N__54486;
    wire N__54485;
    wire N__54482;
    wire N__54475;
    wire N__54472;
    wire N__54467;
    wire N__54460;
    wire N__54455;
    wire N__54452;
    wire N__54451;
    wire N__54448;
    wire N__54445;
    wire N__54442;
    wire N__54441;
    wire N__54440;
    wire N__54437;
    wire N__54434;
    wire N__54433;
    wire N__54430;
    wire N__54427;
    wire N__54424;
    wire N__54421;
    wire N__54416;
    wire N__54399;
    wire N__54394;
    wire N__54389;
    wire N__54388;
    wire N__54387;
    wire N__54384;
    wire N__54381;
    wire N__54376;
    wire N__54373;
    wire N__54372;
    wire N__54369;
    wire N__54368;
    wire N__54367;
    wire N__54364;
    wire N__54361;
    wire N__54358;
    wire N__54355;
    wire N__54352;
    wire N__54341;
    wire N__54336;
    wire N__54329;
    wire N__54318;
    wire N__54315;
    wire N__54312;
    wire N__54309;
    wire N__54306;
    wire N__54301;
    wire N__54298;
    wire N__54295;
    wire N__54288;
    wire N__54285;
    wire N__54280;
    wire N__54275;
    wire N__54268;
    wire N__54263;
    wire N__54260;
    wire N__54253;
    wire N__54250;
    wire N__54249;
    wire N__54246;
    wire N__54245;
    wire N__54244;
    wire N__54241;
    wire N__54240;
    wire N__54239;
    wire N__54238;
    wire N__54235;
    wire N__54228;
    wire N__54223;
    wire N__54220;
    wire N__54211;
    wire N__54200;
    wire N__54193;
    wire N__54184;
    wire N__54177;
    wire N__54176;
    wire N__54175;
    wire N__54172;
    wire N__54169;
    wire N__54166;
    wire N__54157;
    wire N__54154;
    wire N__54143;
    wire N__54138;
    wire N__54135;
    wire N__54132;
    wire N__54127;
    wire N__54106;
    wire N__54105;
    wire N__54104;
    wire N__54103;
    wire N__54102;
    wire N__54101;
    wire N__54100;
    wire N__54099;
    wire N__54098;
    wire N__54097;
    wire N__54096;
    wire N__54095;
    wire N__54094;
    wire N__54093;
    wire N__54092;
    wire N__54091;
    wire N__54090;
    wire N__54089;
    wire N__54088;
    wire N__54087;
    wire N__54086;
    wire N__54085;
    wire N__54084;
    wire N__54083;
    wire N__54082;
    wire N__54081;
    wire N__54080;
    wire N__54079;
    wire N__54076;
    wire N__54067;
    wire N__54064;
    wire N__54061;
    wire N__54052;
    wire N__54051;
    wire N__54048;
    wire N__54045;
    wire N__54042;
    wire N__54039;
    wire N__54036;
    wire N__54035;
    wire N__54034;
    wire N__54033;
    wire N__54032;
    wire N__54031;
    wire N__54028;
    wire N__54027;
    wire N__54010;
    wire N__54005;
    wire N__54002;
    wire N__54001;
    wire N__54000;
    wire N__53997;
    wire N__53988;
    wire N__53987;
    wire N__53986;
    wire N__53985;
    wire N__53984;
    wire N__53983;
    wire N__53982;
    wire N__53981;
    wire N__53980;
    wire N__53979;
    wire N__53978;
    wire N__53977;
    wire N__53976;
    wire N__53975;
    wire N__53972;
    wire N__53967;
    wire N__53964;
    wire N__53961;
    wire N__53958;
    wire N__53957;
    wire N__53956;
    wire N__53953;
    wire N__53950;
    wire N__53949;
    wire N__53948;
    wire N__53947;
    wire N__53946;
    wire N__53945;
    wire N__53944;
    wire N__53943;
    wire N__53942;
    wire N__53941;
    wire N__53940;
    wire N__53939;
    wire N__53938;
    wire N__53937;
    wire N__53936;
    wire N__53935;
    wire N__53932;
    wire N__53929;
    wire N__53926;
    wire N__53923;
    wire N__53920;
    wire N__53913;
    wire N__53910;
    wire N__53909;
    wire N__53908;
    wire N__53905;
    wire N__53904;
    wire N__53903;
    wire N__53902;
    wire N__53901;
    wire N__53900;
    wire N__53895;
    wire N__53892;
    wire N__53889;
    wire N__53886;
    wire N__53885;
    wire N__53884;
    wire N__53883;
    wire N__53882;
    wire N__53881;
    wire N__53878;
    wire N__53875;
    wire N__53874;
    wire N__53873;
    wire N__53872;
    wire N__53871;
    wire N__53854;
    wire N__53851;
    wire N__53848;
    wire N__53843;
    wire N__53840;
    wire N__53839;
    wire N__53838;
    wire N__53837;
    wire N__53834;
    wire N__53831;
    wire N__53830;
    wire N__53829;
    wire N__53828;
    wire N__53823;
    wire N__53806;
    wire N__53791;
    wire N__53780;
    wire N__53777;
    wire N__53774;
    wire N__53771;
    wire N__53768;
    wire N__53765;
    wire N__53756;
    wire N__53753;
    wire N__53750;
    wire N__53743;
    wire N__53742;
    wire N__53741;
    wire N__53740;
    wire N__53733;
    wire N__53728;
    wire N__53723;
    wire N__53720;
    wire N__53713;
    wire N__53704;
    wire N__53701;
    wire N__53696;
    wire N__53693;
    wire N__53688;
    wire N__53687;
    wire N__53686;
    wire N__53685;
    wire N__53682;
    wire N__53681;
    wire N__53680;
    wire N__53679;
    wire N__53676;
    wire N__53673;
    wire N__53670;
    wire N__53659;
    wire N__53658;
    wire N__53657;
    wire N__53656;
    wire N__53655;
    wire N__53654;
    wire N__53645;
    wire N__53638;
    wire N__53637;
    wire N__53630;
    wire N__53623;
    wire N__53608;
    wire N__53601;
    wire N__53592;
    wire N__53587;
    wire N__53582;
    wire N__53571;
    wire N__53568;
    wire N__53565;
    wire N__53562;
    wire N__53555;
    wire N__53536;
    wire N__53533;
    wire N__53532;
    wire N__53531;
    wire N__53530;
    wire N__53529;
    wire N__53526;
    wire N__53523;
    wire N__53522;
    wire N__53521;
    wire N__53518;
    wire N__53513;
    wire N__53512;
    wire N__53511;
    wire N__53510;
    wire N__53509;
    wire N__53506;
    wire N__53503;
    wire N__53500;
    wire N__53499;
    wire N__53498;
    wire N__53497;
    wire N__53496;
    wire N__53495;
    wire N__53494;
    wire N__53493;
    wire N__53492;
    wire N__53491;
    wire N__53490;
    wire N__53489;
    wire N__53488;
    wire N__53487;
    wire N__53486;
    wire N__53485;
    wire N__53482;
    wire N__53479;
    wire N__53476;
    wire N__53475;
    wire N__53474;
    wire N__53467;
    wire N__53466;
    wire N__53463;
    wire N__53462;
    wire N__53461;
    wire N__53454;
    wire N__53451;
    wire N__53450;
    wire N__53449;
    wire N__53448;
    wire N__53439;
    wire N__53438;
    wire N__53437;
    wire N__53432;
    wire N__53421;
    wire N__53418;
    wire N__53417;
    wire N__53414;
    wire N__53411;
    wire N__53408;
    wire N__53403;
    wire N__53398;
    wire N__53395;
    wire N__53392;
    wire N__53389;
    wire N__53384;
    wire N__53379;
    wire N__53372;
    wire N__53371;
    wire N__53368;
    wire N__53365;
    wire N__53362;
    wire N__53361;
    wire N__53358;
    wire N__53353;
    wire N__53350;
    wire N__53345;
    wire N__53340;
    wire N__53337;
    wire N__53332;
    wire N__53327;
    wire N__53324;
    wire N__53321;
    wire N__53318;
    wire N__53311;
    wire N__53308;
    wire N__53303;
    wire N__53300;
    wire N__53291;
    wire N__53288;
    wire N__53285;
    wire N__53266;
    wire N__53263;
    wire N__53260;
    wire N__53259;
    wire N__53258;
    wire N__53255;
    wire N__53250;
    wire N__53247;
    wire N__53244;
    wire N__53239;
    wire N__53236;
    wire N__53233;
    wire N__53230;
    wire N__53229;
    wire N__53228;
    wire N__53225;
    wire N__53222;
    wire N__53219;
    wire N__53212;
    wire N__53209;
    wire N__53206;
    wire N__53203;
    wire N__53200;
    wire N__53199;
    wire N__53194;
    wire N__53193;
    wire N__53190;
    wire N__53187;
    wire N__53184;
    wire N__53181;
    wire N__53176;
    wire N__53173;
    wire N__53170;
    wire N__53167;
    wire N__53164;
    wire N__53161;
    wire N__53160;
    wire N__53157;
    wire N__53154;
    wire N__53149;
    wire N__53148;
    wire N__53145;
    wire N__53142;
    wire N__53139;
    wire N__53136;
    wire N__53131;
    wire N__53128;
    wire N__53125;
    wire N__53122;
    wire N__53119;
    wire N__53116;
    wire N__53113;
    wire N__53110;
    wire N__53107;
    wire N__53104;
    wire N__53103;
    wire N__53100;
    wire N__53097;
    wire N__53094;
    wire N__53089;
    wire N__53088;
    wire N__53085;
    wire N__53082;
    wire N__53079;
    wire N__53074;
    wire N__53071;
    wire N__53068;
    wire N__53067;
    wire N__53064;
    wire N__53061;
    wire N__53058;
    wire N__53053;
    wire N__53052;
    wire N__53049;
    wire N__53046;
    wire N__53043;
    wire N__53038;
    wire N__53035;
    wire N__53032;
    wire N__53029;
    wire N__53026;
    wire N__53025;
    wire N__53022;
    wire N__53019;
    wire N__53018;
    wire N__53015;
    wire N__53012;
    wire N__53009;
    wire N__53006;
    wire N__53005;
    wire N__53002;
    wire N__52999;
    wire N__52996;
    wire N__52993;
    wire N__52990;
    wire N__52985;
    wire N__52982;
    wire N__52979;
    wire N__52976;
    wire N__52969;
    wire N__52966;
    wire N__52963;
    wire N__52960;
    wire N__52957;
    wire N__52954;
    wire N__52953;
    wire N__52952;
    wire N__52949;
    wire N__52946;
    wire N__52943;
    wire N__52942;
    wire N__52941;
    wire N__52938;
    wire N__52933;
    wire N__52930;
    wire N__52927;
    wire N__52924;
    wire N__52917;
    wire N__52914;
    wire N__52911;
    wire N__52906;
    wire N__52903;
    wire N__52900;
    wire N__52897;
    wire N__52894;
    wire N__52891;
    wire N__52888;
    wire N__52887;
    wire N__52886;
    wire N__52883;
    wire N__52880;
    wire N__52879;
    wire N__52878;
    wire N__52877;
    wire N__52874;
    wire N__52873;
    wire N__52868;
    wire N__52865;
    wire N__52862;
    wire N__52861;
    wire N__52860;
    wire N__52857;
    wire N__52854;
    wire N__52851;
    wire N__52844;
    wire N__52841;
    wire N__52838;
    wire N__52837;
    wire N__52836;
    wire N__52835;
    wire N__52832;
    wire N__52831;
    wire N__52830;
    wire N__52829;
    wire N__52828;
    wire N__52823;
    wire N__52816;
    wire N__52813;
    wire N__52812;
    wire N__52811;
    wire N__52810;
    wire N__52809;
    wire N__52806;
    wire N__52805;
    wire N__52804;
    wire N__52803;
    wire N__52802;
    wire N__52801;
    wire N__52800;
    wire N__52799;
    wire N__52796;
    wire N__52795;
    wire N__52794;
    wire N__52793;
    wire N__52792;
    wire N__52791;
    wire N__52788;
    wire N__52785;
    wire N__52784;
    wire N__52781;
    wire N__52780;
    wire N__52777;
    wire N__52776;
    wire N__52773;
    wire N__52766;
    wire N__52763;
    wire N__52762;
    wire N__52759;
    wire N__52758;
    wire N__52755;
    wire N__52754;
    wire N__52751;
    wire N__52750;
    wire N__52749;
    wire N__52748;
    wire N__52747;
    wire N__52744;
    wire N__52737;
    wire N__52728;
    wire N__52725;
    wire N__52724;
    wire N__52723;
    wire N__52720;
    wire N__52719;
    wire N__52716;
    wire N__52715;
    wire N__52712;
    wire N__52711;
    wire N__52708;
    wire N__52707;
    wire N__52704;
    wire N__52701;
    wire N__52686;
    wire N__52683;
    wire N__52668;
    wire N__52667;
    wire N__52664;
    wire N__52663;
    wire N__52660;
    wire N__52659;
    wire N__52656;
    wire N__52655;
    wire N__52652;
    wire N__52649;
    wire N__52644;
    wire N__52641;
    wire N__52638;
    wire N__52635;
    wire N__52632;
    wire N__52615;
    wire N__52610;
    wire N__52605;
    wire N__52588;
    wire N__52585;
    wire N__52582;
    wire N__52577;
    wire N__52574;
    wire N__52571;
    wire N__52568;
    wire N__52561;
    wire N__52556;
    wire N__52551;
    wire N__52546;
    wire N__52543;
    wire N__52534;
    wire N__52531;
    wire N__52528;
    wire N__52525;
    wire N__52522;
    wire N__52519;
    wire N__52518;
    wire N__52515;
    wire N__52512;
    wire N__52507;
    wire N__52504;
    wire N__52501;
    wire N__52498;
    wire N__52497;
    wire N__52494;
    wire N__52491;
    wire N__52486;
    wire N__52483;
    wire N__52482;
    wire N__52479;
    wire N__52476;
    wire N__52471;
    wire N__52468;
    wire N__52465;
    wire N__52462;
    wire N__52461;
    wire N__52458;
    wire N__52455;
    wire N__52452;
    wire N__52449;
    wire N__52444;
    wire N__52443;
    wire N__52442;
    wire N__52441;
    wire N__52438;
    wire N__52437;
    wire N__52434;
    wire N__52431;
    wire N__52430;
    wire N__52427;
    wire N__52426;
    wire N__52425;
    wire N__52424;
    wire N__52421;
    wire N__52418;
    wire N__52417;
    wire N__52416;
    wire N__52415;
    wire N__52414;
    wire N__52413;
    wire N__52408;
    wire N__52407;
    wire N__52404;
    wire N__52401;
    wire N__52398;
    wire N__52395;
    wire N__52392;
    wire N__52391;
    wire N__52386;
    wire N__52383;
    wire N__52380;
    wire N__52379;
    wire N__52376;
    wire N__52375;
    wire N__52372;
    wire N__52369;
    wire N__52368;
    wire N__52365;
    wire N__52364;
    wire N__52361;
    wire N__52360;
    wire N__52353;
    wire N__52348;
    wire N__52345;
    wire N__52340;
    wire N__52337;
    wire N__52334;
    wire N__52331;
    wire N__52328;
    wire N__52323;
    wire N__52320;
    wire N__52319;
    wire N__52316;
    wire N__52313;
    wire N__52310;
    wire N__52307;
    wire N__52304;
    wire N__52293;
    wire N__52288;
    wire N__52283;
    wire N__52280;
    wire N__52277;
    wire N__52274;
    wire N__52267;
    wire N__52264;
    wire N__52257;
    wire N__52246;
    wire N__52243;
    wire N__52240;
    wire N__52237;
    wire N__52234;
    wire N__52233;
    wire N__52232;
    wire N__52229;
    wire N__52226;
    wire N__52223;
    wire N__52220;
    wire N__52217;
    wire N__52214;
    wire N__52211;
    wire N__52208;
    wire N__52205;
    wire N__52198;
    wire N__52195;
    wire N__52194;
    wire N__52193;
    wire N__52192;
    wire N__52191;
    wire N__52190;
    wire N__52189;
    wire N__52186;
    wire N__52185;
    wire N__52182;
    wire N__52181;
    wire N__52178;
    wire N__52177;
    wire N__52176;
    wire N__52175;
    wire N__52174;
    wire N__52173;
    wire N__52172;
    wire N__52171;
    wire N__52170;
    wire N__52169;
    wire N__52168;
    wire N__52167;
    wire N__52166;
    wire N__52163;
    wire N__52162;
    wire N__52161;
    wire N__52160;
    wire N__52159;
    wire N__52158;
    wire N__52151;
    wire N__52148;
    wire N__52147;
    wire N__52140;
    wire N__52135;
    wire N__52132;
    wire N__52125;
    wire N__52124;
    wire N__52123;
    wire N__52120;
    wire N__52117;
    wire N__52114;
    wire N__52113;
    wire N__52112;
    wire N__52111;
    wire N__52110;
    wire N__52109;
    wire N__52108;
    wire N__52105;
    wire N__52102;
    wire N__52099;
    wire N__52096;
    wire N__52093;
    wire N__52092;
    wire N__52091;
    wire N__52088;
    wire N__52087;
    wire N__52084;
    wire N__52081;
    wire N__52078;
    wire N__52077;
    wire N__52074;
    wire N__52069;
    wire N__52066;
    wire N__52065;
    wire N__52064;
    wire N__52063;
    wire N__52062;
    wire N__52061;
    wire N__52060;
    wire N__52059;
    wire N__52050;
    wire N__52047;
    wire N__52044;
    wire N__52043;
    wire N__52042;
    wire N__52037;
    wire N__52034;
    wire N__52033;
    wire N__52030;
    wire N__52027;
    wire N__52024;
    wire N__52017;
    wire N__52012;
    wire N__52007;
    wire N__52004;
    wire N__52001;
    wire N__51998;
    wire N__51995;
    wire N__51986;
    wire N__51985;
    wire N__51984;
    wire N__51983;
    wire N__51980;
    wire N__51979;
    wire N__51978;
    wire N__51977;
    wire N__51976;
    wire N__51975;
    wire N__51974;
    wire N__51971;
    wire N__51968;
    wire N__51963;
    wire N__51958;
    wire N__51955;
    wire N__51952;
    wire N__51951;
    wire N__51950;
    wire N__51945;
    wire N__51942;
    wire N__51937;
    wire N__51934;
    wire N__51931;
    wire N__51930;
    wire N__51929;
    wire N__51924;
    wire N__51921;
    wire N__51920;
    wire N__51919;
    wire N__51916;
    wire N__51915;
    wire N__51914;
    wire N__51907;
    wire N__51900;
    wire N__51895;
    wire N__51894;
    wire N__51893;
    wire N__51888;
    wire N__51885;
    wire N__51882;
    wire N__51881;
    wire N__51878;
    wire N__51873;
    wire N__51870;
    wire N__51861;
    wire N__51852;
    wire N__51849;
    wire N__51842;
    wire N__51835;
    wire N__51826;
    wire N__51823;
    wire N__51818;
    wire N__51815;
    wire N__51812;
    wire N__51807;
    wire N__51800;
    wire N__51795;
    wire N__51792;
    wire N__51787;
    wire N__51786;
    wire N__51783;
    wire N__51782;
    wire N__51763;
    wire N__51758;
    wire N__51755;
    wire N__51752;
    wire N__51747;
    wire N__51740;
    wire N__51737;
    wire N__51734;
    wire N__51731;
    wire N__51728;
    wire N__51725;
    wire N__51716;
    wire N__51703;
    wire N__51700;
    wire N__51697;
    wire N__51694;
    wire N__51691;
    wire N__51688;
    wire N__51685;
    wire N__51684;
    wire N__51681;
    wire N__51678;
    wire N__51677;
    wire N__51674;
    wire N__51671;
    wire N__51668;
    wire N__51665;
    wire N__51660;
    wire N__51659;
    wire N__51656;
    wire N__51653;
    wire N__51650;
    wire N__51643;
    wire N__51642;
    wire N__51641;
    wire N__51640;
    wire N__51639;
    wire N__51638;
    wire N__51633;
    wire N__51632;
    wire N__51631;
    wire N__51630;
    wire N__51629;
    wire N__51628;
    wire N__51627;
    wire N__51626;
    wire N__51625;
    wire N__51624;
    wire N__51623;
    wire N__51622;
    wire N__51621;
    wire N__51620;
    wire N__51619;
    wire N__51610;
    wire N__51607;
    wire N__51606;
    wire N__51605;
    wire N__51604;
    wire N__51601;
    wire N__51592;
    wire N__51583;
    wire N__51580;
    wire N__51579;
    wire N__51578;
    wire N__51577;
    wire N__51570;
    wire N__51567;
    wire N__51564;
    wire N__51561;
    wire N__51554;
    wire N__51551;
    wire N__51544;
    wire N__51541;
    wire N__51538;
    wire N__51537;
    wire N__51534;
    wire N__51533;
    wire N__51530;
    wire N__51529;
    wire N__51526;
    wire N__51519;
    wire N__51518;
    wire N__51517;
    wire N__51516;
    wire N__51515;
    wire N__51510;
    wire N__51505;
    wire N__51498;
    wire N__51495;
    wire N__51492;
    wire N__51487;
    wire N__51478;
    wire N__51473;
    wire N__51460;
    wire N__51457;
    wire N__51454;
    wire N__51451;
    wire N__51448;
    wire N__51445;
    wire N__51442;
    wire N__51439;
    wire N__51438;
    wire N__51435;
    wire N__51432;
    wire N__51431;
    wire N__51430;
    wire N__51429;
    wire N__51428;
    wire N__51425;
    wire N__51420;
    wire N__51417;
    wire N__51414;
    wire N__51411;
    wire N__51406;
    wire N__51403;
    wire N__51400;
    wire N__51397;
    wire N__51394;
    wire N__51391;
    wire N__51386;
    wire N__51383;
    wire N__51376;
    wire N__51375;
    wire N__51372;
    wire N__51369;
    wire N__51364;
    wire N__51361;
    wire N__51358;
    wire N__51355;
    wire N__51352;
    wire N__51349;
    wire N__51346;
    wire N__51343;
    wire N__51342;
    wire N__51339;
    wire N__51336;
    wire N__51331;
    wire N__51330;
    wire N__51327;
    wire N__51326;
    wire N__51323;
    wire N__51320;
    wire N__51317;
    wire N__51310;
    wire N__51307;
    wire N__51304;
    wire N__51301;
    wire N__51298;
    wire N__51297;
    wire N__51294;
    wire N__51293;
    wire N__51290;
    wire N__51287;
    wire N__51286;
    wire N__51285;
    wire N__51284;
    wire N__51283;
    wire N__51282;
    wire N__51279;
    wire N__51276;
    wire N__51273;
    wire N__51268;
    wire N__51265;
    wire N__51264;
    wire N__51263;
    wire N__51262;
    wire N__51261;
    wire N__51260;
    wire N__51259;
    wire N__51254;
    wire N__51251;
    wire N__51244;
    wire N__51241;
    wire N__51240;
    wire N__51239;
    wire N__51238;
    wire N__51235;
    wire N__51234;
    wire N__51231;
    wire N__51230;
    wire N__51229;
    wire N__51228;
    wire N__51227;
    wire N__51226;
    wire N__51225;
    wire N__51222;
    wire N__51221;
    wire N__51220;
    wire N__51219;
    wire N__51218;
    wire N__51217;
    wire N__51214;
    wire N__51211;
    wire N__51210;
    wire N__51209;
    wire N__51208;
    wire N__51207;
    wire N__51206;
    wire N__51205;
    wire N__51204;
    wire N__51201;
    wire N__51200;
    wire N__51199;
    wire N__51198;
    wire N__51197;
    wire N__51196;
    wire N__51193;
    wire N__51186;
    wire N__51181;
    wire N__51178;
    wire N__51169;
    wire N__51166;
    wire N__51163;
    wire N__51156;
    wire N__51153;
    wire N__51150;
    wire N__51143;
    wire N__51134;
    wire N__51129;
    wire N__51126;
    wire N__51123;
    wire N__51118;
    wire N__51115;
    wire N__51112;
    wire N__51111;
    wire N__51110;
    wire N__51107;
    wire N__51106;
    wire N__51105;
    wire N__51104;
    wire N__51101;
    wire N__51096;
    wire N__51087;
    wire N__51084;
    wire N__51075;
    wire N__51074;
    wire N__51073;
    wire N__51070;
    wire N__51063;
    wire N__51062;
    wire N__51061;
    wire N__51058;
    wire N__51049;
    wire N__51044;
    wire N__51041;
    wire N__51038;
    wire N__51033;
    wire N__51022;
    wire N__51017;
    wire N__51014;
    wire N__51011;
    wire N__51006;
    wire N__51001;
    wire N__50980;
    wire N__50977;
    wire N__50974;
    wire N__50971;
    wire N__50968;
    wire N__50965;
    wire N__50964;
    wire N__50963;
    wire N__50962;
    wire N__50961;
    wire N__50960;
    wire N__50957;
    wire N__50956;
    wire N__50955;
    wire N__50954;
    wire N__50953;
    wire N__50952;
    wire N__50951;
    wire N__50950;
    wire N__50949;
    wire N__50948;
    wire N__50945;
    wire N__50938;
    wire N__50937;
    wire N__50936;
    wire N__50935;
    wire N__50934;
    wire N__50931;
    wire N__50922;
    wire N__50921;
    wire N__50920;
    wire N__50919;
    wire N__50916;
    wire N__50915;
    wire N__50914;
    wire N__50913;
    wire N__50912;
    wire N__50911;
    wire N__50910;
    wire N__50909;
    wire N__50908;
    wire N__50907;
    wire N__50906;
    wire N__50903;
    wire N__50896;
    wire N__50893;
    wire N__50888;
    wire N__50885;
    wire N__50884;
    wire N__50883;
    wire N__50882;
    wire N__50881;
    wire N__50880;
    wire N__50877;
    wire N__50872;
    wire N__50867;
    wire N__50860;
    wire N__50857;
    wire N__50856;
    wire N__50855;
    wire N__50852;
    wire N__50849;
    wire N__50844;
    wire N__50841;
    wire N__50838;
    wire N__50837;
    wire N__50836;
    wire N__50835;
    wire N__50834;
    wire N__50831;
    wire N__50830;
    wire N__50825;
    wire N__50822;
    wire N__50821;
    wire N__50818;
    wire N__50813;
    wire N__50810;
    wire N__50805;
    wire N__50802;
    wire N__50801;
    wire N__50798;
    wire N__50793;
    wire N__50788;
    wire N__50781;
    wire N__50776;
    wire N__50771;
    wire N__50766;
    wire N__50763;
    wire N__50760;
    wire N__50759;
    wire N__50756;
    wire N__50753;
    wire N__50750;
    wire N__50749;
    wire N__50748;
    wire N__50747;
    wire N__50746;
    wire N__50741;
    wire N__50736;
    wire N__50733;
    wire N__50730;
    wire N__50725;
    wire N__50724;
    wire N__50723;
    wire N__50718;
    wire N__50717;
    wire N__50716;
    wire N__50715;
    wire N__50714;
    wire N__50713;
    wire N__50712;
    wire N__50711;
    wire N__50710;
    wire N__50707;
    wire N__50704;
    wire N__50695;
    wire N__50692;
    wire N__50689;
    wire N__50686;
    wire N__50681;
    wire N__50666;
    wire N__50663;
    wire N__50660;
    wire N__50657;
    wire N__50652;
    wire N__50651;
    wire N__50650;
    wire N__50649;
    wire N__50648;
    wire N__50647;
    wire N__50646;
    wire N__50645;
    wire N__50642;
    wire N__50639;
    wire N__50636;
    wire N__50619;
    wire N__50614;
    wire N__50611;
    wire N__50606;
    wire N__50603;
    wire N__50594;
    wire N__50589;
    wire N__50582;
    wire N__50573;
    wire N__50548;
    wire N__50547;
    wire N__50544;
    wire N__50541;
    wire N__50540;
    wire N__50537;
    wire N__50532;
    wire N__50527;
    wire N__50526;
    wire N__50523;
    wire N__50520;
    wire N__50519;
    wire N__50518;
    wire N__50517;
    wire N__50516;
    wire N__50515;
    wire N__50514;
    wire N__50513;
    wire N__50512;
    wire N__50507;
    wire N__50502;
    wire N__50501;
    wire N__50500;
    wire N__50497;
    wire N__50496;
    wire N__50495;
    wire N__50494;
    wire N__50493;
    wire N__50492;
    wire N__50491;
    wire N__50486;
    wire N__50483;
    wire N__50480;
    wire N__50479;
    wire N__50476;
    wire N__50471;
    wire N__50470;
    wire N__50469;
    wire N__50466;
    wire N__50463;
    wire N__50460;
    wire N__50459;
    wire N__50458;
    wire N__50457;
    wire N__50456;
    wire N__50455;
    wire N__50454;
    wire N__50453;
    wire N__50448;
    wire N__50443;
    wire N__50438;
    wire N__50431;
    wire N__50428;
    wire N__50425;
    wire N__50422;
    wire N__50419;
    wire N__50418;
    wire N__50417;
    wire N__50416;
    wire N__50415;
    wire N__50412;
    wire N__50409;
    wire N__50406;
    wire N__50403;
    wire N__50390;
    wire N__50387;
    wire N__50378;
    wire N__50373;
    wire N__50370;
    wire N__50367;
    wire N__50358;
    wire N__50353;
    wire N__50350;
    wire N__50347;
    wire N__50336;
    wire N__50323;
    wire N__50322;
    wire N__50319;
    wire N__50316;
    wire N__50315;
    wire N__50312;
    wire N__50309;
    wire N__50306;
    wire N__50299;
    wire N__50296;
    wire N__50293;
    wire N__50292;
    wire N__50289;
    wire N__50286;
    wire N__50285;
    wire N__50282;
    wire N__50279;
    wire N__50276;
    wire N__50273;
    wire N__50266;
    wire N__50263;
    wire N__50260;
    wire N__50257;
    wire N__50256;
    wire N__50255;
    wire N__50252;
    wire N__50249;
    wire N__50246;
    wire N__50239;
    wire N__50236;
    wire N__50233;
    wire N__50230;
    wire N__50227;
    wire N__50224;
    wire N__50221;
    wire N__50220;
    wire N__50217;
    wire N__50214;
    wire N__50211;
    wire N__50206;
    wire N__50205;
    wire N__50202;
    wire N__50199;
    wire N__50194;
    wire N__50191;
    wire N__50190;
    wire N__50187;
    wire N__50184;
    wire N__50183;
    wire N__50182;
    wire N__50181;
    wire N__50178;
    wire N__50175;
    wire N__50172;
    wire N__50169;
    wire N__50166;
    wire N__50163;
    wire N__50158;
    wire N__50155;
    wire N__50148;
    wire N__50145;
    wire N__50142;
    wire N__50137;
    wire N__50136;
    wire N__50133;
    wire N__50132;
    wire N__50129;
    wire N__50126;
    wire N__50123;
    wire N__50120;
    wire N__50115;
    wire N__50110;
    wire N__50107;
    wire N__50104;
    wire N__50101;
    wire N__50100;
    wire N__50099;
    wire N__50098;
    wire N__50097;
    wire N__50096;
    wire N__50095;
    wire N__50094;
    wire N__50089;
    wire N__50088;
    wire N__50087;
    wire N__50082;
    wire N__50079;
    wire N__50078;
    wire N__50077;
    wire N__50076;
    wire N__50075;
    wire N__50070;
    wire N__50069;
    wire N__50068;
    wire N__50067;
    wire N__50064;
    wire N__50061;
    wire N__50058;
    wire N__50055;
    wire N__50050;
    wire N__50047;
    wire N__50040;
    wire N__50037;
    wire N__50030;
    wire N__50027;
    wire N__50016;
    wire N__50011;
    wire N__50010;
    wire N__50009;
    wire N__50008;
    wire N__50007;
    wire N__50006;
    wire N__50003;
    wire N__50002;
    wire N__49999;
    wire N__49994;
    wire N__49989;
    wire N__49986;
    wire N__49981;
    wire N__49978;
    wire N__49975;
    wire N__49968;
    wire N__49957;
    wire N__49954;
    wire N__49951;
    wire N__49948;
    wire N__49947;
    wire N__49944;
    wire N__49941;
    wire N__49940;
    wire N__49939;
    wire N__49936;
    wire N__49933;
    wire N__49930;
    wire N__49927;
    wire N__49918;
    wire N__49915;
    wire N__49914;
    wire N__49911;
    wire N__49910;
    wire N__49909;
    wire N__49908;
    wire N__49905;
    wire N__49902;
    wire N__49897;
    wire N__49894;
    wire N__49891;
    wire N__49888;
    wire N__49883;
    wire N__49876;
    wire N__49873;
    wire N__49870;
    wire N__49869;
    wire N__49864;
    wire N__49861;
    wire N__49860;
    wire N__49859;
    wire N__49858;
    wire N__49855;
    wire N__49850;
    wire N__49847;
    wire N__49846;
    wire N__49839;
    wire N__49836;
    wire N__49831;
    wire N__49828;
    wire N__49825;
    wire N__49822;
    wire N__49821;
    wire N__49818;
    wire N__49815;
    wire N__49812;
    wire N__49809;
    wire N__49804;
    wire N__49801;
    wire N__49800;
    wire N__49799;
    wire N__49798;
    wire N__49797;
    wire N__49796;
    wire N__49795;
    wire N__49792;
    wire N__49791;
    wire N__49790;
    wire N__49783;
    wire N__49782;
    wire N__49781;
    wire N__49778;
    wire N__49775;
    wire N__49774;
    wire N__49771;
    wire N__49770;
    wire N__49769;
    wire N__49768;
    wire N__49767;
    wire N__49764;
    wire N__49759;
    wire N__49756;
    wire N__49755;
    wire N__49752;
    wire N__49751;
    wire N__49750;
    wire N__49747;
    wire N__49744;
    wire N__49735;
    wire N__49730;
    wire N__49727;
    wire N__49722;
    wire N__49719;
    wire N__49712;
    wire N__49709;
    wire N__49700;
    wire N__49699;
    wire N__49696;
    wire N__49693;
    wire N__49690;
    wire N__49683;
    wire N__49680;
    wire N__49677;
    wire N__49674;
    wire N__49671;
    wire N__49666;
    wire N__49661;
    wire N__49656;
    wire N__49653;
    wire N__49650;
    wire N__49645;
    wire N__49642;
    wire N__49641;
    wire N__49640;
    wire N__49639;
    wire N__49636;
    wire N__49635;
    wire N__49634;
    wire N__49633;
    wire N__49632;
    wire N__49629;
    wire N__49628;
    wire N__49627;
    wire N__49626;
    wire N__49625;
    wire N__49624;
    wire N__49619;
    wire N__49616;
    wire N__49613;
    wire N__49610;
    wire N__49605;
    wire N__49602;
    wire N__49593;
    wire N__49590;
    wire N__49573;
    wire N__49570;
    wire N__49567;
    wire N__49564;
    wire N__49561;
    wire N__49558;
    wire N__49555;
    wire N__49552;
    wire N__49549;
    wire N__49546;
    wire N__49543;
    wire N__49540;
    wire N__49539;
    wire N__49538;
    wire N__49537;
    wire N__49536;
    wire N__49535;
    wire N__49534;
    wire N__49533;
    wire N__49532;
    wire N__49531;
    wire N__49530;
    wire N__49529;
    wire N__49526;
    wire N__49525;
    wire N__49524;
    wire N__49523;
    wire N__49522;
    wire N__49521;
    wire N__49520;
    wire N__49515;
    wire N__49514;
    wire N__49513;
    wire N__49506;
    wire N__49503;
    wire N__49500;
    wire N__49493;
    wire N__49492;
    wire N__49489;
    wire N__49486;
    wire N__49481;
    wire N__49476;
    wire N__49471;
    wire N__49468;
    wire N__49467;
    wire N__49464;
    wire N__49463;
    wire N__49462;
    wire N__49459;
    wire N__49456;
    wire N__49451;
    wire N__49448;
    wire N__49445;
    wire N__49442;
    wire N__49435;
    wire N__49430;
    wire N__49429;
    wire N__49426;
    wire N__49423;
    wire N__49420;
    wire N__49417;
    wire N__49414;
    wire N__49407;
    wire N__49404;
    wire N__49397;
    wire N__49396;
    wire N__49395;
    wire N__49392;
    wire N__49387;
    wire N__49384;
    wire N__49375;
    wire N__49372;
    wire N__49367;
    wire N__49364;
    wire N__49361;
    wire N__49348;
    wire N__49345;
    wire N__49344;
    wire N__49341;
    wire N__49338;
    wire N__49335;
    wire N__49332;
    wire N__49327;
    wire N__49324;
    wire N__49323;
    wire N__49320;
    wire N__49317;
    wire N__49314;
    wire N__49311;
    wire N__49306;
    wire N__49303;
    wire N__49302;
    wire N__49299;
    wire N__49298;
    wire N__49295;
    wire N__49292;
    wire N__49289;
    wire N__49288;
    wire N__49281;
    wire N__49278;
    wire N__49275;
    wire N__49270;
    wire N__49267;
    wire N__49264;
    wire N__49261;
    wire N__49258;
    wire N__49255;
    wire N__49252;
    wire N__49249;
    wire N__49246;
    wire N__49243;
    wire N__49240;
    wire N__49239;
    wire N__49238;
    wire N__49237;
    wire N__49236;
    wire N__49235;
    wire N__49232;
    wire N__49229;
    wire N__49226;
    wire N__49223;
    wire N__49220;
    wire N__49217;
    wire N__49216;
    wire N__49215;
    wire N__49212;
    wire N__49211;
    wire N__49210;
    wire N__49207;
    wire N__49200;
    wire N__49193;
    wire N__49190;
    wire N__49187;
    wire N__49186;
    wire N__49185;
    wire N__49182;
    wire N__49179;
    wire N__49176;
    wire N__49169;
    wire N__49164;
    wire N__49159;
    wire N__49154;
    wire N__49147;
    wire N__49144;
    wire N__49141;
    wire N__49140;
    wire N__49135;
    wire N__49132;
    wire N__49129;
    wire N__49126;
    wire N__49123;
    wire N__49120;
    wire N__49117;
    wire N__49114;
    wire N__49113;
    wire N__49110;
    wire N__49107;
    wire N__49102;
    wire N__49099;
    wire N__49096;
    wire N__49093;
    wire N__49090;
    wire N__49087;
    wire N__49084;
    wire N__49081;
    wire N__49078;
    wire N__49077;
    wire N__49074;
    wire N__49071;
    wire N__49070;
    wire N__49067;
    wire N__49064;
    wire N__49061;
    wire N__49058;
    wire N__49055;
    wire N__49048;
    wire N__49045;
    wire N__49042;
    wire N__49041;
    wire N__49038;
    wire N__49035;
    wire N__49032;
    wire N__49029;
    wire N__49026;
    wire N__49025;
    wire N__49022;
    wire N__49019;
    wire N__49016;
    wire N__49009;
    wire N__49008;
    wire N__49005;
    wire N__49004;
    wire N__49001;
    wire N__49000;
    wire N__48999;
    wire N__48998;
    wire N__48997;
    wire N__48994;
    wire N__48991;
    wire N__48990;
    wire N__48987;
    wire N__48984;
    wire N__48979;
    wire N__48976;
    wire N__48975;
    wire N__48970;
    wire N__48969;
    wire N__48968;
    wire N__48967;
    wire N__48966;
    wire N__48963;
    wire N__48962;
    wire N__48961;
    wire N__48960;
    wire N__48959;
    wire N__48954;
    wire N__48953;
    wire N__48948;
    wire N__48945;
    wire N__48942;
    wire N__48939;
    wire N__48936;
    wire N__48931;
    wire N__48928;
    wire N__48923;
    wire N__48918;
    wire N__48915;
    wire N__48912;
    wire N__48911;
    wire N__48910;
    wire N__48905;
    wire N__48898;
    wire N__48895;
    wire N__48894;
    wire N__48893;
    wire N__48892;
    wire N__48887;
    wire N__48884;
    wire N__48879;
    wire N__48874;
    wire N__48873;
    wire N__48870;
    wire N__48867;
    wire N__48864;
    wire N__48859;
    wire N__48856;
    wire N__48847;
    wire N__48844;
    wire N__48829;
    wire N__48828;
    wire N__48825;
    wire N__48822;
    wire N__48821;
    wire N__48818;
    wire N__48815;
    wire N__48812;
    wire N__48809;
    wire N__48806;
    wire N__48799;
    wire N__48798;
    wire N__48795;
    wire N__48792;
    wire N__48789;
    wire N__48786;
    wire N__48785;
    wire N__48782;
    wire N__48779;
    wire N__48776;
    wire N__48769;
    wire N__48766;
    wire N__48763;
    wire N__48760;
    wire N__48757;
    wire N__48754;
    wire N__48751;
    wire N__48748;
    wire N__48745;
    wire N__48744;
    wire N__48741;
    wire N__48738;
    wire N__48737;
    wire N__48734;
    wire N__48731;
    wire N__48728;
    wire N__48725;
    wire N__48720;
    wire N__48717;
    wire N__48714;
    wire N__48709;
    wire N__48706;
    wire N__48703;
    wire N__48700;
    wire N__48699;
    wire N__48696;
    wire N__48693;
    wire N__48688;
    wire N__48685;
    wire N__48682;
    wire N__48681;
    wire N__48678;
    wire N__48675;
    wire N__48672;
    wire N__48667;
    wire N__48664;
    wire N__48663;
    wire N__48662;
    wire N__48659;
    wire N__48656;
    wire N__48655;
    wire N__48652;
    wire N__48649;
    wire N__48646;
    wire N__48643;
    wire N__48640;
    wire N__48635;
    wire N__48632;
    wire N__48631;
    wire N__48628;
    wire N__48623;
    wire N__48620;
    wire N__48617;
    wire N__48614;
    wire N__48611;
    wire N__48604;
    wire N__48603;
    wire N__48600;
    wire N__48597;
    wire N__48596;
    wire N__48593;
    wire N__48590;
    wire N__48587;
    wire N__48586;
    wire N__48583;
    wire N__48580;
    wire N__48577;
    wire N__48574;
    wire N__48565;
    wire N__48564;
    wire N__48561;
    wire N__48558;
    wire N__48557;
    wire N__48554;
    wire N__48551;
    wire N__48548;
    wire N__48545;
    wire N__48542;
    wire N__48535;
    wire N__48534;
    wire N__48533;
    wire N__48530;
    wire N__48527;
    wire N__48526;
    wire N__48525;
    wire N__48524;
    wire N__48521;
    wire N__48518;
    wire N__48515;
    wire N__48512;
    wire N__48511;
    wire N__48510;
    wire N__48509;
    wire N__48508;
    wire N__48507;
    wire N__48506;
    wire N__48505;
    wire N__48504;
    wire N__48499;
    wire N__48496;
    wire N__48495;
    wire N__48494;
    wire N__48493;
    wire N__48492;
    wire N__48489;
    wire N__48484;
    wire N__48481;
    wire N__48480;
    wire N__48479;
    wire N__48478;
    wire N__48469;
    wire N__48464;
    wire N__48461;
    wire N__48456;
    wire N__48453;
    wire N__48448;
    wire N__48445;
    wire N__48440;
    wire N__48439;
    wire N__48438;
    wire N__48437;
    wire N__48432;
    wire N__48427;
    wire N__48422;
    wire N__48419;
    wire N__48416;
    wire N__48413;
    wire N__48408;
    wire N__48405;
    wire N__48402;
    wire N__48399;
    wire N__48396;
    wire N__48389;
    wire N__48386;
    wire N__48383;
    wire N__48378;
    wire N__48375;
    wire N__48358;
    wire N__48355;
    wire N__48352;
    wire N__48351;
    wire N__48350;
    wire N__48349;
    wire N__48348;
    wire N__48347;
    wire N__48346;
    wire N__48343;
    wire N__48336;
    wire N__48335;
    wire N__48332;
    wire N__48329;
    wire N__48326;
    wire N__48325;
    wire N__48324;
    wire N__48323;
    wire N__48322;
    wire N__48321;
    wire N__48320;
    wire N__48319;
    wire N__48316;
    wire N__48315;
    wire N__48314;
    wire N__48311;
    wire N__48308;
    wire N__48305;
    wire N__48302;
    wire N__48293;
    wire N__48288;
    wire N__48287;
    wire N__48286;
    wire N__48285;
    wire N__48284;
    wire N__48283;
    wire N__48282;
    wire N__48281;
    wire N__48280;
    wire N__48275;
    wire N__48272;
    wire N__48269;
    wire N__48266;
    wire N__48265;
    wire N__48264;
    wire N__48263;
    wire N__48262;
    wire N__48259;
    wire N__48256;
    wire N__48251;
    wire N__48248;
    wire N__48245;
    wire N__48242;
    wire N__48235;
    wire N__48232;
    wire N__48229;
    wire N__48226;
    wire N__48225;
    wire N__48224;
    wire N__48223;
    wire N__48220;
    wire N__48219;
    wire N__48218;
    wire N__48217;
    wire N__48216;
    wire N__48209;
    wire N__48206;
    wire N__48205;
    wire N__48204;
    wire N__48203;
    wire N__48202;
    wire N__48199;
    wire N__48198;
    wire N__48197;
    wire N__48196;
    wire N__48195;
    wire N__48194;
    wire N__48191;
    wire N__48188;
    wire N__48185;
    wire N__48184;
    wire N__48183;
    wire N__48182;
    wire N__48181;
    wire N__48180;
    wire N__48179;
    wire N__48178;
    wire N__48177;
    wire N__48176;
    wire N__48175;
    wire N__48174;
    wire N__48173;
    wire N__48166;
    wire N__48157;
    wire N__48144;
    wire N__48139;
    wire N__48136;
    wire N__48131;
    wire N__48128;
    wire N__48125;
    wire N__48118;
    wire N__48117;
    wire N__48114;
    wire N__48113;
    wire N__48112;
    wire N__48109;
    wire N__48098;
    wire N__48081;
    wire N__48076;
    wire N__48065;
    wire N__48060;
    wire N__48051;
    wire N__48048;
    wire N__48043;
    wire N__48042;
    wire N__48041;
    wire N__48040;
    wire N__48039;
    wire N__48038;
    wire N__48037;
    wire N__48036;
    wire N__48035;
    wire N__48032;
    wire N__48025;
    wire N__48018;
    wire N__48013;
    wire N__48010;
    wire N__48003;
    wire N__47994;
    wire N__47985;
    wire N__47968;
    wire N__47967;
    wire N__47964;
    wire N__47961;
    wire N__47958;
    wire N__47955;
    wire N__47952;
    wire N__47949;
    wire N__47948;
    wire N__47945;
    wire N__47942;
    wire N__47939;
    wire N__47932;
    wire N__47929;
    wire N__47928;
    wire N__47925;
    wire N__47924;
    wire N__47921;
    wire N__47918;
    wire N__47915;
    wire N__47908;
    wire N__47905;
    wire N__47902;
    wire N__47899;
    wire N__47898;
    wire N__47895;
    wire N__47892;
    wire N__47889;
    wire N__47886;
    wire N__47881;
    wire N__47880;
    wire N__47877;
    wire N__47874;
    wire N__47873;
    wire N__47870;
    wire N__47867;
    wire N__47864;
    wire N__47861;
    wire N__47854;
    wire N__47851;
    wire N__47850;
    wire N__47849;
    wire N__47848;
    wire N__47847;
    wire N__47846;
    wire N__47845;
    wire N__47844;
    wire N__47843;
    wire N__47840;
    wire N__47837;
    wire N__47836;
    wire N__47835;
    wire N__47834;
    wire N__47833;
    wire N__47832;
    wire N__47831;
    wire N__47830;
    wire N__47829;
    wire N__47826;
    wire N__47825;
    wire N__47824;
    wire N__47823;
    wire N__47822;
    wire N__47821;
    wire N__47820;
    wire N__47817;
    wire N__47814;
    wire N__47811;
    wire N__47806;
    wire N__47803;
    wire N__47800;
    wire N__47797;
    wire N__47794;
    wire N__47791;
    wire N__47790;
    wire N__47789;
    wire N__47788;
    wire N__47787;
    wire N__47786;
    wire N__47785;
    wire N__47784;
    wire N__47783;
    wire N__47782;
    wire N__47781;
    wire N__47780;
    wire N__47779;
    wire N__47778;
    wire N__47775;
    wire N__47774;
    wire N__47771;
    wire N__47768;
    wire N__47763;
    wire N__47758;
    wire N__47755;
    wire N__47754;
    wire N__47753;
    wire N__47752;
    wire N__47749;
    wire N__47748;
    wire N__47747;
    wire N__47746;
    wire N__47745;
    wire N__47744;
    wire N__47743;
    wire N__47742;
    wire N__47741;
    wire N__47738;
    wire N__47737;
    wire N__47734;
    wire N__47731;
    wire N__47728;
    wire N__47727;
    wire N__47726;
    wire N__47721;
    wire N__47718;
    wire N__47705;
    wire N__47702;
    wire N__47701;
    wire N__47700;
    wire N__47699;
    wire N__47698;
    wire N__47697;
    wire N__47696;
    wire N__47695;
    wire N__47694;
    wire N__47691;
    wire N__47688;
    wire N__47683;
    wire N__47674;
    wire N__47665;
    wire N__47662;
    wire N__47659;
    wire N__47654;
    wire N__47649;
    wire N__47646;
    wire N__47643;
    wire N__47640;
    wire N__47637;
    wire N__47634;
    wire N__47631;
    wire N__47628;
    wire N__47623;
    wire N__47618;
    wire N__47615;
    wire N__47612;
    wire N__47609;
    wire N__47606;
    wire N__47601;
    wire N__47598;
    wire N__47593;
    wire N__47584;
    wire N__47581;
    wire N__47580;
    wire N__47579;
    wire N__47578;
    wire N__47573;
    wire N__47568;
    wire N__47565;
    wire N__47562;
    wire N__47559;
    wire N__47556;
    wire N__47545;
    wire N__47542;
    wire N__47533;
    wire N__47520;
    wire N__47509;
    wire N__47508;
    wire N__47503;
    wire N__47498;
    wire N__47495;
    wire N__47488;
    wire N__47479;
    wire N__47464;
    wire N__47461;
    wire N__47456;
    wire N__47443;
    wire N__47440;
    wire N__47437;
    wire N__47434;
    wire N__47431;
    wire N__47428;
    wire N__47425;
    wire N__47422;
    wire N__47419;
    wire N__47416;
    wire N__47413;
    wire N__47412;
    wire N__47409;
    wire N__47406;
    wire N__47403;
    wire N__47402;
    wire N__47399;
    wire N__47396;
    wire N__47393;
    wire N__47390;
    wire N__47387;
    wire N__47380;
    wire N__47377;
    wire N__47376;
    wire N__47373;
    wire N__47370;
    wire N__47369;
    wire N__47366;
    wire N__47363;
    wire N__47360;
    wire N__47357;
    wire N__47354;
    wire N__47347;
    wire N__47344;
    wire N__47343;
    wire N__47340;
    wire N__47337;
    wire N__47336;
    wire N__47333;
    wire N__47330;
    wire N__47327;
    wire N__47324;
    wire N__47321;
    wire N__47314;
    wire N__47311;
    wire N__47308;
    wire N__47307;
    wire N__47304;
    wire N__47301;
    wire N__47298;
    wire N__47297;
    wire N__47292;
    wire N__47289;
    wire N__47286;
    wire N__47281;
    wire N__47278;
    wire N__47275;
    wire N__47274;
    wire N__47271;
    wire N__47268;
    wire N__47267;
    wire N__47264;
    wire N__47261;
    wire N__47258;
    wire N__47255;
    wire N__47252;
    wire N__47245;
    wire N__47242;
    wire N__47241;
    wire N__47240;
    wire N__47237;
    wire N__47234;
    wire N__47231;
    wire N__47224;
    wire N__47221;
    wire N__47218;
    wire N__47217;
    wire N__47214;
    wire N__47211;
    wire N__47208;
    wire N__47203;
    wire N__47200;
    wire N__47197;
    wire N__47196;
    wire N__47193;
    wire N__47190;
    wire N__47187;
    wire N__47182;
    wire N__47179;
    wire N__47176;
    wire N__47173;
    wire N__47172;
    wire N__47169;
    wire N__47166;
    wire N__47163;
    wire N__47158;
    wire N__47155;
    wire N__47152;
    wire N__47149;
    wire N__47146;
    wire N__47143;
    wire N__47140;
    wire N__47137;
    wire N__47136;
    wire N__47135;
    wire N__47132;
    wire N__47129;
    wire N__47128;
    wire N__47125;
    wire N__47124;
    wire N__47119;
    wire N__47116;
    wire N__47113;
    wire N__47110;
    wire N__47105;
    wire N__47104;
    wire N__47101;
    wire N__47098;
    wire N__47095;
    wire N__47092;
    wire N__47085;
    wire N__47082;
    wire N__47081;
    wire N__47078;
    wire N__47075;
    wire N__47072;
    wire N__47065;
    wire N__47062;
    wire N__47061;
    wire N__47058;
    wire N__47057;
    wire N__47056;
    wire N__47053;
    wire N__47052;
    wire N__47049;
    wire N__47048;
    wire N__47045;
    wire N__47042;
    wire N__47039;
    wire N__47036;
    wire N__47033;
    wire N__47030;
    wire N__47027;
    wire N__47024;
    wire N__47019;
    wire N__47014;
    wire N__47011;
    wire N__47006;
    wire N__47003;
    wire N__46996;
    wire N__46993;
    wire N__46990;
    wire N__46987;
    wire N__46986;
    wire N__46983;
    wire N__46980;
    wire N__46977;
    wire N__46976;
    wire N__46975;
    wire N__46972;
    wire N__46969;
    wire N__46968;
    wire N__46963;
    wire N__46960;
    wire N__46957;
    wire N__46956;
    wire N__46953;
    wire N__46946;
    wire N__46943;
    wire N__46936;
    wire N__46935;
    wire N__46932;
    wire N__46929;
    wire N__46928;
    wire N__46923;
    wire N__46920;
    wire N__46917;
    wire N__46912;
    wire N__46909;
    wire N__46908;
    wire N__46907;
    wire N__46904;
    wire N__46901;
    wire N__46898;
    wire N__46895;
    wire N__46892;
    wire N__46885;
    wire N__46882;
    wire N__46881;
    wire N__46878;
    wire N__46875;
    wire N__46872;
    wire N__46871;
    wire N__46866;
    wire N__46863;
    wire N__46860;
    wire N__46855;
    wire N__46852;
    wire N__46851;
    wire N__46848;
    wire N__46845;
    wire N__46842;
    wire N__46839;
    wire N__46838;
    wire N__46835;
    wire N__46832;
    wire N__46829;
    wire N__46826;
    wire N__46823;
    wire N__46816;
    wire N__46813;
    wire N__46812;
    wire N__46809;
    wire N__46806;
    wire N__46803;
    wire N__46802;
    wire N__46797;
    wire N__46794;
    wire N__46791;
    wire N__46786;
    wire N__46783;
    wire N__46782;
    wire N__46779;
    wire N__46776;
    wire N__46773;
    wire N__46772;
    wire N__46767;
    wire N__46764;
    wire N__46761;
    wire N__46756;
    wire N__46753;
    wire N__46750;
    wire N__46747;
    wire N__46744;
    wire N__46741;
    wire N__46738;
    wire N__46735;
    wire N__46734;
    wire N__46731;
    wire N__46728;
    wire N__46725;
    wire N__46720;
    wire N__46717;
    wire N__46714;
    wire N__46711;
    wire N__46708;
    wire N__46707;
    wire N__46704;
    wire N__46701;
    wire N__46700;
    wire N__46697;
    wire N__46694;
    wire N__46691;
    wire N__46688;
    wire N__46683;
    wire N__46680;
    wire N__46677;
    wire N__46674;
    wire N__46671;
    wire N__46666;
    wire N__46665;
    wire N__46664;
    wire N__46661;
    wire N__46658;
    wire N__46655;
    wire N__46654;
    wire N__46651;
    wire N__46648;
    wire N__46647;
    wire N__46646;
    wire N__46643;
    wire N__46640;
    wire N__46637;
    wire N__46634;
    wire N__46631;
    wire N__46628;
    wire N__46625;
    wire N__46622;
    wire N__46619;
    wire N__46614;
    wire N__46611;
    wire N__46606;
    wire N__46597;
    wire N__46594;
    wire N__46591;
    wire N__46588;
    wire N__46585;
    wire N__46582;
    wire N__46581;
    wire N__46578;
    wire N__46575;
    wire N__46570;
    wire N__46567;
    wire N__46564;
    wire N__46561;
    wire N__46558;
    wire N__46555;
    wire N__46552;
    wire N__46549;
    wire N__46546;
    wire N__46543;
    wire N__46540;
    wire N__46537;
    wire N__46534;
    wire N__46531;
    wire N__46528;
    wire N__46525;
    wire N__46522;
    wire N__46519;
    wire N__46516;
    wire N__46513;
    wire N__46510;
    wire N__46507;
    wire N__46504;
    wire N__46501;
    wire N__46500;
    wire N__46497;
    wire N__46494;
    wire N__46491;
    wire N__46488;
    wire N__46483;
    wire N__46480;
    wire N__46477;
    wire N__46474;
    wire N__46471;
    wire N__46468;
    wire N__46467;
    wire N__46462;
    wire N__46459;
    wire N__46456;
    wire N__46453;
    wire N__46450;
    wire N__46447;
    wire N__46444;
    wire N__46441;
    wire N__46438;
    wire N__46435;
    wire N__46432;
    wire N__46429;
    wire N__46426;
    wire N__46423;
    wire N__46422;
    wire N__46419;
    wire N__46416;
    wire N__46413;
    wire N__46408;
    wire N__46405;
    wire N__46402;
    wire N__46399;
    wire N__46398;
    wire N__46395;
    wire N__46392;
    wire N__46387;
    wire N__46384;
    wire N__46381;
    wire N__46378;
    wire N__46377;
    wire N__46376;
    wire N__46375;
    wire N__46374;
    wire N__46373;
    wire N__46372;
    wire N__46371;
    wire N__46370;
    wire N__46367;
    wire N__46364;
    wire N__46349;
    wire N__46342;
    wire N__46339;
    wire N__46336;
    wire N__46333;
    wire N__46332;
    wire N__46331;
    wire N__46330;
    wire N__46329;
    wire N__46328;
    wire N__46327;
    wire N__46326;
    wire N__46323;
    wire N__46308;
    wire N__46303;
    wire N__46300;
    wire N__46297;
    wire N__46294;
    wire N__46293;
    wire N__46290;
    wire N__46287;
    wire N__46282;
    wire N__46279;
    wire N__46276;
    wire N__46273;
    wire N__46270;
    wire N__46269;
    wire N__46266;
    wire N__46263;
    wire N__46258;
    wire N__46257;
    wire N__46254;
    wire N__46251;
    wire N__46246;
    wire N__46243;
    wire N__46242;
    wire N__46239;
    wire N__46236;
    wire N__46231;
    wire N__46228;
    wire N__46227;
    wire N__46224;
    wire N__46221;
    wire N__46216;
    wire N__46213;
    wire N__46210;
    wire N__46207;
    wire N__46206;
    wire N__46203;
    wire N__46200;
    wire N__46195;
    wire N__46192;
    wire N__46191;
    wire N__46188;
    wire N__46185;
    wire N__46180;
    wire N__46179;
    wire N__46176;
    wire N__46173;
    wire N__46168;
    wire N__46165;
    wire N__46162;
    wire N__46159;
    wire N__46156;
    wire N__46155;
    wire N__46152;
    wire N__46149;
    wire N__46146;
    wire N__46143;
    wire N__46138;
    wire N__46137;
    wire N__46134;
    wire N__46131;
    wire N__46128;
    wire N__46125;
    wire N__46120;
    wire N__46117;
    wire N__46114;
    wire N__46111;
    wire N__46108;
    wire N__46105;
    wire N__46102;
    wire N__46099;
    wire N__46096;
    wire N__46093;
    wire N__46090;
    wire N__46087;
    wire N__46084;
    wire N__46081;
    wire N__46078;
    wire N__46077;
    wire N__46074;
    wire N__46071;
    wire N__46066;
    wire N__46063;
    wire N__46060;
    wire N__46057;
    wire N__46054;
    wire N__46053;
    wire N__46050;
    wire N__46047;
    wire N__46042;
    wire N__46039;
    wire N__46038;
    wire N__46037;
    wire N__46034;
    wire N__46031;
    wire N__46028;
    wire N__46021;
    wire N__46020;
    wire N__46019;
    wire N__46018;
    wire N__46017;
    wire N__46016;
    wire N__46015;
    wire N__46014;
    wire N__46013;
    wire N__46010;
    wire N__46007;
    wire N__46006;
    wire N__46005;
    wire N__45994;
    wire N__45991;
    wire N__45988;
    wire N__45987;
    wire N__45982;
    wire N__45977;
    wire N__45974;
    wire N__45969;
    wire N__45966;
    wire N__45965;
    wire N__45960;
    wire N__45953;
    wire N__45950;
    wire N__45947;
    wire N__45942;
    wire N__45937;
    wire N__45934;
    wire N__45933;
    wire N__45930;
    wire N__45927;
    wire N__45924;
    wire N__45921;
    wire N__45916;
    wire N__45915;
    wire N__45914;
    wire N__45913;
    wire N__45912;
    wire N__45911;
    wire N__45908;
    wire N__45905;
    wire N__45902;
    wire N__45901;
    wire N__45900;
    wire N__45897;
    wire N__45896;
    wire N__45895;
    wire N__45892;
    wire N__45891;
    wire N__45888;
    wire N__45877;
    wire N__45876;
    wire N__45871;
    wire N__45868;
    wire N__45865;
    wire N__45862;
    wire N__45859;
    wire N__45856;
    wire N__45853;
    wire N__45850;
    wire N__45847;
    wire N__45844;
    wire N__45841;
    wire N__45840;
    wire N__45839;
    wire N__45838;
    wire N__45835;
    wire N__45830;
    wire N__45829;
    wire N__45822;
    wire N__45819;
    wire N__45816;
    wire N__45811;
    wire N__45810;
    wire N__45807;
    wire N__45804;
    wire N__45801;
    wire N__45798;
    wire N__45795;
    wire N__45790;
    wire N__45787;
    wire N__45772;
    wire N__45769;
    wire N__45768;
    wire N__45767;
    wire N__45766;
    wire N__45765;
    wire N__45762;
    wire N__45759;
    wire N__45756;
    wire N__45753;
    wire N__45750;
    wire N__45747;
    wire N__45744;
    wire N__45741;
    wire N__45738;
    wire N__45735;
    wire N__45728;
    wire N__45727;
    wire N__45724;
    wire N__45721;
    wire N__45718;
    wire N__45715;
    wire N__45712;
    wire N__45709;
    wire N__45706;
    wire N__45697;
    wire N__45696;
    wire N__45695;
    wire N__45694;
    wire N__45693;
    wire N__45692;
    wire N__45691;
    wire N__45688;
    wire N__45681;
    wire N__45678;
    wire N__45677;
    wire N__45676;
    wire N__45675;
    wire N__45674;
    wire N__45673;
    wire N__45668;
    wire N__45661;
    wire N__45658;
    wire N__45657;
    wire N__45656;
    wire N__45655;
    wire N__45650;
    wire N__45647;
    wire N__45644;
    wire N__45641;
    wire N__45638;
    wire N__45635;
    wire N__45632;
    wire N__45629;
    wire N__45626;
    wire N__45621;
    wire N__45616;
    wire N__45611;
    wire N__45608;
    wire N__45595;
    wire N__45592;
    wire N__45591;
    wire N__45588;
    wire N__45585;
    wire N__45582;
    wire N__45581;
    wire N__45578;
    wire N__45575;
    wire N__45572;
    wire N__45567;
    wire N__45562;
    wire N__45561;
    wire N__45558;
    wire N__45555;
    wire N__45552;
    wire N__45549;
    wire N__45546;
    wire N__45543;
    wire N__45538;
    wire N__45535;
    wire N__45534;
    wire N__45531;
    wire N__45528;
    wire N__45525;
    wire N__45522;
    wire N__45519;
    wire N__45516;
    wire N__45511;
    wire N__45510;
    wire N__45507;
    wire N__45504;
    wire N__45501;
    wire N__45498;
    wire N__45497;
    wire N__45494;
    wire N__45491;
    wire N__45488;
    wire N__45483;
    wire N__45478;
    wire N__45477;
    wire N__45474;
    wire N__45471;
    wire N__45470;
    wire N__45467;
    wire N__45464;
    wire N__45461;
    wire N__45456;
    wire N__45451;
    wire N__45448;
    wire N__45445;
    wire N__45442;
    wire N__45439;
    wire N__45436;
    wire N__45433;
    wire N__45432;
    wire N__45431;
    wire N__45428;
    wire N__45425;
    wire N__45422;
    wire N__45419;
    wire N__45414;
    wire N__45411;
    wire N__45408;
    wire N__45403;
    wire N__45400;
    wire N__45397;
    wire N__45394;
    wire N__45391;
    wire N__45388;
    wire N__45385;
    wire N__45382;
    wire N__45381;
    wire N__45380;
    wire N__45377;
    wire N__45376;
    wire N__45373;
    wire N__45370;
    wire N__45367;
    wire N__45364;
    wire N__45361;
    wire N__45356;
    wire N__45353;
    wire N__45350;
    wire N__45347;
    wire N__45344;
    wire N__45341;
    wire N__45338;
    wire N__45331;
    wire N__45330;
    wire N__45329;
    wire N__45328;
    wire N__45327;
    wire N__45324;
    wire N__45317;
    wire N__45314;
    wire N__45311;
    wire N__45310;
    wire N__45307;
    wire N__45304;
    wire N__45301;
    wire N__45298;
    wire N__45293;
    wire N__45292;
    wire N__45289;
    wire N__45286;
    wire N__45283;
    wire N__45280;
    wire N__45279;
    wire N__45276;
    wire N__45273;
    wire N__45268;
    wire N__45265;
    wire N__45256;
    wire N__45255;
    wire N__45254;
    wire N__45251;
    wire N__45248;
    wire N__45245;
    wire N__45242;
    wire N__45235;
    wire N__45232;
    wire N__45231;
    wire N__45228;
    wire N__45227;
    wire N__45224;
    wire N__45221;
    wire N__45218;
    wire N__45211;
    wire N__45208;
    wire N__45205;
    wire N__45202;
    wire N__45201;
    wire N__45198;
    wire N__45195;
    wire N__45192;
    wire N__45189;
    wire N__45186;
    wire N__45183;
    wire N__45180;
    wire N__45179;
    wire N__45176;
    wire N__45173;
    wire N__45170;
    wire N__45163;
    wire N__45160;
    wire N__45159;
    wire N__45156;
    wire N__45155;
    wire N__45152;
    wire N__45149;
    wire N__45144;
    wire N__45139;
    wire N__45138;
    wire N__45135;
    wire N__45132;
    wire N__45129;
    wire N__45126;
    wire N__45123;
    wire N__45120;
    wire N__45117;
    wire N__45114;
    wire N__45113;
    wire N__45110;
    wire N__45107;
    wire N__45104;
    wire N__45101;
    wire N__45098;
    wire N__45091;
    wire N__45088;
    wire N__45087;
    wire N__45086;
    wire N__45083;
    wire N__45080;
    wire N__45077;
    wire N__45074;
    wire N__45067;
    wire N__45064;
    wire N__45061;
    wire N__45058;
    wire N__45055;
    wire N__45052;
    wire N__45049;
    wire N__45046;
    wire N__45043;
    wire N__45040;
    wire N__45039;
    wire N__45034;
    wire N__45031;
    wire N__45028;
    wire N__45025;
    wire N__45022;
    wire N__45019;
    wire N__45016;
    wire N__45013;
    wire N__45010;
    wire N__45007;
    wire N__45004;
    wire N__45001;
    wire N__44998;
    wire N__44995;
    wire N__44992;
    wire N__44989;
    wire N__44988;
    wire N__44985;
    wire N__44982;
    wire N__44979;
    wire N__44974;
    wire N__44971;
    wire N__44968;
    wire N__44967;
    wire N__44964;
    wire N__44961;
    wire N__44956;
    wire N__44953;
    wire N__44952;
    wire N__44949;
    wire N__44946;
    wire N__44943;
    wire N__44938;
    wire N__44935;
    wire N__44932;
    wire N__44931;
    wire N__44928;
    wire N__44925;
    wire N__44920;
    wire N__44917;
    wire N__44914;
    wire N__44911;
    wire N__44910;
    wire N__44907;
    wire N__44906;
    wire N__44903;
    wire N__44902;
    wire N__44899;
    wire N__44896;
    wire N__44893;
    wire N__44890;
    wire N__44887;
    wire N__44884;
    wire N__44879;
    wire N__44872;
    wire N__44871;
    wire N__44868;
    wire N__44865;
    wire N__44862;
    wire N__44857;
    wire N__44854;
    wire N__44851;
    wire N__44850;
    wire N__44849;
    wire N__44848;
    wire N__44847;
    wire N__44846;
    wire N__44843;
    wire N__44840;
    wire N__44837;
    wire N__44834;
    wire N__44831;
    wire N__44828;
    wire N__44825;
    wire N__44822;
    wire N__44819;
    wire N__44812;
    wire N__44809;
    wire N__44806;
    wire N__44801;
    wire N__44800;
    wire N__44799;
    wire N__44796;
    wire N__44793;
    wire N__44790;
    wire N__44785;
    wire N__44782;
    wire N__44779;
    wire N__44776;
    wire N__44767;
    wire N__44764;
    wire N__44761;
    wire N__44758;
    wire N__44755;
    wire N__44754;
    wire N__44751;
    wire N__44748;
    wire N__44745;
    wire N__44744;
    wire N__44741;
    wire N__44738;
    wire N__44735;
    wire N__44732;
    wire N__44725;
    wire N__44722;
    wire N__44719;
    wire N__44718;
    wire N__44717;
    wire N__44714;
    wire N__44709;
    wire N__44704;
    wire N__44703;
    wire N__44700;
    wire N__44697;
    wire N__44692;
    wire N__44689;
    wire N__44688;
    wire N__44685;
    wire N__44682;
    wire N__44679;
    wire N__44674;
    wire N__44671;
    wire N__44670;
    wire N__44667;
    wire N__44664;
    wire N__44661;
    wire N__44656;
    wire N__44653;
    wire N__44650;
    wire N__44649;
    wire N__44646;
    wire N__44643;
    wire N__44640;
    wire N__44635;
    wire N__44632;
    wire N__44631;
    wire N__44628;
    wire N__44625;
    wire N__44620;
    wire N__44617;
    wire N__44616;
    wire N__44613;
    wire N__44610;
    wire N__44605;
    wire N__44602;
    wire N__44601;
    wire N__44598;
    wire N__44595;
    wire N__44590;
    wire N__44587;
    wire N__44586;
    wire N__44583;
    wire N__44580;
    wire N__44575;
    wire N__44572;
    wire N__44571;
    wire N__44568;
    wire N__44565;
    wire N__44562;
    wire N__44557;
    wire N__44554;
    wire N__44553;
    wire N__44550;
    wire N__44547;
    wire N__44542;
    wire N__44539;
    wire N__44536;
    wire N__44535;
    wire N__44532;
    wire N__44529;
    wire N__44524;
    wire N__44521;
    wire N__44520;
    wire N__44517;
    wire N__44514;
    wire N__44509;
    wire N__44506;
    wire N__44505;
    wire N__44502;
    wire N__44499;
    wire N__44496;
    wire N__44491;
    wire N__44488;
    wire N__44487;
    wire N__44484;
    wire N__44481;
    wire N__44476;
    wire N__44473;
    wire N__44472;
    wire N__44469;
    wire N__44466;
    wire N__44463;
    wire N__44458;
    wire N__44455;
    wire N__44454;
    wire N__44451;
    wire N__44448;
    wire N__44443;
    wire N__44440;
    wire N__44437;
    wire N__44434;
    wire N__44431;
    wire N__44428;
    wire N__44425;
    wire N__44422;
    wire N__44419;
    wire N__44418;
    wire N__44415;
    wire N__44412;
    wire N__44411;
    wire N__44408;
    wire N__44405;
    wire N__44402;
    wire N__44401;
    wire N__44400;
    wire N__44397;
    wire N__44392;
    wire N__44389;
    wire N__44386;
    wire N__44379;
    wire N__44374;
    wire N__44371;
    wire N__44368;
    wire N__44365;
    wire N__44362;
    wire N__44359;
    wire N__44356;
    wire N__44353;
    wire N__44350;
    wire N__44347;
    wire N__44344;
    wire N__44341;
    wire N__44338;
    wire N__44335;
    wire N__44332;
    wire N__44329;
    wire N__44326;
    wire N__44323;
    wire N__44322;
    wire N__44319;
    wire N__44316;
    wire N__44311;
    wire N__44310;
    wire N__44307;
    wire N__44304;
    wire N__44301;
    wire N__44298;
    wire N__44295;
    wire N__44292;
    wire N__44287;
    wire N__44284;
    wire N__44283;
    wire N__44282;
    wire N__44279;
    wire N__44276;
    wire N__44273;
    wire N__44272;
    wire N__44271;
    wire N__44270;
    wire N__44263;
    wire N__44260;
    wire N__44257;
    wire N__44254;
    wire N__44251;
    wire N__44242;
    wire N__44239;
    wire N__44236;
    wire N__44233;
    wire N__44232;
    wire N__44231;
    wire N__44228;
    wire N__44225;
    wire N__44222;
    wire N__44219;
    wire N__44216;
    wire N__44213;
    wire N__44210;
    wire N__44207;
    wire N__44204;
    wire N__44197;
    wire N__44194;
    wire N__44191;
    wire N__44188;
    wire N__44185;
    wire N__44182;
    wire N__44179;
    wire N__44176;
    wire N__44173;
    wire N__44170;
    wire N__44167;
    wire N__44164;
    wire N__44161;
    wire N__44158;
    wire N__44155;
    wire N__44152;
    wire N__44149;
    wire N__44148;
    wire N__44147;
    wire N__44146;
    wire N__44143;
    wire N__44140;
    wire N__44137;
    wire N__44134;
    wire N__44131;
    wire N__44128;
    wire N__44127;
    wire N__44124;
    wire N__44121;
    wire N__44116;
    wire N__44113;
    wire N__44112;
    wire N__44109;
    wire N__44108;
    wire N__44107;
    wire N__44104;
    wire N__44101;
    wire N__44098;
    wire N__44095;
    wire N__44092;
    wire N__44089;
    wire N__44086;
    wire N__44085;
    wire N__44084;
    wire N__44081;
    wire N__44076;
    wire N__44073;
    wire N__44066;
    wire N__44061;
    wire N__44058;
    wire N__44053;
    wire N__44050;
    wire N__44047;
    wire N__44040;
    wire N__44035;
    wire N__44032;
    wire N__44031;
    wire N__44028;
    wire N__44025;
    wire N__44022;
    wire N__44019;
    wire N__44016;
    wire N__44013;
    wire N__44010;
    wire N__44009;
    wire N__44006;
    wire N__44003;
    wire N__44000;
    wire N__43997;
    wire N__43990;
    wire N__43987;
    wire N__43984;
    wire N__43981;
    wire N__43980;
    wire N__43977;
    wire N__43974;
    wire N__43969;
    wire N__43966;
    wire N__43963;
    wire N__43960;
    wire N__43957;
    wire N__43954;
    wire N__43951;
    wire N__43948;
    wire N__43945;
    wire N__43942;
    wire N__43939;
    wire N__43936;
    wire N__43933;
    wire N__43930;
    wire N__43927;
    wire N__43924;
    wire N__43923;
    wire N__43920;
    wire N__43917;
    wire N__43914;
    wire N__43911;
    wire N__43908;
    wire N__43905;
    wire N__43902;
    wire N__43899;
    wire N__43896;
    wire N__43893;
    wire N__43890;
    wire N__43887;
    wire N__43884;
    wire N__43881;
    wire N__43878;
    wire N__43873;
    wire N__43872;
    wire N__43871;
    wire N__43866;
    wire N__43865;
    wire N__43864;
    wire N__43861;
    wire N__43858;
    wire N__43855;
    wire N__43852;
    wire N__43849;
    wire N__43848;
    wire N__43847;
    wire N__43842;
    wire N__43837;
    wire N__43834;
    wire N__43831;
    wire N__43822;
    wire N__43821;
    wire N__43818;
    wire N__43817;
    wire N__43816;
    wire N__43813;
    wire N__43810;
    wire N__43807;
    wire N__43806;
    wire N__43803;
    wire N__43802;
    wire N__43797;
    wire N__43796;
    wire N__43793;
    wire N__43790;
    wire N__43787;
    wire N__43784;
    wire N__43781;
    wire N__43778;
    wire N__43775;
    wire N__43772;
    wire N__43769;
    wire N__43768;
    wire N__43761;
    wire N__43760;
    wire N__43755;
    wire N__43752;
    wire N__43749;
    wire N__43746;
    wire N__43743;
    wire N__43740;
    wire N__43735;
    wire N__43732;
    wire N__43729;
    wire N__43726;
    wire N__43723;
    wire N__43720;
    wire N__43711;
    wire N__43710;
    wire N__43707;
    wire N__43704;
    wire N__43701;
    wire N__43698;
    wire N__43695;
    wire N__43692;
    wire N__43687;
    wire N__43686;
    wire N__43685;
    wire N__43678;
    wire N__43677;
    wire N__43674;
    wire N__43673;
    wire N__43670;
    wire N__43667;
    wire N__43664;
    wire N__43661;
    wire N__43658;
    wire N__43655;
    wire N__43652;
    wire N__43645;
    wire N__43642;
    wire N__43641;
    wire N__43638;
    wire N__43635;
    wire N__43630;
    wire N__43627;
    wire N__43624;
    wire N__43621;
    wire N__43618;
    wire N__43615;
    wire N__43612;
    wire N__43609;
    wire N__43606;
    wire N__43603;
    wire N__43600;
    wire N__43597;
    wire N__43594;
    wire N__43591;
    wire N__43588;
    wire N__43585;
    wire N__43582;
    wire N__43579;
    wire N__43576;
    wire N__43573;
    wire N__43570;
    wire N__43569;
    wire N__43566;
    wire N__43563;
    wire N__43562;
    wire N__43559;
    wire N__43556;
    wire N__43553;
    wire N__43546;
    wire N__43545;
    wire N__43542;
    wire N__43539;
    wire N__43534;
    wire N__43533;
    wire N__43532;
    wire N__43529;
    wire N__43526;
    wire N__43525;
    wire N__43524;
    wire N__43521;
    wire N__43520;
    wire N__43517;
    wire N__43514;
    wire N__43511;
    wire N__43508;
    wire N__43505;
    wire N__43504;
    wire N__43501;
    wire N__43496;
    wire N__43493;
    wire N__43488;
    wire N__43487;
    wire N__43484;
    wire N__43481;
    wire N__43478;
    wire N__43475;
    wire N__43474;
    wire N__43471;
    wire N__43468;
    wire N__43465;
    wire N__43462;
    wire N__43461;
    wire N__43456;
    wire N__43453;
    wire N__43450;
    wire N__43447;
    wire N__43444;
    wire N__43441;
    wire N__43438;
    wire N__43435;
    wire N__43428;
    wire N__43417;
    wire N__43414;
    wire N__43413;
    wire N__43410;
    wire N__43409;
    wire N__43406;
    wire N__43403;
    wire N__43400;
    wire N__43397;
    wire N__43390;
    wire N__43387;
    wire N__43384;
    wire N__43383;
    wire N__43382;
    wire N__43379;
    wire N__43376;
    wire N__43375;
    wire N__43374;
    wire N__43371;
    wire N__43366;
    wire N__43363;
    wire N__43360;
    wire N__43357;
    wire N__43354;
    wire N__43351;
    wire N__43348;
    wire N__43347;
    wire N__43344;
    wire N__43339;
    wire N__43336;
    wire N__43333;
    wire N__43328;
    wire N__43321;
    wire N__43320;
    wire N__43319;
    wire N__43316;
    wire N__43313;
    wire N__43310;
    wire N__43305;
    wire N__43300;
    wire N__43299;
    wire N__43296;
    wire N__43295;
    wire N__43292;
    wire N__43291;
    wire N__43288;
    wire N__43285;
    wire N__43284;
    wire N__43281;
    wire N__43278;
    wire N__43277;
    wire N__43276;
    wire N__43275;
    wire N__43274;
    wire N__43273;
    wire N__43268;
    wire N__43265;
    wire N__43260;
    wire N__43257;
    wire N__43254;
    wire N__43249;
    wire N__43246;
    wire N__43243;
    wire N__43228;
    wire N__43225;
    wire N__43222;
    wire N__43219;
    wire N__43218;
    wire N__43213;
    wire N__43210;
    wire N__43207;
    wire N__43204;
    wire N__43201;
    wire N__43198;
    wire N__43195;
    wire N__43192;
    wire N__43189;
    wire N__43186;
    wire N__43183;
    wire N__43180;
    wire N__43177;
    wire N__43174;
    wire N__43171;
    wire N__43168;
    wire N__43165;
    wire N__43162;
    wire N__43159;
    wire N__43158;
    wire N__43155;
    wire N__43152;
    wire N__43149;
    wire N__43146;
    wire N__43143;
    wire N__43140;
    wire N__43137;
    wire N__43134;
    wire N__43131;
    wire N__43128;
    wire N__43125;
    wire N__43122;
    wire N__43119;
    wire N__43116;
    wire N__43113;
    wire N__43108;
    wire N__43105;
    wire N__43104;
    wire N__43101;
    wire N__43098;
    wire N__43097;
    wire N__43094;
    wire N__43091;
    wire N__43088;
    wire N__43085;
    wire N__43082;
    wire N__43079;
    wire N__43076;
    wire N__43073;
    wire N__43066;
    wire N__43065;
    wire N__43062;
    wire N__43059;
    wire N__43056;
    wire N__43055;
    wire N__43050;
    wire N__43047;
    wire N__43044;
    wire N__43039;
    wire N__43038;
    wire N__43035;
    wire N__43032;
    wire N__43029;
    wire N__43024;
    wire N__43023;
    wire N__43020;
    wire N__43017;
    wire N__43014;
    wire N__43009;
    wire N__43006;
    wire N__43003;
    wire N__43000;
    wire N__42997;
    wire N__42994;
    wire N__42991;
    wire N__42988;
    wire N__42985;
    wire N__42982;
    wire N__42979;
    wire N__42976;
    wire N__42973;
    wire N__42970;
    wire N__42967;
    wire N__42966;
    wire N__42963;
    wire N__42960;
    wire N__42957;
    wire N__42954;
    wire N__42951;
    wire N__42948;
    wire N__42945;
    wire N__42942;
    wire N__42939;
    wire N__42936;
    wire N__42933;
    wire N__42930;
    wire N__42927;
    wire N__42924;
    wire N__42921;
    wire N__42916;
    wire N__42915;
    wire N__42912;
    wire N__42909;
    wire N__42906;
    wire N__42901;
    wire N__42898;
    wire N__42895;
    wire N__42892;
    wire N__42889;
    wire N__42886;
    wire N__42885;
    wire N__42882;
    wire N__42879;
    wire N__42874;
    wire N__42873;
    wire N__42870;
    wire N__42867;
    wire N__42864;
    wire N__42859;
    wire N__42856;
    wire N__42855;
    wire N__42852;
    wire N__42849;
    wire N__42846;
    wire N__42841;
    wire N__42840;
    wire N__42839;
    wire N__42836;
    wire N__42833;
    wire N__42830;
    wire N__42823;
    wire N__42822;
    wire N__42819;
    wire N__42816;
    wire N__42815;
    wire N__42812;
    wire N__42809;
    wire N__42808;
    wire N__42805;
    wire N__42804;
    wire N__42801;
    wire N__42798;
    wire N__42795;
    wire N__42792;
    wire N__42789;
    wire N__42788;
    wire N__42785;
    wire N__42782;
    wire N__42779;
    wire N__42774;
    wire N__42771;
    wire N__42768;
    wire N__42759;
    wire N__42754;
    wire N__42753;
    wire N__42750;
    wire N__42747;
    wire N__42746;
    wire N__42743;
    wire N__42740;
    wire N__42737;
    wire N__42732;
    wire N__42727;
    wire N__42726;
    wire N__42725;
    wire N__42720;
    wire N__42717;
    wire N__42712;
    wire N__42711;
    wire N__42708;
    wire N__42705;
    wire N__42702;
    wire N__42701;
    wire N__42698;
    wire N__42695;
    wire N__42692;
    wire N__42689;
    wire N__42682;
    wire N__42679;
    wire N__42678;
    wire N__42677;
    wire N__42674;
    wire N__42671;
    wire N__42668;
    wire N__42663;
    wire N__42658;
    wire N__42655;
    wire N__42654;
    wire N__42651;
    wire N__42648;
    wire N__42645;
    wire N__42644;
    wire N__42641;
    wire N__42638;
    wire N__42635;
    wire N__42632;
    wire N__42625;
    wire N__42624;
    wire N__42623;
    wire N__42620;
    wire N__42619;
    wire N__42616;
    wire N__42615;
    wire N__42612;
    wire N__42609;
    wire N__42606;
    wire N__42603;
    wire N__42600;
    wire N__42597;
    wire N__42596;
    wire N__42593;
    wire N__42590;
    wire N__42587;
    wire N__42584;
    wire N__42581;
    wire N__42578;
    wire N__42575;
    wire N__42570;
    wire N__42567;
    wire N__42562;
    wire N__42559;
    wire N__42556;
    wire N__42551;
    wire N__42544;
    wire N__42543;
    wire N__42540;
    wire N__42537;
    wire N__42534;
    wire N__42531;
    wire N__42530;
    wire N__42527;
    wire N__42524;
    wire N__42521;
    wire N__42518;
    wire N__42515;
    wire N__42508;
    wire N__42507;
    wire N__42506;
    wire N__42503;
    wire N__42500;
    wire N__42497;
    wire N__42490;
    wire N__42489;
    wire N__42484;
    wire N__42481;
    wire N__42478;
    wire N__42475;
    wire N__42472;
    wire N__42471;
    wire N__42468;
    wire N__42465;
    wire N__42460;
    wire N__42459;
    wire N__42456;
    wire N__42453;
    wire N__42450;
    wire N__42447;
    wire N__42444;
    wire N__42439;
    wire N__42436;
    wire N__42435;
    wire N__42432;
    wire N__42429;
    wire N__42426;
    wire N__42423;
    wire N__42420;
    wire N__42417;
    wire N__42412;
    wire N__42409;
    wire N__42408;
    wire N__42405;
    wire N__42402;
    wire N__42397;
    wire N__42396;
    wire N__42393;
    wire N__42390;
    wire N__42387;
    wire N__42382;
    wire N__42381;
    wire N__42376;
    wire N__42373;
    wire N__42370;
    wire N__42367;
    wire N__42364;
    wire N__42361;
    wire N__42358;
    wire N__42357;
    wire N__42354;
    wire N__42353;
    wire N__42350;
    wire N__42347;
    wire N__42346;
    wire N__42345;
    wire N__42344;
    wire N__42343;
    wire N__42342;
    wire N__42341;
    wire N__42340;
    wire N__42339;
    wire N__42336;
    wire N__42333;
    wire N__42330;
    wire N__42327;
    wire N__42324;
    wire N__42321;
    wire N__42318;
    wire N__42315;
    wire N__42312;
    wire N__42309;
    wire N__42306;
    wire N__42303;
    wire N__42300;
    wire N__42297;
    wire N__42288;
    wire N__42279;
    wire N__42268;
    wire N__42265;
    wire N__42262;
    wire N__42259;
    wire N__42256;
    wire N__42253;
    wire N__42250;
    wire N__42247;
    wire N__42244;
    wire N__42241;
    wire N__42238;
    wire N__42235;
    wire N__42232;
    wire N__42229;
    wire N__42226;
    wire N__42223;
    wire N__42220;
    wire N__42217;
    wire N__42216;
    wire N__42213;
    wire N__42210;
    wire N__42207;
    wire N__42204;
    wire N__42201;
    wire N__42198;
    wire N__42195;
    wire N__42192;
    wire N__42189;
    wire N__42186;
    wire N__42183;
    wire N__42180;
    wire N__42177;
    wire N__42172;
    wire N__42169;
    wire N__42166;
    wire N__42163;
    wire N__42160;
    wire N__42157;
    wire N__42154;
    wire N__42151;
    wire N__42148;
    wire N__42145;
    wire N__42144;
    wire N__42143;
    wire N__42140;
    wire N__42139;
    wire N__42136;
    wire N__42135;
    wire N__42132;
    wire N__42127;
    wire N__42126;
    wire N__42123;
    wire N__42120;
    wire N__42119;
    wire N__42116;
    wire N__42113;
    wire N__42110;
    wire N__42105;
    wire N__42102;
    wire N__42095;
    wire N__42090;
    wire N__42087;
    wire N__42084;
    wire N__42081;
    wire N__42076;
    wire N__42075;
    wire N__42074;
    wire N__42071;
    wire N__42068;
    wire N__42065;
    wire N__42062;
    wire N__42057;
    wire N__42054;
    wire N__42051;
    wire N__42046;
    wire N__42045;
    wire N__42044;
    wire N__42041;
    wire N__42038;
    wire N__42035;
    wire N__42030;
    wire N__42025;
    wire N__42024;
    wire N__42021;
    wire N__42020;
    wire N__42019;
    wire N__42016;
    wire N__42009;
    wire N__42008;
    wire N__42007;
    wire N__42006;
    wire N__42005;
    wire N__42004;
    wire N__42001;
    wire N__41998;
    wire N__41993;
    wire N__41992;
    wire N__41991;
    wire N__41990;
    wire N__41989;
    wire N__41988;
    wire N__41987;
    wire N__41980;
    wire N__41973;
    wire N__41968;
    wire N__41959;
    wire N__41950;
    wire N__41947;
    wire N__41944;
    wire N__41943;
    wire N__41940;
    wire N__41937;
    wire N__41932;
    wire N__41929;
    wire N__41926;
    wire N__41923;
    wire N__41920;
    wire N__41917;
    wire N__41914;
    wire N__41913;
    wire N__41912;
    wire N__41909;
    wire N__41904;
    wire N__41899;
    wire N__41896;
    wire N__41895;
    wire N__41892;
    wire N__41891;
    wire N__41888;
    wire N__41885;
    wire N__41882;
    wire N__41875;
    wire N__41872;
    wire N__41869;
    wire N__41866;
    wire N__41863;
    wire N__41862;
    wire N__41861;
    wire N__41858;
    wire N__41855;
    wire N__41852;
    wire N__41847;
    wire N__41842;
    wire N__41841;
    wire N__41836;
    wire N__41833;
    wire N__41830;
    wire N__41827;
    wire N__41826;
    wire N__41825;
    wire N__41822;
    wire N__41819;
    wire N__41816;
    wire N__41813;
    wire N__41808;
    wire N__41805;
    wire N__41802;
    wire N__41797;
    wire N__41796;
    wire N__41791;
    wire N__41788;
    wire N__41785;
    wire N__41782;
    wire N__41781;
    wire N__41778;
    wire N__41775;
    wire N__41772;
    wire N__41769;
    wire N__41766;
    wire N__41763;
    wire N__41760;
    wire N__41757;
    wire N__41752;
    wire N__41751;
    wire N__41748;
    wire N__41745;
    wire N__41744;
    wire N__41741;
    wire N__41738;
    wire N__41735;
    wire N__41732;
    wire N__41729;
    wire N__41722;
    wire N__41719;
    wire N__41718;
    wire N__41715;
    wire N__41714;
    wire N__41711;
    wire N__41708;
    wire N__41705;
    wire N__41698;
    wire N__41695;
    wire N__41692;
    wire N__41691;
    wire N__41688;
    wire N__41685;
    wire N__41684;
    wire N__41681;
    wire N__41678;
    wire N__41675;
    wire N__41672;
    wire N__41669;
    wire N__41664;
    wire N__41661;
    wire N__41656;
    wire N__41653;
    wire N__41650;
    wire N__41647;
    wire N__41646;
    wire N__41643;
    wire N__41642;
    wire N__41639;
    wire N__41636;
    wire N__41633;
    wire N__41626;
    wire N__41623;
    wire N__41622;
    wire N__41619;
    wire N__41616;
    wire N__41615;
    wire N__41614;
    wire N__41609;
    wire N__41606;
    wire N__41603;
    wire N__41596;
    wire N__41593;
    wire N__41592;
    wire N__41591;
    wire N__41588;
    wire N__41585;
    wire N__41582;
    wire N__41579;
    wire N__41576;
    wire N__41569;
    wire N__41566;
    wire N__41565;
    wire N__41562;
    wire N__41561;
    wire N__41558;
    wire N__41555;
    wire N__41552;
    wire N__41545;
    wire N__41544;
    wire N__41541;
    wire N__41536;
    wire N__41535;
    wire N__41532;
    wire N__41529;
    wire N__41528;
    wire N__41527;
    wire N__41526;
    wire N__41523;
    wire N__41518;
    wire N__41515;
    wire N__41512;
    wire N__41507;
    wire N__41506;
    wire N__41503;
    wire N__41500;
    wire N__41497;
    wire N__41494;
    wire N__41491;
    wire N__41488;
    wire N__41485;
    wire N__41482;
    wire N__41477;
    wire N__41470;
    wire N__41469;
    wire N__41466;
    wire N__41463;
    wire N__41460;
    wire N__41457;
    wire N__41452;
    wire N__41449;
    wire N__41446;
    wire N__41443;
    wire N__41440;
    wire N__41437;
    wire N__41436;
    wire N__41433;
    wire N__41430;
    wire N__41427;
    wire N__41426;
    wire N__41425;
    wire N__41422;
    wire N__41419;
    wire N__41416;
    wire N__41413;
    wire N__41410;
    wire N__41405;
    wire N__41402;
    wire N__41399;
    wire N__41396;
    wire N__41393;
    wire N__41390;
    wire N__41387;
    wire N__41386;
    wire N__41383;
    wire N__41378;
    wire N__41375;
    wire N__41372;
    wire N__41365;
    wire N__41364;
    wire N__41363;
    wire N__41360;
    wire N__41357;
    wire N__41356;
    wire N__41355;
    wire N__41354;
    wire N__41351;
    wire N__41348;
    wire N__41347;
    wire N__41342;
    wire N__41339;
    wire N__41336;
    wire N__41333;
    wire N__41330;
    wire N__41327;
    wire N__41324;
    wire N__41321;
    wire N__41318;
    wire N__41315;
    wire N__41312;
    wire N__41309;
    wire N__41306;
    wire N__41303;
    wire N__41300;
    wire N__41293;
    wire N__41284;
    wire N__41283;
    wire N__41280;
    wire N__41277;
    wire N__41274;
    wire N__41269;
    wire N__41266;
    wire N__41263;
    wire N__41260;
    wire N__41259;
    wire N__41256;
    wire N__41253;
    wire N__41248;
    wire N__41245;
    wire N__41242;
    wire N__41239;
    wire N__41236;
    wire N__41233;
    wire N__41230;
    wire N__41227;
    wire N__41224;
    wire N__41221;
    wire N__41218;
    wire N__41215;
    wire N__41212;
    wire N__41209;
    wire N__41206;
    wire N__41203;
    wire N__41200;
    wire N__41197;
    wire N__41196;
    wire N__41193;
    wire N__41190;
    wire N__41189;
    wire N__41186;
    wire N__41183;
    wire N__41180;
    wire N__41177;
    wire N__41170;
    wire N__41169;
    wire N__41166;
    wire N__41165;
    wire N__41164;
    wire N__41161;
    wire N__41158;
    wire N__41153;
    wire N__41150;
    wire N__41143;
    wire N__41142;
    wire N__41141;
    wire N__41138;
    wire N__41135;
    wire N__41134;
    wire N__41133;
    wire N__41132;
    wire N__41131;
    wire N__41130;
    wire N__41129;
    wire N__41126;
    wire N__41123;
    wire N__41120;
    wire N__41117;
    wire N__41116;
    wire N__41115;
    wire N__41112;
    wire N__41109;
    wire N__41106;
    wire N__41103;
    wire N__41100;
    wire N__41099;
    wire N__41098;
    wire N__41097;
    wire N__41094;
    wire N__41087;
    wire N__41084;
    wire N__41083;
    wire N__41082;
    wire N__41081;
    wire N__41080;
    wire N__41079;
    wire N__41076;
    wire N__41073;
    wire N__41070;
    wire N__41067;
    wire N__41062;
    wire N__41059;
    wire N__41056;
    wire N__41053;
    wire N__41046;
    wire N__41043;
    wire N__41040;
    wire N__41037;
    wire N__41034;
    wire N__41031;
    wire N__41026;
    wire N__41017;
    wire N__41012;
    wire N__41009;
    wire N__41006;
    wire N__41003;
    wire N__41000;
    wire N__40997;
    wire N__40994;
    wire N__40987;
    wire N__40984;
    wire N__40979;
    wire N__40970;
    wire N__40967;
    wire N__40962;
    wire N__40961;
    wire N__40958;
    wire N__40955;
    wire N__40952;
    wire N__40945;
    wire N__40942;
    wire N__40939;
    wire N__40938;
    wire N__40935;
    wire N__40932;
    wire N__40929;
    wire N__40928;
    wire N__40925;
    wire N__40922;
    wire N__40919;
    wire N__40916;
    wire N__40913;
    wire N__40910;
    wire N__40907;
    wire N__40906;
    wire N__40901;
    wire N__40898;
    wire N__40895;
    wire N__40888;
    wire N__40885;
    wire N__40882;
    wire N__40881;
    wire N__40878;
    wire N__40875;
    wire N__40872;
    wire N__40869;
    wire N__40864;
    wire N__40861;
    wire N__40860;
    wire N__40857;
    wire N__40854;
    wire N__40853;
    wire N__40850;
    wire N__40847;
    wire N__40844;
    wire N__40841;
    wire N__40838;
    wire N__40831;
    wire N__40828;
    wire N__40825;
    wire N__40822;
    wire N__40819;
    wire N__40816;
    wire N__40813;
    wire N__40810;
    wire N__40807;
    wire N__40804;
    wire N__40801;
    wire N__40798;
    wire N__40795;
    wire N__40792;
    wire N__40789;
    wire N__40786;
    wire N__40785;
    wire N__40784;
    wire N__40781;
    wire N__40778;
    wire N__40775;
    wire N__40772;
    wire N__40769;
    wire N__40766;
    wire N__40763;
    wire N__40760;
    wire N__40757;
    wire N__40750;
    wire N__40747;
    wire N__40744;
    wire N__40741;
    wire N__40738;
    wire N__40735;
    wire N__40732;
    wire N__40729;
    wire N__40726;
    wire N__40723;
    wire N__40720;
    wire N__40717;
    wire N__40714;
    wire N__40711;
    wire N__40708;
    wire N__40705;
    wire N__40702;
    wire N__40699;
    wire N__40696;
    wire N__40693;
    wire N__40690;
    wire N__40687;
    wire N__40684;
    wire N__40683;
    wire N__40680;
    wire N__40677;
    wire N__40674;
    wire N__40671;
    wire N__40668;
    wire N__40665;
    wire N__40660;
    wire N__40657;
    wire N__40654;
    wire N__40651;
    wire N__40648;
    wire N__40645;
    wire N__40642;
    wire N__40641;
    wire N__40638;
    wire N__40635;
    wire N__40632;
    wire N__40629;
    wire N__40626;
    wire N__40621;
    wire N__40618;
    wire N__40615;
    wire N__40612;
    wire N__40609;
    wire N__40606;
    wire N__40603;
    wire N__40600;
    wire N__40597;
    wire N__40594;
    wire N__40591;
    wire N__40588;
    wire N__40585;
    wire N__40582;
    wire N__40579;
    wire N__40576;
    wire N__40573;
    wire N__40570;
    wire N__40567;
    wire N__40564;
    wire N__40561;
    wire N__40558;
    wire N__40555;
    wire N__40552;
    wire N__40551;
    wire N__40548;
    wire N__40545;
    wire N__40542;
    wire N__40539;
    wire N__40536;
    wire N__40533;
    wire N__40530;
    wire N__40527;
    wire N__40524;
    wire N__40523;
    wire N__40520;
    wire N__40517;
    wire N__40514;
    wire N__40511;
    wire N__40508;
    wire N__40501;
    wire N__40498;
    wire N__40495;
    wire N__40492;
    wire N__40489;
    wire N__40486;
    wire N__40483;
    wire N__40480;
    wire N__40477;
    wire N__40474;
    wire N__40471;
    wire N__40468;
    wire N__40465;
    wire N__40462;
    wire N__40459;
    wire N__40456;
    wire N__40453;
    wire N__40450;
    wire N__40447;
    wire N__40446;
    wire N__40443;
    wire N__40440;
    wire N__40437;
    wire N__40434;
    wire N__40431;
    wire N__40428;
    wire N__40425;
    wire N__40422;
    wire N__40419;
    wire N__40416;
    wire N__40413;
    wire N__40412;
    wire N__40409;
    wire N__40406;
    wire N__40403;
    wire N__40400;
    wire N__40397;
    wire N__40390;
    wire N__40387;
    wire N__40384;
    wire N__40381;
    wire N__40378;
    wire N__40375;
    wire N__40374;
    wire N__40373;
    wire N__40370;
    wire N__40367;
    wire N__40364;
    wire N__40361;
    wire N__40358;
    wire N__40355;
    wire N__40352;
    wire N__40349;
    wire N__40342;
    wire N__40339;
    wire N__40336;
    wire N__40333;
    wire N__40330;
    wire N__40329;
    wire N__40326;
    wire N__40323;
    wire N__40320;
    wire N__40317;
    wire N__40316;
    wire N__40315;
    wire N__40314;
    wire N__40311;
    wire N__40308;
    wire N__40305;
    wire N__40302;
    wire N__40299;
    wire N__40288;
    wire N__40285;
    wire N__40282;
    wire N__40279;
    wire N__40276;
    wire N__40275;
    wire N__40274;
    wire N__40271;
    wire N__40266;
    wire N__40261;
    wire N__40260;
    wire N__40257;
    wire N__40256;
    wire N__40253;
    wire N__40250;
    wire N__40247;
    wire N__40242;
    wire N__40239;
    wire N__40234;
    wire N__40231;
    wire N__40230;
    wire N__40229;
    wire N__40226;
    wire N__40223;
    wire N__40220;
    wire N__40213;
    wire N__40210;
    wire N__40209;
    wire N__40206;
    wire N__40203;
    wire N__40200;
    wire N__40197;
    wire N__40192;
    wire N__40189;
    wire N__40186;
    wire N__40185;
    wire N__40182;
    wire N__40179;
    wire N__40174;
    wire N__40171;
    wire N__40168;
    wire N__40165;
    wire N__40162;
    wire N__40159;
    wire N__40156;
    wire N__40153;
    wire N__40150;
    wire N__40147;
    wire N__40144;
    wire N__40141;
    wire N__40138;
    wire N__40135;
    wire N__40132;
    wire N__40129;
    wire N__40126;
    wire N__40125;
    wire N__40122;
    wire N__40119;
    wire N__40116;
    wire N__40113;
    wire N__40110;
    wire N__40107;
    wire N__40104;
    wire N__40101;
    wire N__40098;
    wire N__40097;
    wire N__40094;
    wire N__40091;
    wire N__40088;
    wire N__40085;
    wire N__40082;
    wire N__40079;
    wire N__40074;
    wire N__40069;
    wire N__40066;
    wire N__40063;
    wire N__40060;
    wire N__40057;
    wire N__40054;
    wire N__40051;
    wire N__40048;
    wire N__40045;
    wire N__40042;
    wire N__40039;
    wire N__40036;
    wire N__40033;
    wire N__40030;
    wire N__40027;
    wire N__40024;
    wire N__40021;
    wire N__40020;
    wire N__40017;
    wire N__40014;
    wire N__40011;
    wire N__40008;
    wire N__40005;
    wire N__40002;
    wire N__39999;
    wire N__39996;
    wire N__39993;
    wire N__39990;
    wire N__39987;
    wire N__39986;
    wire N__39983;
    wire N__39980;
    wire N__39977;
    wire N__39972;
    wire N__39967;
    wire N__39964;
    wire N__39961;
    wire N__39958;
    wire N__39955;
    wire N__39952;
    wire N__39949;
    wire N__39946;
    wire N__39943;
    wire N__39940;
    wire N__39937;
    wire N__39934;
    wire N__39931;
    wire N__39928;
    wire N__39925;
    wire N__39922;
    wire N__39919;
    wire N__39916;
    wire N__39915;
    wire N__39912;
    wire N__39909;
    wire N__39906;
    wire N__39903;
    wire N__39900;
    wire N__39897;
    wire N__39894;
    wire N__39891;
    wire N__39888;
    wire N__39885;
    wire N__39882;
    wire N__39881;
    wire N__39878;
    wire N__39875;
    wire N__39872;
    wire N__39869;
    wire N__39866;
    wire N__39859;
    wire N__39856;
    wire N__39853;
    wire N__39850;
    wire N__39847;
    wire N__39844;
    wire N__39841;
    wire N__39838;
    wire N__39835;
    wire N__39832;
    wire N__39829;
    wire N__39826;
    wire N__39823;
    wire N__39820;
    wire N__39817;
    wire N__39814;
    wire N__39813;
    wire N__39810;
    wire N__39807;
    wire N__39804;
    wire N__39801;
    wire N__39798;
    wire N__39795;
    wire N__39792;
    wire N__39789;
    wire N__39786;
    wire N__39783;
    wire N__39780;
    wire N__39779;
    wire N__39776;
    wire N__39773;
    wire N__39770;
    wire N__39767;
    wire N__39764;
    wire N__39757;
    wire N__39754;
    wire N__39751;
    wire N__39748;
    wire N__39745;
    wire N__39742;
    wire N__39739;
    wire N__39736;
    wire N__39733;
    wire N__39730;
    wire N__39727;
    wire N__39724;
    wire N__39721;
    wire N__39718;
    wire N__39715;
    wire N__39712;
    wire N__39709;
    wire N__39706;
    wire N__39705;
    wire N__39702;
    wire N__39699;
    wire N__39696;
    wire N__39693;
    wire N__39690;
    wire N__39687;
    wire N__39684;
    wire N__39681;
    wire N__39678;
    wire N__39675;
    wire N__39672;
    wire N__39671;
    wire N__39668;
    wire N__39665;
    wire N__39662;
    wire N__39659;
    wire N__39656;
    wire N__39649;
    wire N__39646;
    wire N__39643;
    wire N__39640;
    wire N__39637;
    wire N__39634;
    wire N__39631;
    wire N__39628;
    wire N__39625;
    wire N__39622;
    wire N__39619;
    wire N__39616;
    wire N__39613;
    wire N__39610;
    wire N__39607;
    wire N__39604;
    wire N__39601;
    wire N__39598;
    wire N__39597;
    wire N__39594;
    wire N__39591;
    wire N__39588;
    wire N__39585;
    wire N__39582;
    wire N__39579;
    wire N__39576;
    wire N__39573;
    wire N__39570;
    wire N__39567;
    wire N__39564;
    wire N__39563;
    wire N__39560;
    wire N__39557;
    wire N__39554;
    wire N__39551;
    wire N__39548;
    wire N__39541;
    wire N__39538;
    wire N__39535;
    wire N__39532;
    wire N__39529;
    wire N__39526;
    wire N__39523;
    wire N__39520;
    wire N__39517;
    wire N__39514;
    wire N__39511;
    wire N__39508;
    wire N__39505;
    wire N__39502;
    wire N__39499;
    wire N__39496;
    wire N__39493;
    wire N__39492;
    wire N__39489;
    wire N__39486;
    wire N__39483;
    wire N__39480;
    wire N__39477;
    wire N__39474;
    wire N__39471;
    wire N__39468;
    wire N__39465;
    wire N__39462;
    wire N__39459;
    wire N__39458;
    wire N__39455;
    wire N__39452;
    wire N__39449;
    wire N__39446;
    wire N__39443;
    wire N__39436;
    wire N__39433;
    wire N__39430;
    wire N__39427;
    wire N__39424;
    wire N__39421;
    wire N__39418;
    wire N__39415;
    wire N__39412;
    wire N__39409;
    wire N__39406;
    wire N__39403;
    wire N__39400;
    wire N__39397;
    wire N__39394;
    wire N__39391;
    wire N__39390;
    wire N__39387;
    wire N__39384;
    wire N__39381;
    wire N__39378;
    wire N__39375;
    wire N__39372;
    wire N__39369;
    wire N__39366;
    wire N__39363;
    wire N__39360;
    wire N__39357;
    wire N__39356;
    wire N__39353;
    wire N__39350;
    wire N__39347;
    wire N__39344;
    wire N__39341;
    wire N__39334;
    wire N__39331;
    wire N__39330;
    wire N__39329;
    wire N__39328;
    wire N__39327;
    wire N__39324;
    wire N__39323;
    wire N__39318;
    wire N__39317;
    wire N__39316;
    wire N__39315;
    wire N__39314;
    wire N__39313;
    wire N__39308;
    wire N__39303;
    wire N__39300;
    wire N__39293;
    wire N__39288;
    wire N__39287;
    wire N__39286;
    wire N__39285;
    wire N__39280;
    wire N__39277;
    wire N__39274;
    wire N__39273;
    wire N__39272;
    wire N__39269;
    wire N__39262;
    wire N__39255;
    wire N__39250;
    wire N__39241;
    wire N__39240;
    wire N__39239;
    wire N__39238;
    wire N__39237;
    wire N__39236;
    wire N__39233;
    wire N__39226;
    wire N__39223;
    wire N__39220;
    wire N__39219;
    wire N__39212;
    wire N__39209;
    wire N__39206;
    wire N__39205;
    wire N__39198;
    wire N__39195;
    wire N__39190;
    wire N__39187;
    wire N__39184;
    wire N__39183;
    wire N__39180;
    wire N__39177;
    wire N__39174;
    wire N__39171;
    wire N__39168;
    wire N__39165;
    wire N__39160;
    wire N__39157;
    wire N__39156;
    wire N__39153;
    wire N__39152;
    wire N__39151;
    wire N__39150;
    wire N__39143;
    wire N__39142;
    wire N__39141;
    wire N__39138;
    wire N__39137;
    wire N__39134;
    wire N__39131;
    wire N__39128;
    wire N__39123;
    wire N__39122;
    wire N__39119;
    wire N__39116;
    wire N__39109;
    wire N__39108;
    wire N__39107;
    wire N__39106;
    wire N__39105;
    wire N__39102;
    wire N__39099;
    wire N__39094;
    wire N__39089;
    wire N__39086;
    wire N__39081;
    wire N__39076;
    wire N__39073;
    wire N__39064;
    wire N__39063;
    wire N__39058;
    wire N__39057;
    wire N__39054;
    wire N__39051;
    wire N__39048;
    wire N__39043;
    wire N__39040;
    wire N__39037;
    wire N__39034;
    wire N__39031;
    wire N__39028;
    wire N__39025;
    wire N__39022;
    wire N__39019;
    wire N__39016;
    wire N__39013;
    wire N__39010;
    wire N__39007;
    wire N__39004;
    wire N__39001;
    wire N__38998;
    wire N__38995;
    wire N__38992;
    wire N__38991;
    wire N__38988;
    wire N__38985;
    wire N__38982;
    wire N__38979;
    wire N__38976;
    wire N__38973;
    wire N__38970;
    wire N__38967;
    wire N__38964;
    wire N__38961;
    wire N__38958;
    wire N__38955;
    wire N__38952;
    wire N__38949;
    wire N__38946;
    wire N__38941;
    wire N__38938;
    wire N__38937;
    wire N__38936;
    wire N__38935;
    wire N__38932;
    wire N__38929;
    wire N__38926;
    wire N__38923;
    wire N__38920;
    wire N__38917;
    wire N__38914;
    wire N__38907;
    wire N__38902;
    wire N__38899;
    wire N__38898;
    wire N__38897;
    wire N__38894;
    wire N__38891;
    wire N__38888;
    wire N__38885;
    wire N__38882;
    wire N__38879;
    wire N__38874;
    wire N__38869;
    wire N__38866;
    wire N__38865;
    wire N__38862;
    wire N__38859;
    wire N__38856;
    wire N__38855;
    wire N__38852;
    wire N__38849;
    wire N__38846;
    wire N__38843;
    wire N__38838;
    wire N__38833;
    wire N__38830;
    wire N__38827;
    wire N__38826;
    wire N__38825;
    wire N__38822;
    wire N__38817;
    wire N__38812;
    wire N__38809;
    wire N__38808;
    wire N__38805;
    wire N__38802;
    wire N__38799;
    wire N__38794;
    wire N__38791;
    wire N__38790;
    wire N__38787;
    wire N__38784;
    wire N__38781;
    wire N__38776;
    wire N__38773;
    wire N__38770;
    wire N__38767;
    wire N__38764;
    wire N__38763;
    wire N__38760;
    wire N__38759;
    wire N__38756;
    wire N__38753;
    wire N__38750;
    wire N__38747;
    wire N__38744;
    wire N__38741;
    wire N__38734;
    wire N__38733;
    wire N__38732;
    wire N__38731;
    wire N__38730;
    wire N__38729;
    wire N__38726;
    wire N__38723;
    wire N__38720;
    wire N__38719;
    wire N__38716;
    wire N__38713;
    wire N__38712;
    wire N__38709;
    wire N__38706;
    wire N__38703;
    wire N__38700;
    wire N__38697;
    wire N__38694;
    wire N__38691;
    wire N__38688;
    wire N__38685;
    wire N__38682;
    wire N__38679;
    wire N__38676;
    wire N__38673;
    wire N__38668;
    wire N__38665;
    wire N__38662;
    wire N__38659;
    wire N__38654;
    wire N__38651;
    wire N__38650;
    wire N__38645;
    wire N__38640;
    wire N__38635;
    wire N__38632;
    wire N__38623;
    wire N__38620;
    wire N__38617;
    wire N__38614;
    wire N__38613;
    wire N__38612;
    wire N__38609;
    wire N__38606;
    wire N__38603;
    wire N__38600;
    wire N__38597;
    wire N__38590;
    wire N__38587;
    wire N__38584;
    wire N__38581;
    wire N__38580;
    wire N__38577;
    wire N__38574;
    wire N__38571;
    wire N__38568;
    wire N__38565;
    wire N__38562;
    wire N__38557;
    wire N__38554;
    wire N__38551;
    wire N__38550;
    wire N__38547;
    wire N__38546;
    wire N__38545;
    wire N__38544;
    wire N__38541;
    wire N__38540;
    wire N__38537;
    wire N__38534;
    wire N__38533;
    wire N__38530;
    wire N__38527;
    wire N__38524;
    wire N__38523;
    wire N__38520;
    wire N__38515;
    wire N__38512;
    wire N__38509;
    wire N__38504;
    wire N__38501;
    wire N__38498;
    wire N__38497;
    wire N__38494;
    wire N__38487;
    wire N__38482;
    wire N__38479;
    wire N__38470;
    wire N__38469;
    wire N__38466;
    wire N__38463;
    wire N__38460;
    wire N__38457;
    wire N__38454;
    wire N__38451;
    wire N__38446;
    wire N__38443;
    wire N__38442;
    wire N__38439;
    wire N__38436;
    wire N__38433;
    wire N__38430;
    wire N__38427;
    wire N__38422;
    wire N__38419;
    wire N__38418;
    wire N__38417;
    wire N__38414;
    wire N__38411;
    wire N__38408;
    wire N__38405;
    wire N__38402;
    wire N__38395;
    wire N__38394;
    wire N__38391;
    wire N__38390;
    wire N__38387;
    wire N__38384;
    wire N__38379;
    wire N__38374;
    wire N__38373;
    wire N__38372;
    wire N__38369;
    wire N__38364;
    wire N__38359;
    wire N__38356;
    wire N__38353;
    wire N__38350;
    wire N__38347;
    wire N__38346;
    wire N__38343;
    wire N__38340;
    wire N__38337;
    wire N__38334;
    wire N__38329;
    wire N__38326;
    wire N__38323;
    wire N__38320;
    wire N__38319;
    wire N__38316;
    wire N__38313;
    wire N__38308;
    wire N__38305;
    wire N__38304;
    wire N__38303;
    wire N__38300;
    wire N__38297;
    wire N__38294;
    wire N__38291;
    wire N__38288;
    wire N__38285;
    wire N__38282;
    wire N__38275;
    wire N__38272;
    wire N__38269;
    wire N__38266;
    wire N__38263;
    wire N__38260;
    wire N__38259;
    wire N__38256;
    wire N__38253;
    wire N__38250;
    wire N__38245;
    wire N__38242;
    wire N__38239;
    wire N__38236;
    wire N__38233;
    wire N__38230;
    wire N__38227;
    wire N__38224;
    wire N__38221;
    wire N__38218;
    wire N__38215;
    wire N__38212;
    wire N__38209;
    wire N__38208;
    wire N__38203;
    wire N__38202;
    wire N__38201;
    wire N__38198;
    wire N__38193;
    wire N__38190;
    wire N__38185;
    wire N__38182;
    wire N__38179;
    wire N__38176;
    wire N__38175;
    wire N__38172;
    wire N__38169;
    wire N__38166;
    wire N__38163;
    wire N__38162;
    wire N__38159;
    wire N__38156;
    wire N__38153;
    wire N__38148;
    wire N__38143;
    wire N__38140;
    wire N__38137;
    wire N__38134;
    wire N__38131;
    wire N__38128;
    wire N__38125;
    wire N__38122;
    wire N__38119;
    wire N__38116;
    wire N__38113;
    wire N__38110;
    wire N__38107;
    wire N__38104;
    wire N__38101;
    wire N__38098;
    wire N__38095;
    wire N__38092;
    wire N__38089;
    wire N__38086;
    wire N__38083;
    wire N__38080;
    wire N__38077;
    wire N__38076;
    wire N__38073;
    wire N__38070;
    wire N__38067;
    wire N__38064;
    wire N__38061;
    wire N__38056;
    wire N__38053;
    wire N__38050;
    wire N__38047;
    wire N__38044;
    wire N__38041;
    wire N__38038;
    wire N__38035;
    wire N__38032;
    wire N__38029;
    wire N__38026;
    wire N__38023;
    wire N__38022;
    wire N__38019;
    wire N__38018;
    wire N__38017;
    wire N__38016;
    wire N__38013;
    wire N__38010;
    wire N__38007;
    wire N__38004;
    wire N__38001;
    wire N__37996;
    wire N__37995;
    wire N__37994;
    wire N__37991;
    wire N__37988;
    wire N__37985;
    wire N__37982;
    wire N__37981;
    wire N__37978;
    wire N__37975;
    wire N__37972;
    wire N__37969;
    wire N__37966;
    wire N__37963;
    wire N__37960;
    wire N__37957;
    wire N__37954;
    wire N__37953;
    wire N__37948;
    wire N__37941;
    wire N__37938;
    wire N__37935;
    wire N__37932;
    wire N__37921;
    wire N__37920;
    wire N__37917;
    wire N__37914;
    wire N__37909;
    wire N__37906;
    wire N__37905;
    wire N__37902;
    wire N__37899;
    wire N__37894;
    wire N__37891;
    wire N__37888;
    wire N__37885;
    wire N__37884;
    wire N__37879;
    wire N__37878;
    wire N__37877;
    wire N__37876;
    wire N__37875;
    wire N__37874;
    wire N__37873;
    wire N__37872;
    wire N__37871;
    wire N__37870;
    wire N__37869;
    wire N__37868;
    wire N__37865;
    wire N__37860;
    wire N__37851;
    wire N__37848;
    wire N__37845;
    wire N__37844;
    wire N__37841;
    wire N__37840;
    wire N__37839;
    wire N__37838;
    wire N__37837;
    wire N__37836;
    wire N__37835;
    wire N__37834;
    wire N__37833;
    wire N__37832;
    wire N__37827;
    wire N__37824;
    wire N__37817;
    wire N__37814;
    wire N__37811;
    wire N__37808;
    wire N__37801;
    wire N__37788;
    wire N__37787;
    wire N__37786;
    wire N__37785;
    wire N__37784;
    wire N__37783;
    wire N__37782;
    wire N__37781;
    wire N__37780;
    wire N__37779;
    wire N__37776;
    wire N__37771;
    wire N__37766;
    wire N__37759;
    wire N__37752;
    wire N__37739;
    wire N__37726;
    wire N__37723;
    wire N__37720;
    wire N__37719;
    wire N__37718;
    wire N__37715;
    wire N__37712;
    wire N__37709;
    wire N__37702;
    wire N__37699;
    wire N__37696;
    wire N__37693;
    wire N__37690;
    wire N__37689;
    wire N__37686;
    wire N__37683;
    wire N__37678;
    wire N__37675;
    wire N__37672;
    wire N__37669;
    wire N__37666;
    wire N__37663;
    wire N__37662;
    wire N__37659;
    wire N__37656;
    wire N__37653;
    wire N__37650;
    wire N__37645;
    wire N__37642;
    wire N__37639;
    wire N__37636;
    wire N__37633;
    wire N__37630;
    wire N__37629;
    wire N__37628;
    wire N__37625;
    wire N__37620;
    wire N__37617;
    wire N__37614;
    wire N__37609;
    wire N__37606;
    wire N__37605;
    wire N__37604;
    wire N__37603;
    wire N__37602;
    wire N__37599;
    wire N__37596;
    wire N__37595;
    wire N__37594;
    wire N__37593;
    wire N__37590;
    wire N__37587;
    wire N__37584;
    wire N__37583;
    wire N__37582;
    wire N__37581;
    wire N__37580;
    wire N__37577;
    wire N__37574;
    wire N__37569;
    wire N__37566;
    wire N__37559;
    wire N__37550;
    wire N__37547;
    wire N__37540;
    wire N__37537;
    wire N__37528;
    wire N__37525;
    wire N__37522;
    wire N__37519;
    wire N__37516;
    wire N__37515;
    wire N__37512;
    wire N__37509;
    wire N__37506;
    wire N__37501;
    wire N__37498;
    wire N__37497;
    wire N__37494;
    wire N__37491;
    wire N__37488;
    wire N__37483;
    wire N__37482;
    wire N__37479;
    wire N__37476;
    wire N__37473;
    wire N__37470;
    wire N__37467;
    wire N__37464;
    wire N__37459;
    wire N__37456;
    wire N__37453;
    wire N__37452;
    wire N__37449;
    wire N__37446;
    wire N__37445;
    wire N__37444;
    wire N__37439;
    wire N__37436;
    wire N__37433;
    wire N__37426;
    wire N__37425;
    wire N__37424;
    wire N__37421;
    wire N__37418;
    wire N__37415;
    wire N__37412;
    wire N__37407;
    wire N__37404;
    wire N__37401;
    wire N__37396;
    wire N__37395;
    wire N__37392;
    wire N__37391;
    wire N__37388;
    wire N__37383;
    wire N__37378;
    wire N__37377;
    wire N__37376;
    wire N__37369;
    wire N__37366;
    wire N__37363;
    wire N__37360;
    wire N__37357;
    wire N__37356;
    wire N__37355;
    wire N__37350;
    wire N__37347;
    wire N__37346;
    wire N__37343;
    wire N__37342;
    wire N__37339;
    wire N__37336;
    wire N__37333;
    wire N__37330;
    wire N__37325;
    wire N__37322;
    wire N__37317;
    wire N__37314;
    wire N__37311;
    wire N__37308;
    wire N__37305;
    wire N__37300;
    wire N__37297;
    wire N__37294;
    wire N__37291;
    wire N__37288;
    wire N__37287;
    wire N__37284;
    wire N__37281;
    wire N__37278;
    wire N__37273;
    wire N__37270;
    wire N__37269;
    wire N__37266;
    wire N__37263;
    wire N__37258;
    wire N__37255;
    wire N__37252;
    wire N__37251;
    wire N__37248;
    wire N__37245;
    wire N__37240;
    wire N__37237;
    wire N__37236;
    wire N__37233;
    wire N__37230;
    wire N__37225;
    wire N__37222;
    wire N__37219;
    wire N__37218;
    wire N__37215;
    wire N__37212;
    wire N__37207;
    wire N__37204;
    wire N__37203;
    wire N__37200;
    wire N__37197;
    wire N__37192;
    wire N__37189;
    wire N__37186;
    wire N__37185;
    wire N__37182;
    wire N__37179;
    wire N__37174;
    wire N__37171;
    wire N__37170;
    wire N__37167;
    wire N__37164;
    wire N__37159;
    wire N__37156;
    wire N__37153;
    wire N__37150;
    wire N__37147;
    wire N__37144;
    wire N__37141;
    wire N__37138;
    wire N__37135;
    wire N__37132;
    wire N__37129;
    wire N__37126;
    wire N__37125;
    wire N__37122;
    wire N__37119;
    wire N__37114;
    wire N__37111;
    wire N__37110;
    wire N__37107;
    wire N__37104;
    wire N__37099;
    wire N__37096;
    wire N__37093;
    wire N__37092;
    wire N__37089;
    wire N__37086;
    wire N__37081;
    wire N__37078;
    wire N__37077;
    wire N__37074;
    wire N__37071;
    wire N__37066;
    wire N__37063;
    wire N__37062;
    wire N__37059;
    wire N__37056;
    wire N__37053;
    wire N__37050;
    wire N__37047;
    wire N__37042;
    wire N__37039;
    wire N__37038;
    wire N__37035;
    wire N__37032;
    wire N__37029;
    wire N__37024;
    wire N__37021;
    wire N__37018;
    wire N__37017;
    wire N__37014;
    wire N__37011;
    wire N__37006;
    wire N__37003;
    wire N__37000;
    wire N__36997;
    wire N__36994;
    wire N__36991;
    wire N__36988;
    wire N__36985;
    wire N__36982;
    wire N__36979;
    wire N__36978;
    wire N__36977;
    wire N__36974;
    wire N__36969;
    wire N__36964;
    wire N__36961;
    wire N__36958;
    wire N__36955;
    wire N__36952;
    wire N__36949;
    wire N__36948;
    wire N__36947;
    wire N__36944;
    wire N__36941;
    wire N__36938;
    wire N__36935;
    wire N__36932;
    wire N__36925;
    wire N__36922;
    wire N__36921;
    wire N__36920;
    wire N__36917;
    wire N__36914;
    wire N__36911;
    wire N__36908;
    wire N__36905;
    wire N__36898;
    wire N__36897;
    wire N__36896;
    wire N__36895;
    wire N__36894;
    wire N__36891;
    wire N__36888;
    wire N__36885;
    wire N__36882;
    wire N__36881;
    wire N__36880;
    wire N__36877;
    wire N__36874;
    wire N__36871;
    wire N__36868;
    wire N__36865;
    wire N__36862;
    wire N__36859;
    wire N__36858;
    wire N__36855;
    wire N__36850;
    wire N__36843;
    wire N__36840;
    wire N__36837;
    wire N__36834;
    wire N__36831;
    wire N__36826;
    wire N__36823;
    wire N__36814;
    wire N__36811;
    wire N__36808;
    wire N__36807;
    wire N__36804;
    wire N__36803;
    wire N__36800;
    wire N__36797;
    wire N__36796;
    wire N__36795;
    wire N__36792;
    wire N__36791;
    wire N__36790;
    wire N__36787;
    wire N__36784;
    wire N__36781;
    wire N__36780;
    wire N__36777;
    wire N__36774;
    wire N__36771;
    wire N__36768;
    wire N__36761;
    wire N__36758;
    wire N__36755;
    wire N__36752;
    wire N__36749;
    wire N__36742;
    wire N__36737;
    wire N__36734;
    wire N__36731;
    wire N__36724;
    wire N__36721;
    wire N__36718;
    wire N__36717;
    wire N__36714;
    wire N__36713;
    wire N__36710;
    wire N__36707;
    wire N__36704;
    wire N__36697;
    wire N__36694;
    wire N__36691;
    wire N__36688;
    wire N__36685;
    wire N__36682;
    wire N__36679;
    wire N__36678;
    wire N__36675;
    wire N__36672;
    wire N__36669;
    wire N__36664;
    wire N__36661;
    wire N__36658;
    wire N__36657;
    wire N__36654;
    wire N__36653;
    wire N__36650;
    wire N__36647;
    wire N__36644;
    wire N__36637;
    wire N__36636;
    wire N__36631;
    wire N__36628;
    wire N__36627;
    wire N__36624;
    wire N__36621;
    wire N__36618;
    wire N__36613;
    wire N__36612;
    wire N__36609;
    wire N__36606;
    wire N__36603;
    wire N__36598;
    wire N__36595;
    wire N__36592;
    wire N__36589;
    wire N__36588;
    wire N__36587;
    wire N__36584;
    wire N__36579;
    wire N__36574;
    wire N__36571;
    wire N__36568;
    wire N__36565;
    wire N__36564;
    wire N__36563;
    wire N__36560;
    wire N__36557;
    wire N__36554;
    wire N__36551;
    wire N__36548;
    wire N__36545;
    wire N__36538;
    wire N__36535;
    wire N__36532;
    wire N__36529;
    wire N__36526;
    wire N__36523;
    wire N__36520;
    wire N__36517;
    wire N__36514;
    wire N__36511;
    wire N__36508;
    wire N__36505;
    wire N__36502;
    wire N__36499;
    wire N__36496;
    wire N__36493;
    wire N__36490;
    wire N__36487;
    wire N__36484;
    wire N__36481;
    wire N__36478;
    wire N__36477;
    wire N__36474;
    wire N__36471;
    wire N__36468;
    wire N__36465;
    wire N__36462;
    wire N__36459;
    wire N__36456;
    wire N__36453;
    wire N__36450;
    wire N__36447;
    wire N__36444;
    wire N__36441;
    wire N__36438;
    wire N__36433;
    wire N__36430;
    wire N__36427;
    wire N__36426;
    wire N__36423;
    wire N__36420;
    wire N__36417;
    wire N__36412;
    wire N__36411;
    wire N__36408;
    wire N__36405;
    wire N__36402;
    wire N__36397;
    wire N__36396;
    wire N__36395;
    wire N__36394;
    wire N__36391;
    wire N__36388;
    wire N__36385;
    wire N__36382;
    wire N__36379;
    wire N__36378;
    wire N__36375;
    wire N__36370;
    wire N__36367;
    wire N__36364;
    wire N__36361;
    wire N__36358;
    wire N__36353;
    wire N__36346;
    wire N__36345;
    wire N__36340;
    wire N__36337;
    wire N__36334;
    wire N__36333;
    wire N__36330;
    wire N__36327;
    wire N__36324;
    wire N__36319;
    wire N__36318;
    wire N__36315;
    wire N__36312;
    wire N__36309;
    wire N__36304;
    wire N__36303;
    wire N__36302;
    wire N__36299;
    wire N__36296;
    wire N__36293;
    wire N__36290;
    wire N__36287;
    wire N__36280;
    wire N__36277;
    wire N__36274;
    wire N__36271;
    wire N__36268;
    wire N__36265;
    wire N__36262;
    wire N__36259;
    wire N__36256;
    wire N__36255;
    wire N__36254;
    wire N__36253;
    wire N__36252;
    wire N__36249;
    wire N__36246;
    wire N__36243;
    wire N__36242;
    wire N__36241;
    wire N__36238;
    wire N__36237;
    wire N__36234;
    wire N__36233;
    wire N__36228;
    wire N__36225;
    wire N__36222;
    wire N__36219;
    wire N__36216;
    wire N__36213;
    wire N__36210;
    wire N__36207;
    wire N__36204;
    wire N__36199;
    wire N__36188;
    wire N__36185;
    wire N__36182;
    wire N__36179;
    wire N__36176;
    wire N__36171;
    wire N__36166;
    wire N__36165;
    wire N__36164;
    wire N__36161;
    wire N__36154;
    wire N__36151;
    wire N__36148;
    wire N__36145;
    wire N__36144;
    wire N__36143;
    wire N__36140;
    wire N__36137;
    wire N__36134;
    wire N__36131;
    wire N__36124;
    wire N__36121;
    wire N__36118;
    wire N__36115;
    wire N__36112;
    wire N__36109;
    wire N__36108;
    wire N__36105;
    wire N__36104;
    wire N__36101;
    wire N__36098;
    wire N__36095;
    wire N__36088;
    wire N__36085;
    wire N__36082;
    wire N__36079;
    wire N__36076;
    wire N__36073;
    wire N__36070;
    wire N__36067;
    wire N__36064;
    wire N__36061;
    wire N__36058;
    wire N__36055;
    wire N__36052;
    wire N__36049;
    wire N__36046;
    wire N__36043;
    wire N__36040;
    wire N__36039;
    wire N__36036;
    wire N__36033;
    wire N__36030;
    wire N__36025;
    wire N__36022;
    wire N__36019;
    wire N__36016;
    wire N__36013;
    wire N__36010;
    wire N__36007;
    wire N__36004;
    wire N__36001;
    wire N__35998;
    wire N__35995;
    wire N__35992;
    wire N__35991;
    wire N__35988;
    wire N__35985;
    wire N__35982;
    wire N__35979;
    wire N__35978;
    wire N__35977;
    wire N__35972;
    wire N__35971;
    wire N__35968;
    wire N__35967;
    wire N__35964;
    wire N__35961;
    wire N__35958;
    wire N__35955;
    wire N__35952;
    wire N__35951;
    wire N__35948;
    wire N__35943;
    wire N__35938;
    wire N__35935;
    wire N__35934;
    wire N__35933;
    wire N__35930;
    wire N__35927;
    wire N__35922;
    wire N__35919;
    wire N__35916;
    wire N__35905;
    wire N__35902;
    wire N__35899;
    wire N__35896;
    wire N__35895;
    wire N__35892;
    wire N__35889;
    wire N__35886;
    wire N__35881;
    wire N__35878;
    wire N__35875;
    wire N__35872;
    wire N__35869;
    wire N__35866;
    wire N__35863;
    wire N__35860;
    wire N__35857;
    wire N__35856;
    wire N__35855;
    wire N__35852;
    wire N__35849;
    wire N__35846;
    wire N__35843;
    wire N__35838;
    wire N__35833;
    wire N__35830;
    wire N__35827;
    wire N__35824;
    wire N__35821;
    wire N__35818;
    wire N__35815;
    wire N__35812;
    wire N__35811;
    wire N__35810;
    wire N__35807;
    wire N__35806;
    wire N__35803;
    wire N__35802;
    wire N__35799;
    wire N__35798;
    wire N__35795;
    wire N__35792;
    wire N__35789;
    wire N__35786;
    wire N__35783;
    wire N__35780;
    wire N__35779;
    wire N__35776;
    wire N__35773;
    wire N__35770;
    wire N__35767;
    wire N__35762;
    wire N__35759;
    wire N__35758;
    wire N__35757;
    wire N__35754;
    wire N__35751;
    wire N__35748;
    wire N__35745;
    wire N__35742;
    wire N__35739;
    wire N__35736;
    wire N__35733;
    wire N__35716;
    wire N__35713;
    wire N__35710;
    wire N__35707;
    wire N__35704;
    wire N__35701;
    wire N__35698;
    wire N__35695;
    wire N__35692;
    wire N__35689;
    wire N__35686;
    wire N__35683;
    wire N__35680;
    wire N__35677;
    wire N__35674;
    wire N__35671;
    wire N__35668;
    wire N__35665;
    wire N__35664;
    wire N__35663;
    wire N__35662;
    wire N__35661;
    wire N__35658;
    wire N__35655;
    wire N__35652;
    wire N__35649;
    wire N__35646;
    wire N__35641;
    wire N__35640;
    wire N__35637;
    wire N__35636;
    wire N__35633;
    wire N__35628;
    wire N__35625;
    wire N__35622;
    wire N__35619;
    wire N__35618;
    wire N__35617;
    wire N__35614;
    wire N__35611;
    wire N__35608;
    wire N__35603;
    wire N__35600;
    wire N__35597;
    wire N__35584;
    wire N__35581;
    wire N__35578;
    wire N__35575;
    wire N__35572;
    wire N__35569;
    wire N__35568;
    wire N__35567;
    wire N__35564;
    wire N__35563;
    wire N__35560;
    wire N__35559;
    wire N__35558;
    wire N__35555;
    wire N__35552;
    wire N__35549;
    wire N__35546;
    wire N__35543;
    wire N__35540;
    wire N__35537;
    wire N__35534;
    wire N__35531;
    wire N__35530;
    wire N__35525;
    wire N__35522;
    wire N__35519;
    wire N__35514;
    wire N__35511;
    wire N__35510;
    wire N__35509;
    wire N__35502;
    wire N__35497;
    wire N__35494;
    wire N__35491;
    wire N__35482;
    wire N__35479;
    wire N__35476;
    wire N__35473;
    wire N__35470;
    wire N__35467;
    wire N__35464;
    wire N__35461;
    wire N__35458;
    wire N__35455;
    wire N__35452;
    wire N__35451;
    wire N__35450;
    wire N__35449;
    wire N__35448;
    wire N__35445;
    wire N__35442;
    wire N__35441;
    wire N__35438;
    wire N__35433;
    wire N__35428;
    wire N__35425;
    wire N__35422;
    wire N__35421;
    wire N__35420;
    wire N__35417;
    wire N__35414;
    wire N__35411;
    wire N__35408;
    wire N__35405;
    wire N__35402;
    wire N__35401;
    wire N__35398;
    wire N__35395;
    wire N__35392;
    wire N__35387;
    wire N__35384;
    wire N__35381;
    wire N__35368;
    wire N__35365;
    wire N__35362;
    wire N__35359;
    wire N__35356;
    wire N__35353;
    wire N__35350;
    wire N__35347;
    wire N__35344;
    wire N__35341;
    wire N__35338;
    wire N__35335;
    wire N__35332;
    wire N__35329;
    wire N__35326;
    wire N__35325;
    wire N__35322;
    wire N__35319;
    wire N__35316;
    wire N__35313;
    wire N__35308;
    wire N__35305;
    wire N__35302;
    wire N__35301;
    wire N__35298;
    wire N__35295;
    wire N__35292;
    wire N__35289;
    wire N__35284;
    wire N__35283;
    wire N__35280;
    wire N__35277;
    wire N__35276;
    wire N__35273;
    wire N__35270;
    wire N__35267;
    wire N__35264;
    wire N__35261;
    wire N__35258;
    wire N__35255;
    wire N__35252;
    wire N__35245;
    wire N__35242;
    wire N__35239;
    wire N__35236;
    wire N__35233;
    wire N__35230;
    wire N__35227;
    wire N__35224;
    wire N__35221;
    wire N__35218;
    wire N__35215;
    wire N__35212;
    wire N__35209;
    wire N__35206;
    wire N__35203;
    wire N__35200;
    wire N__35197;
    wire N__35194;
    wire N__35191;
    wire N__35188;
    wire N__35185;
    wire N__35182;
    wire N__35179;
    wire N__35176;
    wire N__35173;
    wire N__35170;
    wire N__35167;
    wire N__35164;
    wire N__35161;
    wire N__35158;
    wire N__35155;
    wire N__35152;
    wire N__35149;
    wire N__35146;
    wire N__35143;
    wire N__35140;
    wire N__35137;
    wire N__35134;
    wire N__35131;
    wire N__35128;
    wire N__35125;
    wire N__35122;
    wire N__35119;
    wire N__35116;
    wire N__35113;
    wire N__35110;
    wire N__35107;
    wire N__35104;
    wire N__35101;
    wire N__35098;
    wire N__35095;
    wire N__35092;
    wire N__35089;
    wire N__35086;
    wire N__35083;
    wire N__35082;
    wire N__35079;
    wire N__35076;
    wire N__35073;
    wire N__35070;
    wire N__35067;
    wire N__35062;
    wire N__35059;
    wire N__35056;
    wire N__35053;
    wire N__35050;
    wire N__35047;
    wire N__35044;
    wire N__35041;
    wire N__35038;
    wire N__35035;
    wire N__35032;
    wire N__35029;
    wire N__35026;
    wire N__35023;
    wire N__35020;
    wire N__35017;
    wire N__35014;
    wire N__35011;
    wire N__35008;
    wire N__35005;
    wire N__35002;
    wire N__34999;
    wire N__34996;
    wire N__34995;
    wire N__34994;
    wire N__34991;
    wire N__34988;
    wire N__34985;
    wire N__34980;
    wire N__34975;
    wire N__34974;
    wire N__34971;
    wire N__34970;
    wire N__34967;
    wire N__34964;
    wire N__34963;
    wire N__34962;
    wire N__34959;
    wire N__34956;
    wire N__34953;
    wire N__34950;
    wire N__34947;
    wire N__34936;
    wire N__34935;
    wire N__34932;
    wire N__34931;
    wire N__34930;
    wire N__34927;
    wire N__34922;
    wire N__34919;
    wire N__34918;
    wire N__34915;
    wire N__34914;
    wire N__34913;
    wire N__34908;
    wire N__34905;
    wire N__34902;
    wire N__34897;
    wire N__34894;
    wire N__34885;
    wire N__34882;
    wire N__34879;
    wire N__34878;
    wire N__34877;
    wire N__34876;
    wire N__34873;
    wire N__34872;
    wire N__34869;
    wire N__34866;
    wire N__34865;
    wire N__34864;
    wire N__34861;
    wire N__34858;
    wire N__34855;
    wire N__34850;
    wire N__34847;
    wire N__34846;
    wire N__34845;
    wire N__34844;
    wire N__34841;
    wire N__34838;
    wire N__34835;
    wire N__34832;
    wire N__34827;
    wire N__34820;
    wire N__34817;
    wire N__34812;
    wire N__34805;
    wire N__34802;
    wire N__34799;
    wire N__34796;
    wire N__34793;
    wire N__34790;
    wire N__34787;
    wire N__34784;
    wire N__34779;
    wire N__34774;
    wire N__34773;
    wire N__34772;
    wire N__34771;
    wire N__34770;
    wire N__34769;
    wire N__34768;
    wire N__34765;
    wire N__34762;
    wire N__34755;
    wire N__34752;
    wire N__34751;
    wire N__34748;
    wire N__34747;
    wire N__34746;
    wire N__34745;
    wire N__34744;
    wire N__34743;
    wire N__34742;
    wire N__34741;
    wire N__34740;
    wire N__34739;
    wire N__34736;
    wire N__34731;
    wire N__34728;
    wire N__34725;
    wire N__34724;
    wire N__34723;
    wire N__34720;
    wire N__34717;
    wire N__34716;
    wire N__34713;
    wire N__34712;
    wire N__34709;
    wire N__34704;
    wire N__34701;
    wire N__34698;
    wire N__34693;
    wire N__34686;
    wire N__34679;
    wire N__34674;
    wire N__34667;
    wire N__34648;
    wire N__34645;
    wire N__34642;
    wire N__34641;
    wire N__34640;
    wire N__34639;
    wire N__34638;
    wire N__34637;
    wire N__34636;
    wire N__34635;
    wire N__34634;
    wire N__34633;
    wire N__34632;
    wire N__34631;
    wire N__34630;
    wire N__34629;
    wire N__34628;
    wire N__34627;
    wire N__34626;
    wire N__34625;
    wire N__34624;
    wire N__34621;
    wire N__34620;
    wire N__34617;
    wire N__34602;
    wire N__34595;
    wire N__34594;
    wire N__34593;
    wire N__34590;
    wire N__34589;
    wire N__34588;
    wire N__34585;
    wire N__34584;
    wire N__34575;
    wire N__34574;
    wire N__34573;
    wire N__34572;
    wire N__34571;
    wire N__34570;
    wire N__34569;
    wire N__34568;
    wire N__34567;
    wire N__34566;
    wire N__34565;
    wire N__34564;
    wire N__34563;
    wire N__34562;
    wire N__34561;
    wire N__34556;
    wire N__34553;
    wire N__34546;
    wire N__34541;
    wire N__34536;
    wire N__34533;
    wire N__34530;
    wire N__34527;
    wire N__34524;
    wire N__34507;
    wire N__34504;
    wire N__34503;
    wire N__34500;
    wire N__34497;
    wire N__34494;
    wire N__34491;
    wire N__34490;
    wire N__34489;
    wire N__34488;
    wire N__34487;
    wire N__34486;
    wire N__34485;
    wire N__34482;
    wire N__34479;
    wire N__34476;
    wire N__34467;
    wire N__34466;
    wire N__34465;
    wire N__34456;
    wire N__34453;
    wire N__34446;
    wire N__34443;
    wire N__34436;
    wire N__34425;
    wire N__34418;
    wire N__34413;
    wire N__34406;
    wire N__34393;
    wire N__34390;
    wire N__34387;
    wire N__34386;
    wire N__34385;
    wire N__34384;
    wire N__34381;
    wire N__34376;
    wire N__34375;
    wire N__34374;
    wire N__34373;
    wire N__34372;
    wire N__34371;
    wire N__34370;
    wire N__34369;
    wire N__34368;
    wire N__34367;
    wire N__34366;
    wire N__34365;
    wire N__34364;
    wire N__34363;
    wire N__34362;
    wire N__34361;
    wire N__34360;
    wire N__34357;
    wire N__34356;
    wire N__34355;
    wire N__34350;
    wire N__34347;
    wire N__34336;
    wire N__34333;
    wire N__34330;
    wire N__34317;
    wire N__34314;
    wire N__34311;
    wire N__34308;
    wire N__34307;
    wire N__34306;
    wire N__34305;
    wire N__34304;
    wire N__34303;
    wire N__34302;
    wire N__34301;
    wire N__34300;
    wire N__34299;
    wire N__34296;
    wire N__34295;
    wire N__34294;
    wire N__34293;
    wire N__34292;
    wire N__34291;
    wire N__34290;
    wire N__34289;
    wire N__34286;
    wire N__34281;
    wire N__34276;
    wire N__34273;
    wire N__34268;
    wire N__34263;
    wire N__34262;
    wire N__34261;
    wire N__34260;
    wire N__34259;
    wire N__34258;
    wire N__34257;
    wire N__34256;
    wire N__34255;
    wire N__34252;
    wire N__34239;
    wire N__34236;
    wire N__34233;
    wire N__34224;
    wire N__34215;
    wire N__34210;
    wire N__34201;
    wire N__34184;
    wire N__34181;
    wire N__34162;
    wire N__34159;
    wire N__34158;
    wire N__34157;
    wire N__34156;
    wire N__34155;
    wire N__34154;
    wire N__34153;
    wire N__34152;
    wire N__34151;
    wire N__34150;
    wire N__34149;
    wire N__34148;
    wire N__34147;
    wire N__34142;
    wire N__34141;
    wire N__34136;
    wire N__34133;
    wire N__34128;
    wire N__34123;
    wire N__34122;
    wire N__34121;
    wire N__34120;
    wire N__34115;
    wire N__34114;
    wire N__34113;
    wire N__34112;
    wire N__34109;
    wire N__34106;
    wire N__34103;
    wire N__34100;
    wire N__34097;
    wire N__34096;
    wire N__34095;
    wire N__34094;
    wire N__34089;
    wire N__34086;
    wire N__34083;
    wire N__34080;
    wire N__34077;
    wire N__34074;
    wire N__34071;
    wire N__34066;
    wire N__34063;
    wire N__34060;
    wire N__34057;
    wire N__34052;
    wire N__34045;
    wire N__34042;
    wire N__34037;
    wire N__34012;
    wire N__34009;
    wire N__34006;
    wire N__34003;
    wire N__34000;
    wire N__33997;
    wire N__33994;
    wire N__33991;
    wire N__33988;
    wire N__33985;
    wire N__33982;
    wire N__33979;
    wire N__33976;
    wire N__33973;
    wire N__33970;
    wire N__33967;
    wire N__33964;
    wire N__33961;
    wire N__33960;
    wire N__33957;
    wire N__33954;
    wire N__33951;
    wire N__33948;
    wire N__33945;
    wire N__33940;
    wire N__33937;
    wire N__33936;
    wire N__33933;
    wire N__33930;
    wire N__33927;
    wire N__33924;
    wire N__33923;
    wire N__33918;
    wire N__33915;
    wire N__33914;
    wire N__33911;
    wire N__33908;
    wire N__33905;
    wire N__33898;
    wire N__33895;
    wire N__33894;
    wire N__33891;
    wire N__33888;
    wire N__33885;
    wire N__33882;
    wire N__33877;
    wire N__33874;
    wire N__33871;
    wire N__33868;
    wire N__33865;
    wire N__33864;
    wire N__33861;
    wire N__33858;
    wire N__33857;
    wire N__33854;
    wire N__33851;
    wire N__33848;
    wire N__33843;
    wire N__33838;
    wire N__33835;
    wire N__33832;
    wire N__33829;
    wire N__33826;
    wire N__33823;
    wire N__33820;
    wire N__33819;
    wire N__33818;
    wire N__33815;
    wire N__33812;
    wire N__33809;
    wire N__33802;
    wire N__33799;
    wire N__33796;
    wire N__33793;
    wire N__33790;
    wire N__33787;
    wire N__33784;
    wire N__33781;
    wire N__33780;
    wire N__33777;
    wire N__33774;
    wire N__33769;
    wire N__33766;
    wire N__33763;
    wire N__33760;
    wire N__33757;
    wire N__33754;
    wire N__33753;
    wire N__33750;
    wire N__33747;
    wire N__33744;
    wire N__33739;
    wire N__33736;
    wire N__33733;
    wire N__33730;
    wire N__33729;
    wire N__33726;
    wire N__33723;
    wire N__33720;
    wire N__33715;
    wire N__33712;
    wire N__33709;
    wire N__33706;
    wire N__33703;
    wire N__33700;
    wire N__33697;
    wire N__33696;
    wire N__33693;
    wire N__33690;
    wire N__33687;
    wire N__33682;
    wire N__33679;
    wire N__33676;
    wire N__33675;
    wire N__33672;
    wire N__33669;
    wire N__33666;
    wire N__33661;
    wire N__33658;
    wire N__33655;
    wire N__33654;
    wire N__33651;
    wire N__33648;
    wire N__33645;
    wire N__33640;
    wire N__33637;
    wire N__33634;
    wire N__33631;
    wire N__33630;
    wire N__33627;
    wire N__33624;
    wire N__33621;
    wire N__33616;
    wire N__33613;
    wire N__33610;
    wire N__33607;
    wire N__33606;
    wire N__33603;
    wire N__33600;
    wire N__33597;
    wire N__33592;
    wire N__33589;
    wire N__33586;
    wire N__33583;
    wire N__33580;
    wire N__33577;
    wire N__33574;
    wire N__33571;
    wire N__33568;
    wire N__33565;
    wire N__33562;
    wire N__33559;
    wire N__33558;
    wire N__33555;
    wire N__33552;
    wire N__33549;
    wire N__33546;
    wire N__33541;
    wire N__33538;
    wire N__33535;
    wire N__33534;
    wire N__33533;
    wire N__33530;
    wire N__33527;
    wire N__33524;
    wire N__33521;
    wire N__33514;
    wire N__33511;
    wire N__33508;
    wire N__33505;
    wire N__33502;
    wire N__33499;
    wire N__33496;
    wire N__33493;
    wire N__33492;
    wire N__33489;
    wire N__33486;
    wire N__33481;
    wire N__33478;
    wire N__33475;
    wire N__33472;
    wire N__33469;
    wire N__33466;
    wire N__33463;
    wire N__33462;
    wire N__33461;
    wire N__33458;
    wire N__33455;
    wire N__33452;
    wire N__33449;
    wire N__33442;
    wire N__33439;
    wire N__33438;
    wire N__33435;
    wire N__33432;
    wire N__33429;
    wire N__33426;
    wire N__33421;
    wire N__33418;
    wire N__33415;
    wire N__33412;
    wire N__33409;
    wire N__33406;
    wire N__33403;
    wire N__33400;
    wire N__33397;
    wire N__33394;
    wire N__33391;
    wire N__33390;
    wire N__33387;
    wire N__33384;
    wire N__33381;
    wire N__33376;
    wire N__33373;
    wire N__33370;
    wire N__33367;
    wire N__33364;
    wire N__33361;
    wire N__33358;
    wire N__33355;
    wire N__33354;
    wire N__33353;
    wire N__33350;
    wire N__33345;
    wire N__33340;
    wire N__33337;
    wire N__33336;
    wire N__33333;
    wire N__33330;
    wire N__33325;
    wire N__33322;
    wire N__33319;
    wire N__33316;
    wire N__33313;
    wire N__33310;
    wire N__33307;
    wire N__33304;
    wire N__33301;
    wire N__33298;
    wire N__33295;
    wire N__33292;
    wire N__33289;
    wire N__33286;
    wire N__33283;
    wire N__33280;
    wire N__33277;
    wire N__33274;
    wire N__33271;
    wire N__33268;
    wire N__33265;
    wire N__33262;
    wire N__33261;
    wire N__33258;
    wire N__33255;
    wire N__33252;
    wire N__33249;
    wire N__33244;
    wire N__33241;
    wire N__33238;
    wire N__33235;
    wire N__33232;
    wire N__33229;
    wire N__33226;
    wire N__33223;
    wire N__33220;
    wire N__33217;
    wire N__33214;
    wire N__33211;
    wire N__33208;
    wire N__33207;
    wire N__33204;
    wire N__33201;
    wire N__33198;
    wire N__33195;
    wire N__33190;
    wire N__33187;
    wire N__33184;
    wire N__33181;
    wire N__33178;
    wire N__33175;
    wire N__33172;
    wire N__33169;
    wire N__33166;
    wire N__33163;
    wire N__33162;
    wire N__33159;
    wire N__33156;
    wire N__33151;
    wire N__33148;
    wire N__33145;
    wire N__33142;
    wire N__33139;
    wire N__33136;
    wire N__33133;
    wire N__33130;
    wire N__33127;
    wire N__33124;
    wire N__33121;
    wire N__33118;
    wire N__33115;
    wire N__33112;
    wire N__33109;
    wire N__33106;
    wire N__33103;
    wire N__33100;
    wire N__33097;
    wire N__33094;
    wire N__33091;
    wire N__33088;
    wire N__33085;
    wire N__33082;
    wire N__33079;
    wire N__33076;
    wire N__33075;
    wire N__33072;
    wire N__33069;
    wire N__33066;
    wire N__33061;
    wire N__33058;
    wire N__33055;
    wire N__33052;
    wire N__33049;
    wire N__33046;
    wire N__33043;
    wire N__33040;
    wire N__33037;
    wire N__33034;
    wire N__33033;
    wire N__33032;
    wire N__33031;
    wire N__33024;
    wire N__33021;
    wire N__33016;
    wire N__33015;
    wire N__33012;
    wire N__33011;
    wire N__33010;
    wire N__33009;
    wire N__33006;
    wire N__32997;
    wire N__32994;
    wire N__32989;
    wire N__32988;
    wire N__32987;
    wire N__32984;
    wire N__32979;
    wire N__32976;
    wire N__32971;
    wire N__32968;
    wire N__32965;
    wire N__32962;
    wire N__32959;
    wire N__32956;
    wire N__32953;
    wire N__32952;
    wire N__32951;
    wire N__32948;
    wire N__32943;
    wire N__32938;
    wire N__32935;
    wire N__32932;
    wire N__32931;
    wire N__32930;
    wire N__32927;
    wire N__32924;
    wire N__32921;
    wire N__32914;
    wire N__32913;
    wire N__32912;
    wire N__32909;
    wire N__32908;
    wire N__32905;
    wire N__32904;
    wire N__32903;
    wire N__32900;
    wire N__32897;
    wire N__32896;
    wire N__32895;
    wire N__32894;
    wire N__32893;
    wire N__32890;
    wire N__32887;
    wire N__32886;
    wire N__32885;
    wire N__32884;
    wire N__32881;
    wire N__32880;
    wire N__32877;
    wire N__32874;
    wire N__32873;
    wire N__32872;
    wire N__32871;
    wire N__32868;
    wire N__32865;
    wire N__32862;
    wire N__32861;
    wire N__32858;
    wire N__32855;
    wire N__32850;
    wire N__32847;
    wire N__32846;
    wire N__32843;
    wire N__32842;
    wire N__32839;
    wire N__32836;
    wire N__32833;
    wire N__32830;
    wire N__32827;
    wire N__32824;
    wire N__32821;
    wire N__32818;
    wire N__32815;
    wire N__32810;
    wire N__32807;
    wire N__32806;
    wire N__32801;
    wire N__32796;
    wire N__32793;
    wire N__32790;
    wire N__32787;
    wire N__32784;
    wire N__32779;
    wire N__32778;
    wire N__32775;
    wire N__32770;
    wire N__32765;
    wire N__32762;
    wire N__32757;
    wire N__32754;
    wire N__32751;
    wire N__32746;
    wire N__32741;
    wire N__32736;
    wire N__32733;
    wire N__32728;
    wire N__32727;
    wire N__32724;
    wire N__32719;
    wire N__32716;
    wire N__32711;
    wire N__32704;
    wire N__32701;
    wire N__32698;
    wire N__32693;
    wire N__32688;
    wire N__32685;
    wire N__32680;
    wire N__32671;
    wire N__32668;
    wire N__32665;
    wire N__32662;
    wire N__32659;
    wire N__32656;
    wire N__32653;
    wire N__32650;
    wire N__32647;
    wire N__32644;
    wire N__32641;
    wire N__32640;
    wire N__32637;
    wire N__32634;
    wire N__32633;
    wire N__32632;
    wire N__32629;
    wire N__32626;
    wire N__32625;
    wire N__32622;
    wire N__32619;
    wire N__32616;
    wire N__32613;
    wire N__32610;
    wire N__32599;
    wire N__32596;
    wire N__32595;
    wire N__32592;
    wire N__32591;
    wire N__32590;
    wire N__32589;
    wire N__32586;
    wire N__32583;
    wire N__32580;
    wire N__32575;
    wire N__32566;
    wire N__32563;
    wire N__32560;
    wire N__32557;
    wire N__32554;
    wire N__32551;
    wire N__32548;
    wire N__32547;
    wire N__32546;
    wire N__32543;
    wire N__32542;
    wire N__32541;
    wire N__32538;
    wire N__32535;
    wire N__32532;
    wire N__32527;
    wire N__32518;
    wire N__32515;
    wire N__32512;
    wire N__32511;
    wire N__32510;
    wire N__32509;
    wire N__32506;
    wire N__32505;
    wire N__32502;
    wire N__32499;
    wire N__32496;
    wire N__32493;
    wire N__32488;
    wire N__32479;
    wire N__32476;
    wire N__32473;
    wire N__32470;
    wire N__32467;
    wire N__32466;
    wire N__32465;
    wire N__32464;
    wire N__32463;
    wire N__32460;
    wire N__32457;
    wire N__32450;
    wire N__32447;
    wire N__32440;
    wire N__32437;
    wire N__32436;
    wire N__32435;
    wire N__32432;
    wire N__32429;
    wire N__32426;
    wire N__32419;
    wire N__32416;
    wire N__32413;
    wire N__32410;
    wire N__32409;
    wire N__32404;
    wire N__32401;
    wire N__32398;
    wire N__32395;
    wire N__32392;
    wire N__32389;
    wire N__32386;
    wire N__32383;
    wire N__32382;
    wire N__32379;
    wire N__32376;
    wire N__32371;
    wire N__32370;
    wire N__32367;
    wire N__32366;
    wire N__32363;
    wire N__32360;
    wire N__32355;
    wire N__32350;
    wire N__32347;
    wire N__32344;
    wire N__32341;
    wire N__32338;
    wire N__32337;
    wire N__32336;
    wire N__32333;
    wire N__32330;
    wire N__32327;
    wire N__32320;
    wire N__32317;
    wire N__32314;
    wire N__32311;
    wire N__32310;
    wire N__32307;
    wire N__32304;
    wire N__32301;
    wire N__32300;
    wire N__32297;
    wire N__32294;
    wire N__32291;
    wire N__32288;
    wire N__32281;
    wire N__32278;
    wire N__32275;
    wire N__32272;
    wire N__32271;
    wire N__32268;
    wire N__32265;
    wire N__32262;
    wire N__32259;
    wire N__32258;
    wire N__32255;
    wire N__32252;
    wire N__32249;
    wire N__32246;
    wire N__32239;
    wire N__32238;
    wire N__32235;
    wire N__32232;
    wire N__32231;
    wire N__32228;
    wire N__32225;
    wire N__32222;
    wire N__32219;
    wire N__32212;
    wire N__32209;
    wire N__32206;
    wire N__32203;
    wire N__32200;
    wire N__32197;
    wire N__32194;
    wire N__32191;
    wire N__32188;
    wire N__32185;
    wire N__32182;
    wire N__32181;
    wire N__32180;
    wire N__32179;
    wire N__32178;
    wire N__32173;
    wire N__32170;
    wire N__32165;
    wire N__32164;
    wire N__32163;
    wire N__32162;
    wire N__32161;
    wire N__32160;
    wire N__32159;
    wire N__32158;
    wire N__32157;
    wire N__32156;
    wire N__32155;
    wire N__32152;
    wire N__32147;
    wire N__32138;
    wire N__32131;
    wire N__32128;
    wire N__32125;
    wire N__32122;
    wire N__32117;
    wire N__32108;
    wire N__32101;
    wire N__32100;
    wire N__32099;
    wire N__32096;
    wire N__32095;
    wire N__32094;
    wire N__32091;
    wire N__32088;
    wire N__32087;
    wire N__32084;
    wire N__32079;
    wire N__32074;
    wire N__32071;
    wire N__32070;
    wire N__32069;
    wire N__32068;
    wire N__32067;
    wire N__32064;
    wire N__32061;
    wire N__32058;
    wire N__32055;
    wire N__32052;
    wire N__32045;
    wire N__32032;
    wire N__32029;
    wire N__32026;
    wire N__32023;
    wire N__32020;
    wire N__32017;
    wire N__32016;
    wire N__32013;
    wire N__32012;
    wire N__32009;
    wire N__32006;
    wire N__32003;
    wire N__31998;
    wire N__31995;
    wire N__31990;
    wire N__31987;
    wire N__31986;
    wire N__31983;
    wire N__31980;
    wire N__31979;
    wire N__31976;
    wire N__31973;
    wire N__31970;
    wire N__31965;
    wire N__31960;
    wire N__31957;
    wire N__31954;
    wire N__31951;
    wire N__31948;
    wire N__31945;
    wire N__31942;
    wire N__31939;
    wire N__31936;
    wire N__31933;
    wire N__31932;
    wire N__31931;
    wire N__31928;
    wire N__31925;
    wire N__31922;
    wire N__31917;
    wire N__31914;
    wire N__31911;
    wire N__31906;
    wire N__31905;
    wire N__31904;
    wire N__31899;
    wire N__31896;
    wire N__31891;
    wire N__31888;
    wire N__31885;
    wire N__31884;
    wire N__31883;
    wire N__31882;
    wire N__31879;
    wire N__31876;
    wire N__31873;
    wire N__31870;
    wire N__31861;
    wire N__31860;
    wire N__31859;
    wire N__31858;
    wire N__31855;
    wire N__31852;
    wire N__31847;
    wire N__31840;
    wire N__31837;
    wire N__31834;
    wire N__31831;
    wire N__31828;
    wire N__31827;
    wire N__31824;
    wire N__31821;
    wire N__31820;
    wire N__31815;
    wire N__31812;
    wire N__31809;
    wire N__31804;
    wire N__31801;
    wire N__31798;
    wire N__31795;
    wire N__31792;
    wire N__31789;
    wire N__31786;
    wire N__31783;
    wire N__31780;
    wire N__31777;
    wire N__31776;
    wire N__31773;
    wire N__31770;
    wire N__31769;
    wire N__31768;
    wire N__31767;
    wire N__31766;
    wire N__31763;
    wire N__31760;
    wire N__31757;
    wire N__31754;
    wire N__31753;
    wire N__31752;
    wire N__31751;
    wire N__31750;
    wire N__31747;
    wire N__31744;
    wire N__31741;
    wire N__31736;
    wire N__31733;
    wire N__31730;
    wire N__31727;
    wire N__31726;
    wire N__31723;
    wire N__31720;
    wire N__31719;
    wire N__31716;
    wire N__31713;
    wire N__31708;
    wire N__31703;
    wire N__31700;
    wire N__31697;
    wire N__31694;
    wire N__31691;
    wire N__31688;
    wire N__31685;
    wire N__31682;
    wire N__31677;
    wire N__31672;
    wire N__31665;
    wire N__31662;
    wire N__31659;
    wire N__31654;
    wire N__31651;
    wire N__31648;
    wire N__31641;
    wire N__31636;
    wire N__31633;
    wire N__31630;
    wire N__31627;
    wire N__31624;
    wire N__31621;
    wire N__31618;
    wire N__31615;
    wire N__31612;
    wire N__31609;
    wire N__31606;
    wire N__31603;
    wire N__31600;
    wire N__31597;
    wire N__31594;
    wire N__31591;
    wire N__31588;
    wire N__31587;
    wire N__31584;
    wire N__31581;
    wire N__31578;
    wire N__31575;
    wire N__31572;
    wire N__31569;
    wire N__31566;
    wire N__31563;
    wire N__31560;
    wire N__31557;
    wire N__31554;
    wire N__31551;
    wire N__31548;
    wire N__31545;
    wire N__31542;
    wire N__31537;
    wire N__31534;
    wire N__31533;
    wire N__31530;
    wire N__31529;
    wire N__31526;
    wire N__31523;
    wire N__31520;
    wire N__31513;
    wire N__31510;
    wire N__31507;
    wire N__31504;
    wire N__31501;
    wire N__31498;
    wire N__31495;
    wire N__31492;
    wire N__31489;
    wire N__31488;
    wire N__31483;
    wire N__31480;
    wire N__31477;
    wire N__31474;
    wire N__31471;
    wire N__31468;
    wire N__31465;
    wire N__31462;
    wire N__31459;
    wire N__31456;
    wire N__31453;
    wire N__31450;
    wire N__31447;
    wire N__31444;
    wire N__31441;
    wire N__31438;
    wire N__31435;
    wire N__31434;
    wire N__31431;
    wire N__31428;
    wire N__31425;
    wire N__31422;
    wire N__31419;
    wire N__31416;
    wire N__31413;
    wire N__31410;
    wire N__31407;
    wire N__31404;
    wire N__31401;
    wire N__31398;
    wire N__31395;
    wire N__31392;
    wire N__31389;
    wire N__31384;
    wire N__31381;
    wire N__31378;
    wire N__31377;
    wire N__31376;
    wire N__31373;
    wire N__31370;
    wire N__31367;
    wire N__31364;
    wire N__31357;
    wire N__31356;
    wire N__31353;
    wire N__31350;
    wire N__31347;
    wire N__31342;
    wire N__31339;
    wire N__31336;
    wire N__31333;
    wire N__31332;
    wire N__31329;
    wire N__31326;
    wire N__31323;
    wire N__31320;
    wire N__31317;
    wire N__31312;
    wire N__31309;
    wire N__31306;
    wire N__31303;
    wire N__31302;
    wire N__31299;
    wire N__31296;
    wire N__31293;
    wire N__31288;
    wire N__31287;
    wire N__31284;
    wire N__31281;
    wire N__31278;
    wire N__31273;
    wire N__31270;
    wire N__31267;
    wire N__31264;
    wire N__31261;
    wire N__31258;
    wire N__31255;
    wire N__31252;
    wire N__31249;
    wire N__31246;
    wire N__31243;
    wire N__31240;
    wire N__31237;
    wire N__31234;
    wire N__31231;
    wire N__31228;
    wire N__31225;
    wire N__31222;
    wire N__31221;
    wire N__31218;
    wire N__31215;
    wire N__31212;
    wire N__31207;
    wire N__31204;
    wire N__31201;
    wire N__31198;
    wire N__31195;
    wire N__31194;
    wire N__31191;
    wire N__31188;
    wire N__31185;
    wire N__31180;
    wire N__31177;
    wire N__31176;
    wire N__31173;
    wire N__31170;
    wire N__31167;
    wire N__31164;
    wire N__31159;
    wire N__31156;
    wire N__31153;
    wire N__31150;
    wire N__31147;
    wire N__31146;
    wire N__31143;
    wire N__31140;
    wire N__31137;
    wire N__31134;
    wire N__31131;
    wire N__31126;
    wire N__31123;
    wire N__31120;
    wire N__31117;
    wire N__31114;
    wire N__31111;
    wire N__31108;
    wire N__31105;
    wire N__31102;
    wire N__31099;
    wire N__31096;
    wire N__31093;
    wire N__31090;
    wire N__31087;
    wire N__31084;
    wire N__31081;
    wire N__31078;
    wire N__31075;
    wire N__31072;
    wire N__31069;
    wire N__31066;
    wire N__31063;
    wire N__31060;
    wire N__31057;
    wire N__31054;
    wire N__31051;
    wire N__31048;
    wire N__31045;
    wire N__31042;
    wire N__31039;
    wire N__31036;
    wire N__31033;
    wire N__31030;
    wire N__31027;
    wire N__31024;
    wire N__31021;
    wire N__31018;
    wire N__31015;
    wire N__31012;
    wire N__31009;
    wire N__31006;
    wire N__31003;
    wire N__31000;
    wire N__30999;
    wire N__30994;
    wire N__30993;
    wire N__30992;
    wire N__30991;
    wire N__30990;
    wire N__30989;
    wire N__30986;
    wire N__30983;
    wire N__30980;
    wire N__30977;
    wire N__30972;
    wire N__30969;
    wire N__30966;
    wire N__30959;
    wire N__30956;
    wire N__30953;
    wire N__30950;
    wire N__30943;
    wire N__30940;
    wire N__30939;
    wire N__30936;
    wire N__30933;
    wire N__30932;
    wire N__30931;
    wire N__30930;
    wire N__30929;
    wire N__30928;
    wire N__30925;
    wire N__30922;
    wire N__30917;
    wire N__30912;
    wire N__30909;
    wire N__30898;
    wire N__30895;
    wire N__30892;
    wire N__30889;
    wire N__30886;
    wire N__30883;
    wire N__30880;
    wire N__30877;
    wire N__30874;
    wire N__30871;
    wire N__30868;
    wire N__30865;
    wire N__30862;
    wire N__30859;
    wire N__30856;
    wire N__30853;
    wire N__30850;
    wire N__30847;
    wire N__30844;
    wire N__30841;
    wire N__30838;
    wire N__30835;
    wire N__30832;
    wire N__30829;
    wire N__30826;
    wire N__30823;
    wire N__30820;
    wire N__30817;
    wire N__30814;
    wire N__30811;
    wire N__30810;
    wire N__30807;
    wire N__30804;
    wire N__30803;
    wire N__30800;
    wire N__30797;
    wire N__30794;
    wire N__30791;
    wire N__30788;
    wire N__30785;
    wire N__30778;
    wire N__30775;
    wire N__30772;
    wire N__30771;
    wire N__30770;
    wire N__30767;
    wire N__30764;
    wire N__30761;
    wire N__30754;
    wire N__30751;
    wire N__30748;
    wire N__30745;
    wire N__30744;
    wire N__30741;
    wire N__30740;
    wire N__30739;
    wire N__30736;
    wire N__30729;
    wire N__30724;
    wire N__30723;
    wire N__30722;
    wire N__30721;
    wire N__30718;
    wire N__30711;
    wire N__30706;
    wire N__30703;
    wire N__30702;
    wire N__30701;
    wire N__30698;
    wire N__30693;
    wire N__30688;
    wire N__30685;
    wire N__30682;
    wire N__30679;
    wire N__30676;
    wire N__30673;
    wire N__30670;
    wire N__30667;
    wire N__30664;
    wire N__30663;
    wire N__30660;
    wire N__30657;
    wire N__30654;
    wire N__30649;
    wire N__30646;
    wire N__30643;
    wire N__30640;
    wire N__30637;
    wire N__30636;
    wire N__30633;
    wire N__30630;
    wire N__30625;
    wire N__30624;
    wire N__30623;
    wire N__30616;
    wire N__30613;
    wire N__30610;
    wire N__30607;
    wire N__30604;
    wire N__30601;
    wire N__30598;
    wire N__30595;
    wire N__30594;
    wire N__30591;
    wire N__30588;
    wire N__30583;
    wire N__30580;
    wire N__30579;
    wire N__30576;
    wire N__30573;
    wire N__30568;
    wire N__30567;
    wire N__30564;
    wire N__30561;
    wire N__30558;
    wire N__30553;
    wire N__30550;
    wire N__30549;
    wire N__30546;
    wire N__30543;
    wire N__30538;
    wire N__30535;
    wire N__30532;
    wire N__30529;
    wire N__30528;
    wire N__30525;
    wire N__30522;
    wire N__30519;
    wire N__30516;
    wire N__30511;
    wire N__30508;
    wire N__30505;
    wire N__30502;
    wire N__30499;
    wire N__30496;
    wire N__30493;
    wire N__30490;
    wire N__30487;
    wire N__30484;
    wire N__30481;
    wire N__30478;
    wire N__30475;
    wire N__30472;
    wire N__30469;
    wire N__30466;
    wire N__30463;
    wire N__30462;
    wire N__30461;
    wire N__30458;
    wire N__30455;
    wire N__30454;
    wire N__30451;
    wire N__30448;
    wire N__30443;
    wire N__30442;
    wire N__30439;
    wire N__30436;
    wire N__30433;
    wire N__30430;
    wire N__30427;
    wire N__30422;
    wire N__30415;
    wire N__30412;
    wire N__30409;
    wire N__30406;
    wire N__30403;
    wire N__30400;
    wire N__30397;
    wire N__30394;
    wire N__30391;
    wire N__30390;
    wire N__30387;
    wire N__30384;
    wire N__30379;
    wire N__30378;
    wire N__30375;
    wire N__30372;
    wire N__30367;
    wire N__30366;
    wire N__30363;
    wire N__30360;
    wire N__30357;
    wire N__30354;
    wire N__30349;
    wire N__30348;
    wire N__30345;
    wire N__30342;
    wire N__30337;
    wire N__30334;
    wire N__30333;
    wire N__30330;
    wire N__30327;
    wire N__30322;
    wire N__30319;
    wire N__30318;
    wire N__30315;
    wire N__30312;
    wire N__30307;
    wire N__30306;
    wire N__30303;
    wire N__30300;
    wire N__30297;
    wire N__30292;
    wire N__30291;
    wire N__30288;
    wire N__30285;
    wire N__30280;
    wire N__30277;
    wire N__30274;
    wire N__30271;
    wire N__30270;
    wire N__30267;
    wire N__30264;
    wire N__30259;
    wire N__30258;
    wire N__30255;
    wire N__30252;
    wire N__30247;
    wire N__30246;
    wire N__30243;
    wire N__30240;
    wire N__30237;
    wire N__30232;
    wire N__30231;
    wire N__30228;
    wire N__30225;
    wire N__30220;
    wire N__30217;
    wire N__30214;
    wire N__30211;
    wire N__30208;
    wire N__30205;
    wire N__30204;
    wire N__30203;
    wire N__30200;
    wire N__30197;
    wire N__30194;
    wire N__30187;
    wire N__30186;
    wire N__30185;
    wire N__30182;
    wire N__30179;
    wire N__30176;
    wire N__30173;
    wire N__30170;
    wire N__30163;
    wire N__30160;
    wire N__30157;
    wire N__30154;
    wire N__30151;
    wire N__30148;
    wire N__30145;
    wire N__30142;
    wire N__30141;
    wire N__30140;
    wire N__30139;
    wire N__30134;
    wire N__30133;
    wire N__30128;
    wire N__30125;
    wire N__30122;
    wire N__30119;
    wire N__30116;
    wire N__30111;
    wire N__30106;
    wire N__30103;
    wire N__30100;
    wire N__30099;
    wire N__30096;
    wire N__30093;
    wire N__30090;
    wire N__30087;
    wire N__30084;
    wire N__30079;
    wire N__30078;
    wire N__30075;
    wire N__30072;
    wire N__30069;
    wire N__30064;
    wire N__30061;
    wire N__30058;
    wire N__30055;
    wire N__30052;
    wire N__30049;
    wire N__30046;
    wire N__30045;
    wire N__30042;
    wire N__30041;
    wire N__30038;
    wire N__30035;
    wire N__30032;
    wire N__30029;
    wire N__30022;
    wire N__30021;
    wire N__30018;
    wire N__30015;
    wire N__30014;
    wire N__30013;
    wire N__30012;
    wire N__30009;
    wire N__30006;
    wire N__30005;
    wire N__30004;
    wire N__30003;
    wire N__30000;
    wire N__29999;
    wire N__29996;
    wire N__29995;
    wire N__29994;
    wire N__29991;
    wire N__29990;
    wire N__29987;
    wire N__29984;
    wire N__29981;
    wire N__29974;
    wire N__29961;
    wire N__29950;
    wire N__29949;
    wire N__29946;
    wire N__29943;
    wire N__29940;
    wire N__29937;
    wire N__29936;
    wire N__29935;
    wire N__29934;
    wire N__29933;
    wire N__29932;
    wire N__29931;
    wire N__29930;
    wire N__29929;
    wire N__29928;
    wire N__29927;
    wire N__29924;
    wire N__29921;
    wire N__29918;
    wire N__29909;
    wire N__29898;
    wire N__29887;
    wire N__29886;
    wire N__29883;
    wire N__29880;
    wire N__29879;
    wire N__29876;
    wire N__29873;
    wire N__29870;
    wire N__29863;
    wire N__29862;
    wire N__29859;
    wire N__29858;
    wire N__29857;
    wire N__29856;
    wire N__29855;
    wire N__29854;
    wire N__29851;
    wire N__29848;
    wire N__29847;
    wire N__29846;
    wire N__29845;
    wire N__29842;
    wire N__29841;
    wire N__29838;
    wire N__29837;
    wire N__29830;
    wire N__29827;
    wire N__29824;
    wire N__29819;
    wire N__29808;
    wire N__29805;
    wire N__29794;
    wire N__29793;
    wire N__29792;
    wire N__29791;
    wire N__29788;
    wire N__29787;
    wire N__29784;
    wire N__29783;
    wire N__29782;
    wire N__29781;
    wire N__29776;
    wire N__29773;
    wire N__29768;
    wire N__29767;
    wire N__29766;
    wire N__29765;
    wire N__29764;
    wire N__29757;
    wire N__29754;
    wire N__29749;
    wire N__29742;
    wire N__29739;
    wire N__29736;
    wire N__29725;
    wire N__29722;
    wire N__29719;
    wire N__29716;
    wire N__29715;
    wire N__29712;
    wire N__29709;
    wire N__29706;
    wire N__29705;
    wire N__29702;
    wire N__29699;
    wire N__29696;
    wire N__29693;
    wire N__29686;
    wire N__29683;
    wire N__29680;
    wire N__29677;
    wire N__29674;
    wire N__29671;
    wire N__29668;
    wire N__29665;
    wire N__29662;
    wire N__29659;
    wire N__29656;
    wire N__29653;
    wire N__29650;
    wire N__29647;
    wire N__29644;
    wire N__29641;
    wire N__29638;
    wire N__29635;
    wire N__29632;
    wire N__29629;
    wire N__29626;
    wire N__29623;
    wire N__29620;
    wire N__29617;
    wire N__29614;
    wire N__29611;
    wire N__29608;
    wire N__29607;
    wire N__29604;
    wire N__29601;
    wire N__29598;
    wire N__29595;
    wire N__29590;
    wire N__29587;
    wire N__29586;
    wire N__29583;
    wire N__29580;
    wire N__29577;
    wire N__29576;
    wire N__29573;
    wire N__29570;
    wire N__29567;
    wire N__29562;
    wire N__29557;
    wire N__29556;
    wire N__29555;
    wire N__29552;
    wire N__29549;
    wire N__29546;
    wire N__29543;
    wire N__29536;
    wire N__29533;
    wire N__29530;
    wire N__29527;
    wire N__29524;
    wire N__29521;
    wire N__29518;
    wire N__29515;
    wire N__29512;
    wire N__29509;
    wire N__29508;
    wire N__29505;
    wire N__29502;
    wire N__29499;
    wire N__29498;
    wire N__29493;
    wire N__29490;
    wire N__29487;
    wire N__29482;
    wire N__29479;
    wire N__29476;
    wire N__29475;
    wire N__29474;
    wire N__29473;
    wire N__29472;
    wire N__29471;
    wire N__29470;
    wire N__29459;
    wire N__29454;
    wire N__29449;
    wire N__29448;
    wire N__29447;
    wire N__29440;
    wire N__29437;
    wire N__29436;
    wire N__29433;
    wire N__29432;
    wire N__29425;
    wire N__29422;
    wire N__29421;
    wire N__29420;
    wire N__29417;
    wire N__29412;
    wire N__29407;
    wire N__29404;
    wire N__29401;
    wire N__29398;
    wire N__29397;
    wire N__29394;
    wire N__29393;
    wire N__29390;
    wire N__29387;
    wire N__29384;
    wire N__29377;
    wire N__29374;
    wire N__29371;
    wire N__29368;
    wire N__29365;
    wire N__29362;
    wire N__29359;
    wire N__29356;
    wire N__29353;
    wire N__29350;
    wire N__29347;
    wire N__29344;
    wire N__29341;
    wire N__29338;
    wire N__29335;
    wire N__29332;
    wire N__29329;
    wire N__29326;
    wire N__29325;
    wire N__29322;
    wire N__29319;
    wire N__29318;
    wire N__29317;
    wire N__29314;
    wire N__29311;
    wire N__29308;
    wire N__29305;
    wire N__29300;
    wire N__29297;
    wire N__29296;
    wire N__29293;
    wire N__29288;
    wire N__29285;
    wire N__29282;
    wire N__29275;
    wire N__29272;
    wire N__29271;
    wire N__29268;
    wire N__29265;
    wire N__29260;
    wire N__29257;
    wire N__29254;
    wire N__29253;
    wire N__29250;
    wire N__29247;
    wire N__29244;
    wire N__29239;
    wire N__29236;
    wire N__29235;
    wire N__29232;
    wire N__29229;
    wire N__29224;
    wire N__29221;
    wire N__29220;
    wire N__29217;
    wire N__29214;
    wire N__29209;
    wire N__29206;
    wire N__29203;
    wire N__29202;
    wire N__29199;
    wire N__29196;
    wire N__29191;
    wire N__29190;
    wire N__29187;
    wire N__29186;
    wire N__29183;
    wire N__29180;
    wire N__29179;
    wire N__29178;
    wire N__29177;
    wire N__29174;
    wire N__29169;
    wire N__29166;
    wire N__29163;
    wire N__29162;
    wire N__29159;
    wire N__29152;
    wire N__29149;
    wire N__29146;
    wire N__29143;
    wire N__29140;
    wire N__29135;
    wire N__29134;
    wire N__29131;
    wire N__29128;
    wire N__29125;
    wire N__29122;
    wire N__29113;
    wire N__29110;
    wire N__29109;
    wire N__29108;
    wire N__29105;
    wire N__29104;
    wire N__29103;
    wire N__29100;
    wire N__29099;
    wire N__29096;
    wire N__29095;
    wire N__29092;
    wire N__29089;
    wire N__29086;
    wire N__29083;
    wire N__29080;
    wire N__29077;
    wire N__29074;
    wire N__29069;
    wire N__29066;
    wire N__29061;
    wire N__29056;
    wire N__29051;
    wire N__29048;
    wire N__29045;
    wire N__29042;
    wire N__29035;
    wire N__29032;
    wire N__29029;
    wire N__29026;
    wire N__29023;
    wire N__29020;
    wire N__29017;
    wire N__29014;
    wire N__29011;
    wire N__29008;
    wire N__29005;
    wire N__29002;
    wire N__28999;
    wire N__28996;
    wire N__28993;
    wire N__28990;
    wire N__28987;
    wire N__28984;
    wire N__28981;
    wire N__28980;
    wire N__28979;
    wire N__28978;
    wire N__28977;
    wire N__28976;
    wire N__28975;
    wire N__28974;
    wire N__28973;
    wire N__28968;
    wire N__28955;
    wire N__28954;
    wire N__28953;
    wire N__28952;
    wire N__28951;
    wire N__28950;
    wire N__28949;
    wire N__28948;
    wire N__28947;
    wire N__28944;
    wire N__28943;
    wire N__28942;
    wire N__28941;
    wire N__28940;
    wire N__28937;
    wire N__28934;
    wire N__28931;
    wire N__28916;
    wire N__28913;
    wire N__28910;
    wire N__28909;
    wire N__28908;
    wire N__28907;
    wire N__28904;
    wire N__28899;
    wire N__28892;
    wire N__28889;
    wire N__28884;
    wire N__28881;
    wire N__28880;
    wire N__28877;
    wire N__28876;
    wire N__28873;
    wire N__28870;
    wire N__28867;
    wire N__28866;
    wire N__28865;
    wire N__28860;
    wire N__28855;
    wire N__28852;
    wire N__28849;
    wire N__28846;
    wire N__28841;
    wire N__28838;
    wire N__28833;
    wire N__28830;
    wire N__28827;
    wire N__28810;
    wire N__28809;
    wire N__28808;
    wire N__28807;
    wire N__28806;
    wire N__28805;
    wire N__28804;
    wire N__28803;
    wire N__28802;
    wire N__28801;
    wire N__28800;
    wire N__28799;
    wire N__28798;
    wire N__28797;
    wire N__28796;
    wire N__28795;
    wire N__28788;
    wire N__28777;
    wire N__28776;
    wire N__28775;
    wire N__28774;
    wire N__28773;
    wire N__28756;
    wire N__28751;
    wire N__28750;
    wire N__28749;
    wire N__28748;
    wire N__28747;
    wire N__28746;
    wire N__28743;
    wire N__28740;
    wire N__28737;
    wire N__28736;
    wire N__28733;
    wire N__28728;
    wire N__28725;
    wire N__28716;
    wire N__28711;
    wire N__28708;
    wire N__28705;
    wire N__28702;
    wire N__28699;
    wire N__28694;
    wire N__28689;
    wire N__28678;
    wire N__28677;
    wire N__28674;
    wire N__28671;
    wire N__28668;
    wire N__28665;
    wire N__28664;
    wire N__28661;
    wire N__28658;
    wire N__28655;
    wire N__28654;
    wire N__28649;
    wire N__28646;
    wire N__28643;
    wire N__28640;
    wire N__28637;
    wire N__28634;
    wire N__28631;
    wire N__28628;
    wire N__28621;
    wire N__28618;
    wire N__28617;
    wire N__28614;
    wire N__28613;
    wire N__28612;
    wire N__28611;
    wire N__28608;
    wire N__28607;
    wire N__28604;
    wire N__28601;
    wire N__28598;
    wire N__28595;
    wire N__28594;
    wire N__28593;
    wire N__28592;
    wire N__28591;
    wire N__28588;
    wire N__28585;
    wire N__28582;
    wire N__28575;
    wire N__28566;
    wire N__28555;
    wire N__28552;
    wire N__28551;
    wire N__28548;
    wire N__28545;
    wire N__28540;
    wire N__28537;
    wire N__28534;
    wire N__28531;
    wire N__28530;
    wire N__28527;
    wire N__28524;
    wire N__28519;
    wire N__28516;
    wire N__28515;
    wire N__28512;
    wire N__28509;
    wire N__28506;
    wire N__28501;
    wire N__28498;
    wire N__28497;
    wire N__28494;
    wire N__28491;
    wire N__28486;
    wire N__28483;
    wire N__28482;
    wire N__28479;
    wire N__28476;
    wire N__28473;
    wire N__28468;
    wire N__28465;
    wire N__28464;
    wire N__28461;
    wire N__28458;
    wire N__28453;
    wire N__28450;
    wire N__28449;
    wire N__28446;
    wire N__28443;
    wire N__28438;
    wire N__28435;
    wire N__28434;
    wire N__28431;
    wire N__28428;
    wire N__28423;
    wire N__28420;
    wire N__28419;
    wire N__28418;
    wire N__28417;
    wire N__28416;
    wire N__28415;
    wire N__28414;
    wire N__28399;
    wire N__28398;
    wire N__28397;
    wire N__28394;
    wire N__28391;
    wire N__28390;
    wire N__28389;
    wire N__28388;
    wire N__28385;
    wire N__28382;
    wire N__28373;
    wire N__28372;
    wire N__28371;
    wire N__28370;
    wire N__28369;
    wire N__28368;
    wire N__28367;
    wire N__28366;
    wire N__28365;
    wire N__28364;
    wire N__28363;
    wire N__28362;
    wire N__28361;
    wire N__28354;
    wire N__28337;
    wire N__28330;
    wire N__28327;
    wire N__28324;
    wire N__28321;
    wire N__28318;
    wire N__28315;
    wire N__28312;
    wire N__28307;
    wire N__28300;
    wire N__28297;
    wire N__28294;
    wire N__28291;
    wire N__28288;
    wire N__28285;
    wire N__28282;
    wire N__28279;
    wire N__28276;
    wire N__28273;
    wire N__28270;
    wire N__28267;
    wire N__28264;
    wire N__28261;
    wire N__28258;
    wire N__28255;
    wire N__28252;
    wire N__28249;
    wire N__28246;
    wire N__28243;
    wire N__28240;
    wire N__28237;
    wire N__28234;
    wire N__28231;
    wire N__28228;
    wire N__28225;
    wire N__28222;
    wire N__28219;
    wire N__28216;
    wire N__28213;
    wire N__28212;
    wire N__28211;
    wire N__28208;
    wire N__28205;
    wire N__28202;
    wire N__28195;
    wire N__28192;
    wire N__28189;
    wire N__28186;
    wire N__28183;
    wire N__28180;
    wire N__28177;
    wire N__28174;
    wire N__28171;
    wire N__28168;
    wire N__28165;
    wire N__28162;
    wire N__28161;
    wire N__28158;
    wire N__28157;
    wire N__28154;
    wire N__28151;
    wire N__28146;
    wire N__28143;
    wire N__28138;
    wire N__28135;
    wire N__28134;
    wire N__28131;
    wire N__28128;
    wire N__28125;
    wire N__28122;
    wire N__28121;
    wire N__28118;
    wire N__28115;
    wire N__28112;
    wire N__28109;
    wire N__28106;
    wire N__28099;
    wire N__28096;
    wire N__28093;
    wire N__28090;
    wire N__28087;
    wire N__28086;
    wire N__28085;
    wire N__28082;
    wire N__28079;
    wire N__28076;
    wire N__28073;
    wire N__28070;
    wire N__28067;
    wire N__28060;
    wire N__28057;
    wire N__28054;
    wire N__28051;
    wire N__28050;
    wire N__28047;
    wire N__28046;
    wire N__28043;
    wire N__28040;
    wire N__28037;
    wire N__28034;
    wire N__28027;
    wire N__28024;
    wire N__28021;
    wire N__28018;
    wire N__28015;
    wire N__28014;
    wire N__28013;
    wire N__28010;
    wire N__28007;
    wire N__28004;
    wire N__27997;
    wire N__27994;
    wire N__27993;
    wire N__27992;
    wire N__27989;
    wire N__27986;
    wire N__27983;
    wire N__27980;
    wire N__27977;
    wire N__27974;
    wire N__27971;
    wire N__27964;
    wire N__27963;
    wire N__27960;
    wire N__27959;
    wire N__27956;
    wire N__27953;
    wire N__27950;
    wire N__27943;
    wire N__27940;
    wire N__27937;
    wire N__27934;
    wire N__27931;
    wire N__27928;
    wire N__27925;
    wire N__27922;
    wire N__27921;
    wire N__27920;
    wire N__27917;
    wire N__27914;
    wire N__27911;
    wire N__27908;
    wire N__27901;
    wire N__27898;
    wire N__27895;
    wire N__27892;
    wire N__27889;
    wire N__27886;
    wire N__27883;
    wire N__27880;
    wire N__27877;
    wire N__27874;
    wire N__27873;
    wire N__27870;
    wire N__27867;
    wire N__27864;
    wire N__27861;
    wire N__27858;
    wire N__27857;
    wire N__27854;
    wire N__27851;
    wire N__27848;
    wire N__27845;
    wire N__27838;
    wire N__27835;
    wire N__27832;
    wire N__27829;
    wire N__27826;
    wire N__27825;
    wire N__27824;
    wire N__27821;
    wire N__27816;
    wire N__27811;
    wire N__27808;
    wire N__27805;
    wire N__27802;
    wire N__27801;
    wire N__27800;
    wire N__27797;
    wire N__27794;
    wire N__27791;
    wire N__27788;
    wire N__27785;
    wire N__27778;
    wire N__27777;
    wire N__27774;
    wire N__27773;
    wire N__27770;
    wire N__27767;
    wire N__27764;
    wire N__27757;
    wire N__27756;
    wire N__27753;
    wire N__27750;
    wire N__27747;
    wire N__27746;
    wire N__27743;
    wire N__27740;
    wire N__27737;
    wire N__27730;
    wire N__27727;
    wire N__27726;
    wire N__27723;
    wire N__27720;
    wire N__27717;
    wire N__27714;
    wire N__27709;
    wire N__27706;
    wire N__27703;
    wire N__27700;
    wire N__27697;
    wire N__27694;
    wire N__27691;
    wire N__27688;
    wire N__27685;
    wire N__27682;
    wire N__27679;
    wire N__27676;
    wire N__27673;
    wire N__27670;
    wire N__27667;
    wire N__27664;
    wire N__27661;
    wire N__27658;
    wire N__27655;
    wire N__27652;
    wire N__27649;
    wire N__27646;
    wire N__27643;
    wire N__27640;
    wire N__27637;
    wire N__27634;
    wire N__27631;
    wire N__27628;
    wire N__27625;
    wire N__27622;
    wire N__27619;
    wire N__27616;
    wire N__27613;
    wire N__27610;
    wire N__27609;
    wire N__27608;
    wire N__27605;
    wire N__27602;
    wire N__27599;
    wire N__27596;
    wire N__27589;
    wire N__27588;
    wire N__27587;
    wire N__27584;
    wire N__27581;
    wire N__27578;
    wire N__27571;
    wire N__27570;
    wire N__27567;
    wire N__27566;
    wire N__27563;
    wire N__27560;
    wire N__27557;
    wire N__27554;
    wire N__27551;
    wire N__27544;
    wire N__27541;
    wire N__27538;
    wire N__27535;
    wire N__27532;
    wire N__27529;
    wire N__27526;
    wire N__27523;
    wire N__27520;
    wire N__27517;
    wire N__27514;
    wire N__27513;
    wire N__27512;
    wire N__27509;
    wire N__27506;
    wire N__27505;
    wire N__27504;
    wire N__27501;
    wire N__27496;
    wire N__27493;
    wire N__27490;
    wire N__27487;
    wire N__27484;
    wire N__27481;
    wire N__27478;
    wire N__27469;
    wire N__27466;
    wire N__27465;
    wire N__27464;
    wire N__27461;
    wire N__27458;
    wire N__27455;
    wire N__27454;
    wire N__27453;
    wire N__27448;
    wire N__27445;
    wire N__27442;
    wire N__27439;
    wire N__27436;
    wire N__27433;
    wire N__27430;
    wire N__27427;
    wire N__27418;
    wire N__27415;
    wire N__27412;
    wire N__27409;
    wire N__27406;
    wire N__27403;
    wire N__27400;
    wire N__27397;
    wire N__27394;
    wire N__27391;
    wire N__27388;
    wire N__27385;
    wire N__27382;
    wire N__27379;
    wire N__27376;
    wire N__27373;
    wire N__27370;
    wire N__27367;
    wire N__27364;
    wire N__27361;
    wire N__27358;
    wire N__27355;
    wire N__27352;
    wire N__27349;
    wire N__27346;
    wire N__27343;
    wire N__27340;
    wire N__27337;
    wire N__27334;
    wire N__27331;
    wire N__27328;
    wire N__27325;
    wire N__27322;
    wire N__27319;
    wire N__27316;
    wire N__27313;
    wire N__27310;
    wire N__27307;
    wire N__27304;
    wire N__27301;
    wire N__27300;
    wire N__27297;
    wire N__27294;
    wire N__27291;
    wire N__27288;
    wire N__27287;
    wire N__27284;
    wire N__27281;
    wire N__27278;
    wire N__27275;
    wire N__27272;
    wire N__27265;
    wire N__27262;
    wire N__27259;
    wire N__27256;
    wire N__27253;
    wire N__27250;
    wire N__27247;
    wire N__27244;
    wire N__27241;
    wire N__27238;
    wire N__27235;
    wire N__27232;
    wire N__27229;
    wire N__27226;
    wire N__27223;
    wire N__27220;
    wire N__27217;
    wire N__27214;
    wire N__27211;
    wire N__27208;
    wire N__27205;
    wire N__27202;
    wire N__27199;
    wire N__27196;
    wire N__27193;
    wire N__27190;
    wire N__27187;
    wire N__27184;
    wire N__27181;
    wire N__27178;
    wire N__27175;
    wire N__27172;
    wire N__27169;
    wire N__27166;
    wire N__27163;
    wire N__27160;
    wire N__27157;
    wire N__27154;
    wire N__27151;
    wire N__27148;
    wire N__27145;
    wire N__27142;
    wire N__27139;
    wire N__27136;
    wire N__27133;
    wire N__27130;
    wire N__27127;
    wire N__27124;
    wire N__27121;
    wire N__27118;
    wire N__27115;
    wire N__27114;
    wire N__27111;
    wire N__27108;
    wire N__27103;
    wire N__27102;
    wire N__27099;
    wire N__27096;
    wire N__27091;
    wire N__27088;
    wire N__27087;
    wire N__27084;
    wire N__27081;
    wire N__27076;
    wire N__27073;
    wire N__27070;
    wire N__27067;
    wire N__27064;
    wire N__27061;
    wire N__27058;
    wire N__27055;
    wire N__27052;
    wire N__27049;
    wire N__27048;
    wire N__27047;
    wire N__27044;
    wire N__27041;
    wire N__27038;
    wire N__27031;
    wire N__27028;
    wire N__27025;
    wire N__27022;
    wire N__27019;
    wire N__27016;
    wire N__27013;
    wire N__27010;
    wire N__27007;
    wire N__27004;
    wire N__27001;
    wire N__26998;
    wire N__26995;
    wire N__26992;
    wire N__26989;
    wire N__26988;
    wire N__26985;
    wire N__26984;
    wire N__26981;
    wire N__26978;
    wire N__26975;
    wire N__26972;
    wire N__26969;
    wire N__26966;
    wire N__26959;
    wire N__26958;
    wire N__26957;
    wire N__26954;
    wire N__26949;
    wire N__26946;
    wire N__26941;
    wire N__26938;
    wire N__26935;
    wire N__26932;
    wire N__26931;
    wire N__26928;
    wire N__26925;
    wire N__26920;
    wire N__26919;
    wire N__26916;
    wire N__26915;
    wire N__26912;
    wire N__26909;
    wire N__26906;
    wire N__26903;
    wire N__26896;
    wire N__26895;
    wire N__26892;
    wire N__26891;
    wire N__26890;
    wire N__26889;
    wire N__26888;
    wire N__26885;
    wire N__26884;
    wire N__26883;
    wire N__26882;
    wire N__26881;
    wire N__26880;
    wire N__26879;
    wire N__26878;
    wire N__26875;
    wire N__26864;
    wire N__26861;
    wire N__26858;
    wire N__26855;
    wire N__26852;
    wire N__26851;
    wire N__26850;
    wire N__26847;
    wire N__26846;
    wire N__26843;
    wire N__26842;
    wire N__26841;
    wire N__26838;
    wire N__26837;
    wire N__26836;
    wire N__26831;
    wire N__26818;
    wire N__26805;
    wire N__26802;
    wire N__26799;
    wire N__26798;
    wire N__26797;
    wire N__26792;
    wire N__26789;
    wire N__26780;
    wire N__26773;
    wire N__26770;
    wire N__26769;
    wire N__26768;
    wire N__26765;
    wire N__26762;
    wire N__26759;
    wire N__26756;
    wire N__26753;
    wire N__26746;
    wire N__26745;
    wire N__26742;
    wire N__26739;
    wire N__26734;
    wire N__26731;
    wire N__26728;
    wire N__26727;
    wire N__26724;
    wire N__26721;
    wire N__26718;
    wire N__26715;
    wire N__26710;
    wire N__26709;
    wire N__26706;
    wire N__26703;
    wire N__26698;
    wire N__26695;
    wire N__26692;
    wire N__26691;
    wire N__26688;
    wire N__26685;
    wire N__26682;
    wire N__26679;
    wire N__26674;
    wire N__26671;
    wire N__26670;
    wire N__26667;
    wire N__26664;
    wire N__26659;
    wire N__26658;
    wire N__26655;
    wire N__26652;
    wire N__26647;
    wire N__26646;
    wire N__26643;
    wire N__26640;
    wire N__26635;
    wire N__26632;
    wire N__26629;
    wire N__26628;
    wire N__26625;
    wire N__26622;
    wire N__26619;
    wire N__26616;
    wire N__26611;
    wire N__26610;
    wire N__26609;
    wire N__26606;
    wire N__26603;
    wire N__26600;
    wire N__26597;
    wire N__26590;
    wire N__26587;
    wire N__26586;
    wire N__26585;
    wire N__26582;
    wire N__26577;
    wire N__26574;
    wire N__26569;
    wire N__26568;
    wire N__26565;
    wire N__26564;
    wire N__26561;
    wire N__26558;
    wire N__26555;
    wire N__26552;
    wire N__26545;
    wire N__26542;
    wire N__26539;
    wire N__26536;
    wire N__26533;
    wire N__26532;
    wire N__26529;
    wire N__26528;
    wire N__26525;
    wire N__26522;
    wire N__26519;
    wire N__26514;
    wire N__26509;
    wire N__26508;
    wire N__26505;
    wire N__26504;
    wire N__26501;
    wire N__26498;
    wire N__26495;
    wire N__26492;
    wire N__26485;
    wire N__26482;
    wire N__26481;
    wire N__26480;
    wire N__26477;
    wire N__26474;
    wire N__26471;
    wire N__26468;
    wire N__26465;
    wire N__26458;
    wire N__26455;
    wire N__26452;
    wire N__26451;
    wire N__26450;
    wire N__26447;
    wire N__26444;
    wire N__26441;
    wire N__26438;
    wire N__26435;
    wire N__26428;
    wire N__26427;
    wire N__26426;
    wire N__26423;
    wire N__26418;
    wire N__26415;
    wire N__26410;
    wire N__26409;
    wire N__26408;
    wire N__26405;
    wire N__26402;
    wire N__26399;
    wire N__26396;
    wire N__26389;
    wire N__26388;
    wire N__26387;
    wire N__26384;
    wire N__26381;
    wire N__26378;
    wire N__26375;
    wire N__26372;
    wire N__26365;
    wire N__26364;
    wire N__26363;
    wire N__26360;
    wire N__26357;
    wire N__26354;
    wire N__26351;
    wire N__26348;
    wire N__26345;
    wire N__26342;
    wire N__26335;
    wire N__26332;
    wire N__26329;
    wire N__26326;
    wire N__26323;
    wire N__26320;
    wire N__26317;
    wire N__26314;
    wire N__26311;
    wire N__26308;
    wire N__26307;
    wire N__26304;
    wire N__26301;
    wire N__26296;
    wire N__26293;
    wire N__26292;
    wire N__26289;
    wire N__26286;
    wire N__26283;
    wire N__26280;
    wire N__26275;
    wire N__26272;
    wire N__26269;
    wire N__26266;
    wire N__26263;
    wire N__26262;
    wire N__26259;
    wire N__26258;
    wire N__26255;
    wire N__26252;
    wire N__26247;
    wire N__26242;
    wire N__26239;
    wire N__26236;
    wire N__26233;
    wire N__26230;
    wire N__26227;
    wire N__26224;
    wire N__26221;
    wire N__26218;
    wire N__26215;
    wire N__26212;
    wire N__26209;
    wire N__26208;
    wire N__26207;
    wire N__26204;
    wire N__26199;
    wire N__26194;
    wire N__26191;
    wire N__26188;
    wire N__26185;
    wire N__26184;
    wire N__26181;
    wire N__26178;
    wire N__26175;
    wire N__26172;
    wire N__26167;
    wire N__26164;
    wire N__26161;
    wire N__26158;
    wire N__26155;
    wire N__26152;
    wire N__26149;
    wire N__26148;
    wire N__26145;
    wire N__26142;
    wire N__26139;
    wire N__26136;
    wire N__26133;
    wire N__26130;
    wire N__26127;
    wire N__26124;
    wire N__26119;
    wire N__26116;
    wire N__26113;
    wire N__26110;
    wire N__26107;
    wire N__26104;
    wire N__26101;
    wire N__26100;
    wire N__26097;
    wire N__26096;
    wire N__26093;
    wire N__26090;
    wire N__26087;
    wire N__26084;
    wire N__26077;
    wire N__26074;
    wire N__26071;
    wire N__26070;
    wire N__26069;
    wire N__26066;
    wire N__26063;
    wire N__26060;
    wire N__26057;
    wire N__26054;
    wire N__26047;
    wire N__26044;
    wire N__26041;
    wire N__26038;
    wire N__26035;
    wire N__26032;
    wire N__26031;
    wire N__26028;
    wire N__26027;
    wire N__26024;
    wire N__26021;
    wire N__26016;
    wire N__26011;
    wire N__26008;
    wire N__26005;
    wire N__26002;
    wire N__25999;
    wire N__25996;
    wire N__25993;
    wire N__25992;
    wire N__25989;
    wire N__25986;
    wire N__25983;
    wire N__25982;
    wire N__25977;
    wire N__25974;
    wire N__25969;
    wire N__25968;
    wire N__25965;
    wire N__25962;
    wire N__25961;
    wire N__25958;
    wire N__25955;
    wire N__25952;
    wire N__25949;
    wire N__25946;
    wire N__25939;
    wire N__25938;
    wire N__25937;
    wire N__25934;
    wire N__25931;
    wire N__25930;
    wire N__25927;
    wire N__25920;
    wire N__25917;
    wire N__25912;
    wire N__25911;
    wire N__25910;
    wire N__25905;
    wire N__25902;
    wire N__25897;
    wire N__25894;
    wire N__25893;
    wire N__25890;
    wire N__25889;
    wire N__25886;
    wire N__25883;
    wire N__25880;
    wire N__25873;
    wire N__25872;
    wire N__25869;
    wire N__25866;
    wire N__25863;
    wire N__25860;
    wire N__25857;
    wire N__25856;
    wire N__25853;
    wire N__25850;
    wire N__25847;
    wire N__25840;
    wire N__25837;
    wire N__25834;
    wire N__25831;
    wire N__25828;
    wire N__25825;
    wire N__25822;
    wire N__25819;
    wire N__25816;
    wire N__25813;
    wire N__25812;
    wire N__25809;
    wire N__25808;
    wire N__25805;
    wire N__25802;
    wire N__25799;
    wire N__25796;
    wire N__25793;
    wire N__25786;
    wire N__25785;
    wire N__25782;
    wire N__25779;
    wire N__25774;
    wire N__25771;
    wire N__25768;
    wire N__25765;
    wire N__25762;
    wire N__25759;
    wire N__25756;
    wire N__25753;
    wire N__25750;
    wire N__25747;
    wire N__25746;
    wire N__25743;
    wire N__25740;
    wire N__25737;
    wire N__25734;
    wire N__25729;
    wire N__25726;
    wire N__25723;
    wire N__25720;
    wire N__25717;
    wire N__25714;
    wire N__25711;
    wire N__25710;
    wire N__25707;
    wire N__25706;
    wire N__25703;
    wire N__25700;
    wire N__25697;
    wire N__25694;
    wire N__25691;
    wire N__25688;
    wire N__25685;
    wire N__25682;
    wire N__25675;
    wire N__25672;
    wire N__25669;
    wire N__25668;
    wire N__25665;
    wire N__25662;
    wire N__25659;
    wire N__25656;
    wire N__25651;
    wire N__25648;
    wire N__25645;
    wire N__25642;
    wire N__25639;
    wire N__25636;
    wire N__25633;
    wire N__25630;
    wire N__25627;
    wire N__25624;
    wire N__25621;
    wire N__25618;
    wire N__25615;
    wire N__25612;
    wire N__25609;
    wire N__25606;
    wire N__25603;
    wire N__25600;
    wire N__25597;
    wire N__25594;
    wire N__25591;
    wire N__25588;
    wire N__25585;
    wire N__25582;
    wire N__25579;
    wire N__25578;
    wire N__25575;
    wire N__25572;
    wire N__25567;
    wire N__25564;
    wire N__25563;
    wire N__25560;
    wire N__25557;
    wire N__25552;
    wire N__25549;
    wire N__25548;
    wire N__25545;
    wire N__25542;
    wire N__25537;
    wire N__25534;
    wire N__25533;
    wire N__25530;
    wire N__25527;
    wire N__25522;
    wire N__25519;
    wire N__25518;
    wire N__25515;
    wire N__25512;
    wire N__25507;
    wire N__25504;
    wire N__25503;
    wire N__25500;
    wire N__25497;
    wire N__25492;
    wire N__25489;
    wire N__25486;
    wire N__25483;
    wire N__25480;
    wire N__25477;
    wire N__25474;
    wire N__25471;
    wire N__25468;
    wire N__25465;
    wire N__25464;
    wire N__25463;
    wire N__25460;
    wire N__25457;
    wire N__25454;
    wire N__25451;
    wire N__25444;
    wire N__25443;
    wire N__25440;
    wire N__25437;
    wire N__25432;
    wire N__25429;
    wire N__25428;
    wire N__25425;
    wire N__25424;
    wire N__25421;
    wire N__25418;
    wire N__25415;
    wire N__25412;
    wire N__25405;
    wire N__25402;
    wire N__25401;
    wire N__25398;
    wire N__25395;
    wire N__25392;
    wire N__25389;
    wire N__25386;
    wire N__25381;
    wire N__25378;
    wire N__25377;
    wire N__25374;
    wire N__25371;
    wire N__25366;
    wire N__25363;
    wire N__25362;
    wire N__25359;
    wire N__25356;
    wire N__25351;
    wire N__25348;
    wire N__25347;
    wire N__25344;
    wire N__25341;
    wire N__25336;
    wire N__25333;
    wire N__25332;
    wire N__25329;
    wire N__25326;
    wire N__25321;
    wire N__25318;
    wire N__25317;
    wire N__25314;
    wire N__25311;
    wire N__25306;
    wire N__25303;
    wire N__25302;
    wire N__25299;
    wire N__25296;
    wire N__25291;
    wire N__25288;
    wire N__25287;
    wire N__25286;
    wire N__25283;
    wire N__25278;
    wire N__25275;
    wire N__25270;
    wire N__25267;
    wire N__25266;
    wire N__25263;
    wire N__25260;
    wire N__25255;
    wire N__25252;
    wire N__25249;
    wire N__25248;
    wire N__25247;
    wire N__25244;
    wire N__25241;
    wire N__25238;
    wire N__25235;
    wire N__25232;
    wire N__25229;
    wire N__25222;
    wire N__25221;
    wire N__25218;
    wire N__25215;
    wire N__25210;
    wire N__25207;
    wire N__25204;
    wire N__25201;
    wire N__25198;
    wire N__25197;
    wire N__25194;
    wire N__25193;
    wire N__25190;
    wire N__25187;
    wire N__25184;
    wire N__25181;
    wire N__25174;
    wire N__25171;
    wire N__25168;
    wire N__25165;
    wire N__25162;
    wire N__25159;
    wire N__25156;
    wire N__25153;
    wire N__25150;
    wire N__25149;
    wire N__25148;
    wire N__25145;
    wire N__25140;
    wire N__25137;
    wire N__25132;
    wire N__25129;
    wire N__25126;
    wire N__25123;
    wire N__25122;
    wire N__25121;
    wire N__25118;
    wire N__25113;
    wire N__25110;
    wire N__25105;
    wire N__25102;
    wire N__25099;
    wire N__25096;
    wire N__25093;
    wire N__25090;
    wire N__25087;
    wire N__25084;
    wire N__25081;
    wire N__25078;
    wire N__25077;
    wire N__25076;
    wire N__25071;
    wire N__25068;
    wire N__25063;
    wire N__25060;
    wire N__25057;
    wire N__25054;
    wire N__25051;
    wire N__25048;
    wire N__25045;
    wire N__25042;
    wire N__25041;
    wire N__25038;
    wire N__25035;
    wire N__25032;
    wire N__25027;
    wire N__25024;
    wire N__25021;
    wire N__25018;
    wire N__25015;
    wire N__25012;
    wire N__25009;
    wire N__25008;
    wire N__25007;
    wire N__25004;
    wire N__25001;
    wire N__24998;
    wire N__24997;
    wire N__24990;
    wire N__24989;
    wire N__24986;
    wire N__24983;
    wire N__24978;
    wire N__24975;
    wire N__24972;
    wire N__24969;
    wire N__24966;
    wire N__24963;
    wire N__24958;
    wire N__24955;
    wire N__24952;
    wire N__24949;
    wire N__24946;
    wire N__24943;
    wire N__24940;
    wire N__24937;
    wire N__24934;
    wire N__24931;
    wire N__24928;
    wire N__24925;
    wire N__24922;
    wire N__24919;
    wire N__24916;
    wire N__24913;
    wire N__24910;
    wire N__24907;
    wire N__24904;
    wire N__24903;
    wire N__24900;
    wire N__24899;
    wire N__24896;
    wire N__24891;
    wire N__24886;
    wire N__24885;
    wire N__24882;
    wire N__24879;
    wire N__24874;
    wire N__24871;
    wire N__24870;
    wire N__24867;
    wire N__24864;
    wire N__24859;
    wire N__24856;
    wire N__24855;
    wire N__24850;
    wire N__24847;
    wire N__24844;
    wire N__24841;
    wire N__24838;
    wire N__24837;
    wire N__24834;
    wire N__24831;
    wire N__24828;
    wire N__24825;
    wire N__24820;
    wire N__24817;
    wire N__24814;
    wire N__24811;
    wire N__24808;
    wire N__24807;
    wire N__24804;
    wire N__24801;
    wire N__24796;
    wire N__24795;
    wire N__24792;
    wire N__24789;
    wire N__24784;
    wire N__24783;
    wire N__24780;
    wire N__24777;
    wire N__24774;
    wire N__24769;
    wire N__24768;
    wire N__24765;
    wire N__24762;
    wire N__24757;
    wire N__24756;
    wire N__24753;
    wire N__24750;
    wire N__24745;
    wire N__24744;
    wire N__24741;
    wire N__24738;
    wire N__24733;
    wire N__24730;
    wire N__24729;
    wire N__24726;
    wire N__24723;
    wire N__24718;
    wire N__24715;
    wire N__24712;
    wire N__24711;
    wire N__24708;
    wire N__24705;
    wire N__24700;
    wire N__24697;
    wire N__24694;
    wire N__24691;
    wire N__24690;
    wire N__24687;
    wire N__24684;
    wire N__24683;
    wire N__24678;
    wire N__24675;
    wire N__24672;
    wire N__24667;
    wire N__24666;
    wire N__24661;
    wire N__24658;
    wire N__24657;
    wire N__24654;
    wire N__24651;
    wire N__24646;
    wire N__24645;
    wire N__24644;
    wire N__24641;
    wire N__24638;
    wire N__24635;
    wire N__24632;
    wire N__24629;
    wire N__24626;
    wire N__24623;
    wire N__24616;
    wire N__24613;
    wire N__24612;
    wire N__24611;
    wire N__24608;
    wire N__24605;
    wire N__24602;
    wire N__24595;
    wire N__24592;
    wire N__24589;
    wire N__24586;
    wire N__24583;
    wire N__24580;
    wire N__24577;
    wire N__24574;
    wire N__24573;
    wire N__24570;
    wire N__24567;
    wire N__24562;
    wire N__24559;
    wire N__24558;
    wire N__24553;
    wire N__24550;
    wire N__24547;
    wire N__24544;
    wire N__24541;
    wire N__24538;
    wire N__24535;
    wire N__24532;
    wire N__24529;
    wire N__24526;
    wire N__24523;
    wire N__24520;
    wire N__24517;
    wire N__24514;
    wire N__24513;
    wire N__24510;
    wire N__24507;
    wire N__24504;
    wire N__24501;
    wire N__24498;
    wire N__24495;
    wire N__24492;
    wire N__24489;
    wire N__24486;
    wire N__24483;
    wire N__24480;
    wire N__24477;
    wire N__24474;
    wire N__24471;
    wire N__24468;
    wire N__24465;
    wire N__24462;
    wire N__24457;
    wire N__24454;
    wire N__24453;
    wire N__24450;
    wire N__24447;
    wire N__24446;
    wire N__24443;
    wire N__24438;
    wire N__24433;
    wire N__24432;
    wire N__24427;
    wire N__24424;
    wire N__24421;
    wire N__24420;
    wire N__24417;
    wire N__24414;
    wire N__24413;
    wire N__24410;
    wire N__24407;
    wire N__24404;
    wire N__24399;
    wire N__24394;
    wire N__24391;
    wire N__24388;
    wire N__24385;
    wire N__24382;
    wire N__24379;
    wire N__24376;
    wire N__24373;
    wire N__24370;
    wire N__24367;
    wire N__24364;
    wire N__24361;
    wire N__24358;
    wire N__24355;
    wire N__24352;
    wire N__24349;
    wire N__24346;
    wire N__24343;
    wire N__24342;
    wire N__24339;
    wire N__24338;
    wire N__24335;
    wire N__24332;
    wire N__24329;
    wire N__24326;
    wire N__24323;
    wire N__24320;
    wire N__24315;
    wire N__24310;
    wire N__24309;
    wire N__24306;
    wire N__24303;
    wire N__24300;
    wire N__24297;
    wire N__24292;
    wire N__24289;
    wire N__24286;
    wire N__24283;
    wire N__24280;
    wire N__24279;
    wire N__24276;
    wire N__24273;
    wire N__24268;
    wire N__24265;
    wire N__24262;
    wire N__24259;
    wire N__24256;
    wire N__24255;
    wire N__24252;
    wire N__24251;
    wire N__24248;
    wire N__24245;
    wire N__24242;
    wire N__24235;
    wire N__24234;
    wire N__24231;
    wire N__24230;
    wire N__24227;
    wire N__24224;
    wire N__24221;
    wire N__24214;
    wire N__24211;
    wire N__24208;
    wire N__24205;
    wire N__24202;
    wire N__24199;
    wire N__24196;
    wire N__24195;
    wire N__24194;
    wire N__24191;
    wire N__24188;
    wire N__24185;
    wire N__24182;
    wire N__24179;
    wire N__24176;
    wire N__24175;
    wire N__24172;
    wire N__24167;
    wire N__24166;
    wire N__24163;
    wire N__24160;
    wire N__24157;
    wire N__24154;
    wire N__24151;
    wire N__24142;
    wire N__24139;
    wire N__24138;
    wire N__24135;
    wire N__24132;
    wire N__24129;
    wire N__24128;
    wire N__24125;
    wire N__24122;
    wire N__24119;
    wire N__24112;
    wire N__24111;
    wire N__24110;
    wire N__24107;
    wire N__24102;
    wire N__24097;
    wire N__24094;
    wire N__24091;
    wire N__24090;
    wire N__24089;
    wire N__24086;
    wire N__24081;
    wire N__24076;
    wire N__24073;
    wire N__24072;
    wire N__24069;
    wire N__24066;
    wire N__24063;
    wire N__24060;
    wire N__24055;
    wire N__24052;
    wire N__24049;
    wire N__24046;
    wire N__24045;
    wire N__24044;
    wire N__24041;
    wire N__24036;
    wire N__24031;
    wire N__24030;
    wire N__24027;
    wire N__24024;
    wire N__24021;
    wire N__24020;
    wire N__24017;
    wire N__24014;
    wire N__24011;
    wire N__24004;
    wire N__24001;
    wire N__23998;
    wire N__23995;
    wire N__23992;
    wire N__23989;
    wire N__23986;
    wire N__23985;
    wire N__23982;
    wire N__23979;
    wire N__23976;
    wire N__23973;
    wire N__23968;
    wire N__23965;
    wire N__23962;
    wire N__23961;
    wire N__23960;
    wire N__23957;
    wire N__23954;
    wire N__23951;
    wire N__23946;
    wire N__23941;
    wire N__23938;
    wire N__23935;
    wire N__23932;
    wire N__23929;
    wire N__23926;
    wire N__23923;
    wire N__23920;
    wire N__23917;
    wire N__23914;
    wire N__23911;
    wire N__23908;
    wire N__23905;
    wire N__23902;
    wire N__23899;
    wire N__23896;
    wire N__23893;
    wire N__23890;
    wire N__23887;
    wire N__23884;
    wire N__23881;
    wire N__23878;
    wire N__23875;
    wire N__23874;
    wire N__23871;
    wire N__23868;
    wire N__23865;
    wire N__23862;
    wire N__23857;
    wire N__23856;
    wire N__23853;
    wire N__23852;
    wire N__23849;
    wire N__23846;
    wire N__23843;
    wire N__23840;
    wire N__23837;
    wire N__23830;
    wire N__23827;
    wire N__23824;
    wire N__23823;
    wire N__23820;
    wire N__23819;
    wire N__23816;
    wire N__23813;
    wire N__23810;
    wire N__23807;
    wire N__23806;
    wire N__23805;
    wire N__23800;
    wire N__23797;
    wire N__23792;
    wire N__23785;
    wire N__23782;
    wire N__23779;
    wire N__23778;
    wire N__23777;
    wire N__23774;
    wire N__23771;
    wire N__23768;
    wire N__23767;
    wire N__23764;
    wire N__23763;
    wire N__23760;
    wire N__23755;
    wire N__23752;
    wire N__23749;
    wire N__23744;
    wire N__23737;
    wire N__23734;
    wire N__23733;
    wire N__23732;
    wire N__23729;
    wire N__23724;
    wire N__23719;
    wire N__23718;
    wire N__23717;
    wire N__23714;
    wire N__23711;
    wire N__23708;
    wire N__23701;
    wire N__23698;
    wire N__23697;
    wire N__23694;
    wire N__23691;
    wire N__23688;
    wire N__23683;
    wire N__23682;
    wire N__23681;
    wire N__23680;
    wire N__23677;
    wire N__23674;
    wire N__23671;
    wire N__23668;
    wire N__23659;
    wire N__23656;
    wire N__23653;
    wire N__23650;
    wire N__23647;
    wire N__23646;
    wire N__23643;
    wire N__23640;
    wire N__23635;
    wire N__23632;
    wire N__23629;
    wire N__23628;
    wire N__23627;
    wire N__23624;
    wire N__23621;
    wire N__23618;
    wire N__23615;
    wire N__23612;
    wire N__23609;
    wire N__23606;
    wire N__23603;
    wire N__23596;
    wire N__23593;
    wire N__23590;
    wire N__23587;
    wire N__23584;
    wire N__23581;
    wire N__23578;
    wire N__23577;
    wire N__23574;
    wire N__23571;
    wire N__23568;
    wire N__23565;
    wire N__23560;
    wire N__23557;
    wire N__23554;
    wire N__23553;
    wire N__23550;
    wire N__23547;
    wire N__23542;
    wire N__23541;
    wire N__23538;
    wire N__23535;
    wire N__23532;
    wire N__23529;
    wire N__23524;
    wire N__23523;
    wire N__23520;
    wire N__23517;
    wire N__23514;
    wire N__23511;
    wire N__23508;
    wire N__23505;
    wire N__23500;
    wire N__23499;
    wire N__23496;
    wire N__23493;
    wire N__23490;
    wire N__23487;
    wire N__23482;
    wire N__23479;
    wire N__23478;
    wire N__23477;
    wire N__23474;
    wire N__23471;
    wire N__23468;
    wire N__23463;
    wire N__23458;
    wire N__23457;
    wire N__23454;
    wire N__23451;
    wire N__23450;
    wire N__23447;
    wire N__23444;
    wire N__23441;
    wire N__23436;
    wire N__23431;
    wire N__23428;
    wire N__23425;
    wire N__23422;
    wire N__23419;
    wire N__23416;
    wire N__23415;
    wire N__23412;
    wire N__23409;
    wire N__23404;
    wire N__23401;
    wire N__23398;
    wire N__23395;
    wire N__23392;
    wire N__23391;
    wire N__23388;
    wire N__23385;
    wire N__23382;
    wire N__23379;
    wire N__23374;
    wire N__23371;
    wire N__23368;
    wire N__23367;
    wire N__23364;
    wire N__23361;
    wire N__23358;
    wire N__23355;
    wire N__23350;
    wire N__23347;
    wire N__23344;
    wire N__23343;
    wire N__23340;
    wire N__23337;
    wire N__23334;
    wire N__23331;
    wire N__23326;
    wire N__23325;
    wire N__23322;
    wire N__23319;
    wire N__23316;
    wire N__23313;
    wire N__23308;
    wire N__23307;
    wire N__23304;
    wire N__23301;
    wire N__23298;
    wire N__23295;
    wire N__23290;
    wire N__23287;
    wire N__23286;
    wire N__23283;
    wire N__23280;
    wire N__23277;
    wire N__23274;
    wire N__23269;
    wire N__23266;
    wire N__23263;
    wire N__23260;
    wire N__23257;
    wire N__23254;
    wire N__23251;
    wire N__23248;
    wire N__23245;
    wire N__23242;
    wire N__23239;
    wire N__23236;
    wire N__23233;
    wire N__23232;
    wire N__23231;
    wire N__23230;
    wire N__23229;
    wire N__23226;
    wire N__23219;
    wire N__23216;
    wire N__23209;
    wire N__23206;
    wire N__23205;
    wire N__23202;
    wire N__23199;
    wire N__23194;
    wire N__23191;
    wire N__23188;
    wire N__23185;
    wire N__23182;
    wire N__23179;
    wire N__23176;
    wire N__23173;
    wire N__23172;
    wire N__23169;
    wire N__23166;
    wire N__23163;
    wire N__23160;
    wire N__23155;
    wire N__23152;
    wire N__23149;
    wire N__23146;
    wire N__23143;
    wire N__23140;
    wire N__23137;
    wire N__23134;
    wire N__23133;
    wire N__23130;
    wire N__23127;
    wire N__23122;
    wire N__23119;
    wire N__23118;
    wire N__23115;
    wire N__23112;
    wire N__23107;
    wire N__23104;
    wire N__23103;
    wire N__23100;
    wire N__23097;
    wire N__23094;
    wire N__23089;
    wire N__23086;
    wire N__23085;
    wire N__23082;
    wire N__23079;
    wire N__23074;
    wire N__23071;
    wire N__23070;
    wire N__23067;
    wire N__23064;
    wire N__23059;
    wire N__23056;
    wire N__23053;
    wire N__23052;
    wire N__23049;
    wire N__23046;
    wire N__23041;
    wire N__23038;
    wire N__23035;
    wire N__23032;
    wire N__23029;
    wire N__23026;
    wire N__23023;
    wire N__23020;
    wire N__23017;
    wire N__23014;
    wire N__23011;
    wire N__23008;
    wire N__23005;
    wire N__23002;
    wire N__22999;
    wire N__22998;
    wire N__22995;
    wire N__22994;
    wire N__22993;
    wire N__22988;
    wire N__22983;
    wire N__22982;
    wire N__22977;
    wire N__22974;
    wire N__22971;
    wire N__22968;
    wire N__22965;
    wire N__22962;
    wire N__22957;
    wire N__22954;
    wire N__22951;
    wire N__22948;
    wire N__22945;
    wire N__22942;
    wire N__22941;
    wire N__22938;
    wire N__22935;
    wire N__22930;
    wire N__22927;
    wire N__22926;
    wire N__22923;
    wire N__22920;
    wire N__22917;
    wire N__22912;
    wire N__22909;
    wire N__22906;
    wire N__22905;
    wire N__22900;
    wire N__22897;
    wire N__22896;
    wire N__22891;
    wire N__22888;
    wire N__22887;
    wire N__22882;
    wire N__22879;
    wire N__22876;
    wire N__22875;
    wire N__22872;
    wire N__22869;
    wire N__22864;
    wire N__22861;
    wire N__22858;
    wire N__22855;
    wire N__22852;
    wire N__22849;
    wire N__22846;
    wire N__22845;
    wire N__22842;
    wire N__22839;
    wire N__22838;
    wire N__22835;
    wire N__22830;
    wire N__22825;
    wire N__22822;
    wire N__22819;
    wire N__22818;
    wire N__22815;
    wire N__22812;
    wire N__22807;
    wire N__22804;
    wire N__22803;
    wire N__22800;
    wire N__22797;
    wire N__22796;
    wire N__22793;
    wire N__22788;
    wire N__22783;
    wire N__22782;
    wire N__22779;
    wire N__22776;
    wire N__22775;
    wire N__22768;
    wire N__22765;
    wire N__22762;
    wire N__22759;
    wire N__22756;
    wire N__22753;
    wire N__22750;
    wire N__22747;
    wire N__22744;
    wire N__22741;
    wire N__22740;
    wire N__22739;
    wire N__22734;
    wire N__22731;
    wire N__22726;
    wire N__22725;
    wire N__22724;
    wire N__22721;
    wire N__22716;
    wire N__22711;
    wire N__22708;
    wire N__22705;
    wire N__22704;
    wire N__22703;
    wire N__22700;
    wire N__22697;
    wire N__22694;
    wire N__22691;
    wire N__22688;
    wire N__22681;
    wire N__22678;
    wire N__22677;
    wire N__22674;
    wire N__22673;
    wire N__22670;
    wire N__22667;
    wire N__22664;
    wire N__22657;
    wire N__22656;
    wire N__22653;
    wire N__22652;
    wire N__22649;
    wire N__22646;
    wire N__22643;
    wire N__22640;
    wire N__22637;
    wire N__22634;
    wire N__22627;
    wire N__22626;
    wire N__22623;
    wire N__22620;
    wire N__22619;
    wire N__22614;
    wire N__22611;
    wire N__22606;
    wire N__22605;
    wire N__22600;
    wire N__22597;
    wire N__22596;
    wire N__22595;
    wire N__22592;
    wire N__22589;
    wire N__22586;
    wire N__22583;
    wire N__22580;
    wire N__22577;
    wire N__22570;
    wire N__22567;
    wire N__22566;
    wire N__22563;
    wire N__22560;
    wire N__22559;
    wire N__22556;
    wire N__22553;
    wire N__22550;
    wire N__22543;
    wire N__22540;
    wire N__22537;
    wire N__22534;
    wire N__22531;
    wire N__22528;
    wire N__22525;
    wire N__22522;
    wire N__22519;
    wire N__22518;
    wire N__22515;
    wire N__22512;
    wire N__22509;
    wire N__22506;
    wire N__22501;
    wire N__22498;
    wire N__22495;
    wire N__22492;
    wire N__22491;
    wire N__22490;
    wire N__22487;
    wire N__22484;
    wire N__22481;
    wire N__22478;
    wire N__22475;
    wire N__22468;
    wire N__22465;
    wire N__22462;
    wire N__22459;
    wire N__22456;
    wire N__22453;
    wire N__22452;
    wire N__22449;
    wire N__22446;
    wire N__22443;
    wire N__22440;
    wire N__22435;
    wire N__22432;
    wire N__22429;
    wire N__22426;
    wire N__22425;
    wire N__22424;
    wire N__22421;
    wire N__22416;
    wire N__22411;
    wire N__22410;
    wire N__22409;
    wire N__22408;
    wire N__22405;
    wire N__22404;
    wire N__22403;
    wire N__22402;
    wire N__22399;
    wire N__22396;
    wire N__22395;
    wire N__22394;
    wire N__22393;
    wire N__22390;
    wire N__22389;
    wire N__22388;
    wire N__22387;
    wire N__22384;
    wire N__22381;
    wire N__22378;
    wire N__22375;
    wire N__22362;
    wire N__22361;
    wire N__22360;
    wire N__22359;
    wire N__22356;
    wire N__22355;
    wire N__22354;
    wire N__22353;
    wire N__22352;
    wire N__22351;
    wire N__22350;
    wire N__22345;
    wire N__22342;
    wire N__22337;
    wire N__22334;
    wire N__22333;
    wire N__22330;
    wire N__22325;
    wire N__22324;
    wire N__22323;
    wire N__22316;
    wire N__22313;
    wire N__22310;
    wire N__22303;
    wire N__22294;
    wire N__22291;
    wire N__22286;
    wire N__22281;
    wire N__22278;
    wire N__22261;
    wire N__22260;
    wire N__22259;
    wire N__22258;
    wire N__22257;
    wire N__22256;
    wire N__22255;
    wire N__22254;
    wire N__22253;
    wire N__22252;
    wire N__22249;
    wire N__22248;
    wire N__22247;
    wire N__22246;
    wire N__22243;
    wire N__22240;
    wire N__22237;
    wire N__22224;
    wire N__22223;
    wire N__22222;
    wire N__22221;
    wire N__22220;
    wire N__22219;
    wire N__22212;
    wire N__22209;
    wire N__22204;
    wire N__22199;
    wire N__22196;
    wire N__22195;
    wire N__22194;
    wire N__22193;
    wire N__22192;
    wire N__22191;
    wire N__22190;
    wire N__22187;
    wire N__22182;
    wire N__22179;
    wire N__22176;
    wire N__22169;
    wire N__22166;
    wire N__22163;
    wire N__22158;
    wire N__22151;
    wire N__22132;
    wire N__22131;
    wire N__22130;
    wire N__22129;
    wire N__22128;
    wire N__22127;
    wire N__22126;
    wire N__22125;
    wire N__22124;
    wire N__22123;
    wire N__22122;
    wire N__22121;
    wire N__22120;
    wire N__22119;
    wire N__22118;
    wire N__22117;
    wire N__22116;
    wire N__22115;
    wire N__22114;
    wire N__22113;
    wire N__22110;
    wire N__22109;
    wire N__22106;
    wire N__22105;
    wire N__22104;
    wire N__22103;
    wire N__22102;
    wire N__22101;
    wire N__22100;
    wire N__22099;
    wire N__22096;
    wire N__22095;
    wire N__22094;
    wire N__22093;
    wire N__22088;
    wire N__22085;
    wire N__22076;
    wire N__22069;
    wire N__22064;
    wire N__22057;
    wire N__22044;
    wire N__22041;
    wire N__22038;
    wire N__22037;
    wire N__22036;
    wire N__22035;
    wire N__22034;
    wire N__22033;
    wire N__22032;
    wire N__22031;
    wire N__22030;
    wire N__22027;
    wire N__22026;
    wire N__22025;
    wire N__22018;
    wire N__22015;
    wire N__22008;
    wire N__21999;
    wire N__21992;
    wire N__21991;
    wire N__21990;
    wire N__21989;
    wire N__21984;
    wire N__21983;
    wire N__21968;
    wire N__21965;
    wire N__21962;
    wire N__21959;
    wire N__21956;
    wire N__21953;
    wire N__21944;
    wire N__21937;
    wire N__21934;
    wire N__21931;
    wire N__21910;
    wire N__21907;
    wire N__21904;
    wire N__21903;
    wire N__21900;
    wire N__21897;
    wire N__21892;
    wire N__21889;
    wire N__21886;
    wire N__21883;
    wire N__21880;
    wire N__21877;
    wire N__21874;
    wire N__21871;
    wire N__21868;
    wire N__21867;
    wire N__21864;
    wire N__21861;
    wire N__21856;
    wire N__21853;
    wire N__21852;
    wire N__21849;
    wire N__21846;
    wire N__21843;
    wire N__21840;
    wire N__21839;
    wire N__21834;
    wire N__21831;
    wire N__21828;
    wire N__21823;
    wire N__21820;
    wire N__21817;
    wire N__21814;
    wire N__21813;
    wire N__21810;
    wire N__21807;
    wire N__21802;
    wire N__21801;
    wire N__21798;
    wire N__21795;
    wire N__21794;
    wire N__21791;
    wire N__21786;
    wire N__21781;
    wire N__21778;
    wire N__21777;
    wire N__21776;
    wire N__21773;
    wire N__21770;
    wire N__21767;
    wire N__21760;
    wire N__21759;
    wire N__21756;
    wire N__21753;
    wire N__21752;
    wire N__21749;
    wire N__21746;
    wire N__21743;
    wire N__21736;
    wire N__21733;
    wire N__21732;
    wire N__21729;
    wire N__21726;
    wire N__21725;
    wire N__21722;
    wire N__21719;
    wire N__21716;
    wire N__21709;
    wire N__21706;
    wire N__21703;
    wire N__21700;
    wire N__21697;
    wire N__21696;
    wire N__21695;
    wire N__21692;
    wire N__21687;
    wire N__21684;
    wire N__21681;
    wire N__21676;
    wire N__21673;
    wire N__21672;
    wire N__21671;
    wire N__21668;
    wire N__21665;
    wire N__21662;
    wire N__21659;
    wire N__21656;
    wire N__21649;
    wire N__21646;
    wire N__21643;
    wire N__21640;
    wire N__21637;
    wire N__21634;
    wire N__21631;
    wire N__21628;
    wire N__21625;
    wire N__21622;
    wire N__21619;
    wire N__21616;
    wire N__21613;
    wire N__21610;
    wire N__21607;
    wire N__21604;
    wire N__21603;
    wire N__21600;
    wire N__21597;
    wire N__21594;
    wire N__21591;
    wire N__21586;
    wire N__21583;
    wire N__21580;
    wire N__21579;
    wire N__21576;
    wire N__21573;
    wire N__21568;
    wire N__21567;
    wire N__21564;
    wire N__21561;
    wire N__21558;
    wire N__21557;
    wire N__21554;
    wire N__21551;
    wire N__21548;
    wire N__21541;
    wire N__21540;
    wire N__21537;
    wire N__21534;
    wire N__21533;
    wire N__21530;
    wire N__21527;
    wire N__21524;
    wire N__21517;
    wire N__21514;
    wire N__21513;
    wire N__21510;
    wire N__21507;
    wire N__21502;
    wire N__21501;
    wire N__21496;
    wire N__21493;
    wire N__21490;
    wire N__21487;
    wire N__21484;
    wire N__21481;
    wire N__21478;
    wire N__21475;
    wire N__21474;
    wire N__21473;
    wire N__21470;
    wire N__21467;
    wire N__21464;
    wire N__21461;
    wire N__21458;
    wire N__21451;
    wire N__21448;
    wire N__21447;
    wire N__21446;
    wire N__21443;
    wire N__21440;
    wire N__21437;
    wire N__21434;
    wire N__21431;
    wire N__21428;
    wire N__21421;
    wire N__21420;
    wire N__21417;
    wire N__21414;
    wire N__21413;
    wire N__21406;
    wire N__21403;
    wire N__21400;
    wire N__21397;
    wire N__21394;
    wire N__21391;
    wire N__21388;
    wire N__21387;
    wire N__21386;
    wire N__21383;
    wire N__21378;
    wire N__21373;
    wire N__21370;
    wire N__21367;
    wire N__21366;
    wire N__21363;
    wire N__21360;
    wire N__21357;
    wire N__21354;
    wire N__21349;
    wire N__21346;
    wire N__21345;
    wire N__21342;
    wire N__21339;
    wire N__21338;
    wire N__21335;
    wire N__21332;
    wire N__21329;
    wire N__21322;
    wire N__21321;
    wire N__21318;
    wire N__21315;
    wire N__21314;
    wire N__21311;
    wire N__21308;
    wire N__21305;
    wire N__21298;
    wire N__21297;
    wire N__21294;
    wire N__21291;
    wire N__21290;
    wire N__21287;
    wire N__21282;
    wire N__21277;
    wire N__21276;
    wire N__21273;
    wire N__21270;
    wire N__21269;
    wire N__21266;
    wire N__21263;
    wire N__21260;
    wire N__21253;
    wire N__21252;
    wire N__21251;
    wire N__21246;
    wire N__21243;
    wire N__21238;
    wire N__21237;
    wire N__21234;
    wire N__21231;
    wire N__21230;
    wire N__21227;
    wire N__21224;
    wire N__21221;
    wire N__21214;
    wire N__21213;
    wire N__21210;
    wire N__21207;
    wire N__21202;
    wire N__21199;
    wire N__21196;
    wire N__21195;
    wire N__21190;
    wire N__21187;
    wire N__21186;
    wire N__21185;
    wire N__21184;
    wire N__21183;
    wire N__21182;
    wire N__21181;
    wire N__21170;
    wire N__21165;
    wire N__21160;
    wire N__21159;
    wire N__21158;
    wire N__21157;
    wire N__21156;
    wire N__21155;
    wire N__21154;
    wire N__21153;
    wire N__21152;
    wire N__21149;
    wire N__21146;
    wire N__21141;
    wire N__21134;
    wire N__21131;
    wire N__21128;
    wire N__21115;
    wire N__21114;
    wire N__21111;
    wire N__21108;
    wire N__21103;
    wire N__21100;
    wire N__21097;
    wire N__21096;
    wire N__21093;
    wire N__21090;
    wire N__21087;
    wire N__21084;
    wire N__21079;
    wire N__21076;
    wire N__21073;
    wire N__21070;
    wire N__21069;
    wire N__21066;
    wire N__21065;
    wire N__21062;
    wire N__21059;
    wire N__21056;
    wire N__21049;
    wire N__21046;
    wire N__21043;
    wire N__21042;
    wire N__21039;
    wire N__21038;
    wire N__21035;
    wire N__21032;
    wire N__21029;
    wire N__21022;
    wire N__21019;
    wire N__21016;
    wire N__21013;
    wire N__21010;
    wire N__21007;
    wire N__21004;
    wire N__21001;
    wire N__20998;
    wire N__20995;
    wire N__20994;
    wire N__20991;
    wire N__20988;
    wire N__20983;
    wire N__20980;
    wire N__20977;
    wire N__20974;
    wire N__20971;
    wire N__20970;
    wire N__20969;
    wire N__20968;
    wire N__20967;
    wire N__20966;
    wire N__20965;
    wire N__20964;
    wire N__20963;
    wire N__20960;
    wire N__20949;
    wire N__20946;
    wire N__20945;
    wire N__20944;
    wire N__20943;
    wire N__20942;
    wire N__20941;
    wire N__20940;
    wire N__20939;
    wire N__20938;
    wire N__20937;
    wire N__20936;
    wire N__20935;
    wire N__20934;
    wire N__20933;
    wire N__20932;
    wire N__20929;
    wire N__20928;
    wire N__20927;
    wire N__20926;
    wire N__20925;
    wire N__20924;
    wire N__20923;
    wire N__20920;
    wire N__20915;
    wire N__20914;
    wire N__20913;
    wire N__20910;
    wire N__20907;
    wire N__20898;
    wire N__20897;
    wire N__20896;
    wire N__20895;
    wire N__20894;
    wire N__20893;
    wire N__20890;
    wire N__20873;
    wire N__20870;
    wire N__20867;
    wire N__20856;
    wire N__20851;
    wire N__20846;
    wire N__20839;
    wire N__20828;
    wire N__20809;
    wire N__20806;
    wire N__20805;
    wire N__20800;
    wire N__20797;
    wire N__20794;
    wire N__20791;
    wire N__20790;
    wire N__20787;
    wire N__20784;
    wire N__20779;
    wire N__20776;
    wire N__20773;
    wire N__20770;
    wire N__20767;
    wire N__20764;
    wire N__20761;
    wire N__20758;
    wire N__20755;
    wire N__20752;
    wire N__20749;
    wire N__20746;
    wire N__20743;
    wire N__20740;
    wire N__20737;
    wire N__20734;
    wire N__20731;
    wire N__20730;
    wire N__20727;
    wire N__20724;
    wire N__20719;
    wire N__20716;
    wire N__20713;
    wire N__20710;
    wire N__20707;
    wire N__20704;
    wire N__20701;
    wire N__20698;
    wire N__20695;
    wire N__20692;
    wire N__20689;
    wire N__20686;
    wire N__20683;
    wire N__20680;
    wire N__20679;
    wire N__20676;
    wire N__20673;
    wire N__20668;
    wire N__20665;
    wire N__20662;
    wire N__20659;
    wire N__20656;
    wire N__20653;
    wire N__20650;
    wire N__20647;
    wire N__20644;
    wire N__20641;
    wire N__20640;
    wire N__20637;
    wire N__20634;
    wire N__20631;
    wire N__20628;
    wire N__20625;
    wire N__20620;
    wire N__20617;
    wire N__20616;
    wire N__20615;
    wire N__20614;
    wire N__20611;
    wire N__20606;
    wire N__20603;
    wire N__20596;
    wire N__20595;
    wire N__20592;
    wire N__20589;
    wire N__20588;
    wire N__20587;
    wire N__20586;
    wire N__20583;
    wire N__20576;
    wire N__20573;
    wire N__20566;
    wire N__20563;
    wire N__20562;
    wire N__20561;
    wire N__20558;
    wire N__20555;
    wire N__20552;
    wire N__20545;
    wire N__20544;
    wire N__20541;
    wire N__20540;
    wire N__20537;
    wire N__20534;
    wire N__20531;
    wire N__20524;
    wire N__20521;
    wire N__20520;
    wire N__20519;
    wire N__20518;
    wire N__20517;
    wire N__20514;
    wire N__20511;
    wire N__20508;
    wire N__20505;
    wire N__20502;
    wire N__20493;
    wire N__20490;
    wire N__20487;
    wire N__20482;
    wire N__20479;
    wire N__20476;
    wire N__20475;
    wire N__20472;
    wire N__20469;
    wire N__20466;
    wire N__20461;
    wire N__20458;
    wire N__20457;
    wire N__20454;
    wire N__20453;
    wire N__20450;
    wire N__20449;
    wire N__20446;
    wire N__20439;
    wire N__20436;
    wire N__20431;
    wire N__20430;
    wire N__20429;
    wire N__20426;
    wire N__20421;
    wire N__20418;
    wire N__20413;
    wire N__20410;
    wire N__20407;
    wire N__20404;
    wire N__20401;
    wire N__20398;
    wire N__20395;
    wire N__20392;
    wire N__20389;
    wire N__20386;
    wire N__20383;
    wire N__20380;
    wire N__20377;
    wire N__20374;
    wire N__20371;
    wire N__20368;
    wire N__20367;
    wire N__20364;
    wire N__20361;
    wire N__20358;
    wire N__20355;
    wire N__20352;
    wire N__20349;
    wire N__20346;
    wire N__20343;
    wire N__20340;
    wire N__20337;
    wire N__20334;
    wire N__20331;
    wire N__20328;
    wire N__20325;
    wire N__20322;
    wire N__20319;
    wire N__20316;
    wire N__20313;
    wire N__20310;
    wire N__20305;
    wire N__20304;
    wire N__20301;
    wire N__20300;
    wire N__20293;
    wire N__20290;
    wire N__20287;
    wire N__20284;
    wire N__20281;
    wire N__20280;
    wire N__20277;
    wire N__20274;
    wire N__20271;
    wire N__20268;
    wire N__20263;
    wire N__20260;
    wire N__20257;
    wire N__20254;
    wire N__20251;
    wire N__20248;
    wire N__20245;
    wire N__20244;
    wire N__20241;
    wire N__20238;
    wire N__20235;
    wire N__20232;
    wire N__20227;
    wire N__20224;
    wire N__20221;
    wire N__20218;
    wire N__20217;
    wire N__20214;
    wire N__20211;
    wire N__20208;
    wire N__20205;
    wire N__20200;
    wire N__20197;
    wire N__20194;
    wire N__20191;
    wire N__20190;
    wire N__20189;
    wire N__20186;
    wire N__20181;
    wire N__20176;
    wire N__20173;
    wire N__20170;
    wire N__20167;
    wire N__20164;
    wire N__20161;
    wire N__20158;
    wire N__20155;
    wire N__20152;
    wire N__20149;
    wire N__20146;
    wire N__20145;
    wire N__20144;
    wire N__20143;
    wire N__20142;
    wire N__20139;
    wire N__20136;
    wire N__20133;
    wire N__20130;
    wire N__20127;
    wire N__20120;
    wire N__20113;
    wire N__20110;
    wire N__20107;
    wire N__20104;
    wire N__20103;
    wire N__20102;
    wire N__20099;
    wire N__20098;
    wire N__20093;
    wire N__20088;
    wire N__20085;
    wire N__20082;
    wire N__20077;
    wire N__20074;
    wire N__20071;
    wire N__20070;
    wire N__20065;
    wire N__20062;
    wire N__20061;
    wire N__20056;
    wire N__20053;
    wire N__20052;
    wire N__20047;
    wire N__20044;
    wire N__20041;
    wire N__20038;
    wire N__20035;
    wire N__20034;
    wire N__20029;
    wire N__20026;
    wire N__20023;
    wire N__20022;
    wire N__20019;
    wire N__20016;
    wire N__20013;
    wire N__20010;
    wire N__20005;
    wire N__20002;
    wire N__19999;
    wire N__19996;
    wire N__19993;
    wire N__19992;
    wire N__19989;
    wire N__19986;
    wire N__19981;
    wire N__19980;
    wire N__19977;
    wire N__19974;
    wire N__19971;
    wire N__19966;
    wire N__19963;
    wire N__19960;
    wire N__19957;
    wire N__19954;
    wire N__19953;
    wire N__19950;
    wire N__19947;
    wire N__19942;
    wire N__19939;
    wire N__19936;
    wire N__19933;
    wire N__19930;
    wire N__19929;
    wire N__19928;
    wire N__19925;
    wire N__19922;
    wire N__19919;
    wire N__19912;
    wire N__19909;
    wire N__19906;
    wire N__19903;
    wire N__19900;
    wire N__19897;
    wire N__19894;
    wire N__19893;
    wire N__19892;
    wire N__19891;
    wire N__19890;
    wire N__19889;
    wire N__19888;
    wire N__19885;
    wire N__19872;
    wire N__19867;
    wire N__19864;
    wire N__19863;
    wire N__19860;
    wire N__19859;
    wire N__19854;
    wire N__19851;
    wire N__19848;
    wire N__19843;
    wire N__19840;
    wire N__19837;
    wire N__19834;
    wire N__19831;
    wire N__19828;
    wire N__19825;
    wire N__19822;
    wire N__19819;
    wire N__19816;
    wire N__19813;
    wire N__19812;
    wire N__19809;
    wire N__19806;
    wire N__19801;
    wire N__19798;
    wire N__19795;
    wire N__19792;
    wire N__19789;
    wire N__19786;
    wire N__19783;
    wire N__19780;
    wire N__19777;
    wire N__19774;
    wire N__19771;
    wire N__19768;
    wire N__19765;
    wire N__19762;
    wire N__19759;
    wire N__19758;
    wire N__19757;
    wire N__19756;
    wire N__19755;
    wire N__19752;
    wire N__19751;
    wire N__19750;
    wire N__19749;
    wire N__19746;
    wire N__19745;
    wire N__19744;
    wire N__19741;
    wire N__19738;
    wire N__19737;
    wire N__19736;
    wire N__19735;
    wire N__19734;
    wire N__19733;
    wire N__19732;
    wire N__19729;
    wire N__19726;
    wire N__19723;
    wire N__19720;
    wire N__19717;
    wire N__19712;
    wire N__19703;
    wire N__19692;
    wire N__19689;
    wire N__19674;
    wire N__19669;
    wire N__19666;
    wire N__19663;
    wire N__19660;
    wire N__19657;
    wire N__19654;
    wire N__19653;
    wire N__19652;
    wire N__19651;
    wire N__19648;
    wire N__19645;
    wire N__19642;
    wire N__19641;
    wire N__19640;
    wire N__19637;
    wire N__19626;
    wire N__19623;
    wire N__19618;
    wire N__19617;
    wire N__19616;
    wire N__19613;
    wire N__19610;
    wire N__19607;
    wire N__19600;
    wire N__19597;
    wire N__19596;
    wire N__19595;
    wire N__19592;
    wire N__19589;
    wire N__19586;
    wire N__19579;
    wire N__19578;
    wire N__19577;
    wire N__19576;
    wire N__19575;
    wire N__19574;
    wire N__19569;
    wire N__19568;
    wire N__19563;
    wire N__19562;
    wire N__19561;
    wire N__19560;
    wire N__19559;
    wire N__19558;
    wire N__19553;
    wire N__19552;
    wire N__19551;
    wire N__19550;
    wire N__19547;
    wire N__19544;
    wire N__19541;
    wire N__19530;
    wire N__19527;
    wire N__19520;
    wire N__19507;
    wire N__19506;
    wire N__19505;
    wire N__19500;
    wire N__19497;
    wire N__19492;
    wire N__19491;
    wire N__19488;
    wire N__19487;
    wire N__19484;
    wire N__19479;
    wire N__19474;
    wire N__19473;
    wire N__19472;
    wire N__19469;
    wire N__19468;
    wire N__19467;
    wire N__19466;
    wire N__19461;
    wire N__19460;
    wire N__19459;
    wire N__19458;
    wire N__19457;
    wire N__19448;
    wire N__19447;
    wire N__19444;
    wire N__19437;
    wire N__19434;
    wire N__19433;
    wire N__19432;
    wire N__19431;
    wire N__19430;
    wire N__19427;
    wire N__19424;
    wire N__19417;
    wire N__19410;
    wire N__19407;
    wire N__19396;
    wire N__19393;
    wire N__19390;
    wire N__19389;
    wire N__19386;
    wire N__19383;
    wire N__19378;
    wire N__19377;
    wire N__19376;
    wire N__19373;
    wire N__19370;
    wire N__19367;
    wire N__19360;
    wire N__19359;
    wire N__19356;
    wire N__19355;
    wire N__19348;
    wire N__19345;
    wire N__19344;
    wire N__19339;
    wire N__19336;
    wire N__19335;
    wire N__19330;
    wire N__19327;
    wire N__19326;
    wire N__19323;
    wire N__19318;
    wire N__19315;
    wire N__19314;
    wire N__19309;
    wire N__19306;
    wire N__19303;
    wire N__19302;
    wire N__19299;
    wire N__19294;
    wire N__19291;
    wire N__19290;
    wire N__19287;
    wire N__19286;
    wire N__19283;
    wire N__19280;
    wire N__19277;
    wire N__19270;
    wire N__19269;
    wire N__19268;
    wire N__19265;
    wire N__19262;
    wire N__19259;
    wire N__19256;
    wire N__19251;
    wire N__19246;
    wire N__19243;
    wire N__19240;
    wire N__19239;
    wire N__19238;
    wire N__19233;
    wire N__19230;
    wire N__19225;
    wire N__19224;
    wire N__19219;
    wire N__19216;
    wire N__19213;
    wire N__19210;
    wire N__19209;
    wire N__19208;
    wire N__19205;
    wire N__19202;
    wire N__19199;
    wire N__19192;
    wire N__19191;
    wire N__19190;
    wire N__19187;
    wire N__19182;
    wire N__19177;
    wire N__19176;
    wire N__19175;
    wire N__19172;
    wire N__19167;
    wire N__19162;
    wire N__19161;
    wire N__19158;
    wire N__19157;
    wire N__19154;
    wire N__19149;
    wire N__19144;
    wire N__19141;
    wire N__19140;
    wire N__19135;
    wire N__19134;
    wire N__19131;
    wire N__19128;
    wire N__19123;
    wire N__19122;
    wire N__19119;
    wire N__19116;
    wire N__19115;
    wire N__19112;
    wire N__19109;
    wire N__19106;
    wire N__19099;
    wire N__19096;
    wire N__19093;
    wire N__19090;
    wire N__19087;
    wire N__19084;
    wire N__19081;
    wire N__19078;
    wire N__19075;
    wire N__19072;
    wire N__19069;
    wire N__19066;
    wire N__19063;
    wire N__19060;
    wire N__19057;
    wire N__19054;
    wire N__19051;
    wire N__19048;
    wire N__19045;
    wire N__19042;
    wire N__19039;
    wire N__19036;
    wire N__19033;
    wire N__19030;
    wire N__19027;
    wire N__19024;
    wire N__19021;
    wire N__19018;
    wire N__19015;
    wire N__19012;
    wire N__19009;
    wire N__19006;
    wire N__19003;
    wire N__19000;
    wire N__18997;
    wire N__18994;
    wire N__18991;
    wire N__18988;
    wire N__18985;
    wire ICE_GPMO_2;
    wire VCCG0;
    wire INViac_raw_buf_vac_raw_buf_merged11WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged3WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged10WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged8WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged4WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged9WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged5WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged0WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged6WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged1WCLKN_net;
    wire ICE_SYSCLK;
    wire INViac_raw_buf_vac_raw_buf_merged7WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged2WCLKN_net;
    wire RTD_SCLK;
    wire \RTD.n8 ;
    wire RTD_CS;
    wire \RTD.n11673 ;
    wire n13279_cascade_;
    wire RTD_SDO;
    wire read_buf_0;
    wire read_buf_5;
    wire read_buf_12;
    wire read_buf_6;
    wire read_buf_7;
    wire read_buf_11;
    wire n11700_cascade_;
    wire read_buf_14;
    wire read_buf_15;
    wire read_buf_1;
    wire read_buf_13;
    wire read_buf_9;
    wire adress_1;
    wire adress_2;
    wire adress_3;
    wire adress_4;
    wire adress_5;
    wire read_buf_10;
    wire n14465;
    wire read_buf_8;
    wire read_buf_4;
    wire n13279;
    wire read_buf_2;
    wire read_buf_3;
    wire n11700;
    wire \RTD.n11726 ;
    wire \RTD.n15050 ;
    wire RTD_SDI;
    wire \RTD.n11704 ;
    wire \RTD.n33_cascade_ ;
    wire n1_adj_1575;
    wire \RTD.n16614 ;
    wire \RTD.n16614_cascade_ ;
    wire \RTD.n19482 ;
    wire \RTD.n19482_cascade_ ;
    wire \RTD.n7285_cascade_ ;
    wire \RTD.n21_cascade_ ;
    wire \RTD.n4 ;
    wire \RTD.n20969_cascade_ ;
    wire \RTD.n32 ;
    wire adress_6;
    wire \RTD.adress_7 ;
    wire adress_0;
    wire \RTD.n19855 ;
    wire \RTD.adress_7_N_1331_7_cascade_ ;
    wire RTD_DRDY;
    wire \RTD.n11_cascade_ ;
    wire \RTD.n19_cascade_ ;
    wire n13151;
    wire \RTD.n1_adj_1393 ;
    wire \RTD.adress_7_N_1331_7 ;
    wire \RTD.n16 ;
    wire \RTD.mode ;
    wire \RTD.n10 ;
    wire \RTD.cfg_buf_2 ;
    wire \RTD.cfg_buf_4 ;
    wire \RTD.cfg_buf_7 ;
    wire \RTD.n12 ;
    wire cfg_buf_1;
    wire buf_readRTD_7;
    wire n19_adj_1622_cascade_;
    wire buf_adcdata_vac_15;
    wire buf_data_iac_3;
    wire buf_data_iac_21;
    wire cmd_rdadctmp_28_adj_1415;
    wire buf_readRTD_5;
    wire n14_adj_1577;
    wire n20573_cascade_;
    wire VAC_CS;
    wire VAC_SCLK;
    wire buf_data_iac_8;
    wire data_index_9_N_212_7;
    wire \CLK_DDS.n9 ;
    wire \RTD.bit_cnt_1 ;
    wire \RTD.bit_cnt_0 ;
    wire \RTD.bit_cnt_2 ;
    wire \RTD.n17638 ;
    wire \RTD.bit_cnt_3 ;
    wire \RTD.n17638_cascade_ ;
    wire \RTD.n1_adj_1392 ;
    wire \RTD.n21063_cascade_ ;
    wire bit_cnt_1;
    wire bit_cnt_2;
    wire n8_adj_1409;
    wire \CLK_DDS.n16711 ;
    wire \RTD.n7285 ;
    wire \RTD.n11_adj_1394 ;
    wire \RTD.n21091 ;
    wire \RTD.n33 ;
    wire \RTD.n17676 ;
    wire \RTD.n7_adj_1395 ;
    wire \RTD.n11712 ;
    wire \RTD.cfg_tmp_1 ;
    wire \RTD.cfg_tmp_2 ;
    wire \RTD.cfg_tmp_3 ;
    wire \RTD.cfg_tmp_4 ;
    wire \RTD.cfg_tmp_5 ;
    wire \RTD.cfg_tmp_6 ;
    wire \RTD.cfg_tmp_7 ;
    wire \RTD.cfg_tmp_0 ;
    wire \RTD.adc_state_0 ;
    wire n18586_cascade_;
    wire cfg_buf_0;
    wire \RTD.n9 ;
    wire \RTD.n11 ;
    wire \RTD.n14 ;
    wire \RTD.n20722_cascade_ ;
    wire \RTD.n13198 ;
    wire \RTD.n13198_cascade_ ;
    wire \RTD.n14984 ;
    wire \RTD.cfg_buf_5 ;
    wire \RTD.n11_adj_1396 ;
    wire \RTD.cfg_buf_3 ;
    wire n18586;
    wire n13162;
    wire \RTD.cfg_buf_6 ;
    wire buf_readRTD_11;
    wire n22099_cascade_;
    wire n22102_cascade_;
    wire buf_adcdata_vac_19;
    wire n19_adj_1610_cascade_;
    wire buf_adcdata_iac_3;
    wire n22_adj_1611;
    wire cmd_rdadctmp_29_adj_1414;
    wire cmd_rdadctmp_10;
    wire cmd_rdadctmp_26_adj_1417;
    wire cmd_rdadctmp_27_adj_1416;
    wire cmd_rdadctmp_9;
    wire cmd_rdadctmp_23_adj_1420;
    wire buf_adcdata_vac_3;
    wire cmd_rdadctmp_8;
    wire cmd_rdadctmp_22_adj_1421;
    wire n19_adj_1487;
    wire buf_adcdata_vac_8;
    wire buf_readRTD_0;
    wire n19_adj_1479_cascade_;
    wire n23_adj_1512_cascade_;
    wire cmd_rdadctmp_6_adj_1437;
    wire cmd_rdadctmp_21_adj_1422;
    wire buf_adcdata_vac_13;
    wire cmd_rdadctmp_4_adj_1439;
    wire cmd_rdadctmp_5_adj_1438;
    wire buf_data_iac_14;
    wire cmd_rdadctmp_20;
    wire cmd_rdadctmp_21;
    wire cmd_rdadctmp_19;
    wire cmd_rdadctmp_18;
    wire buf_data_iac_11;
    wire cmd_rdadctmp_17;
    wire buf_adcdata_iac_9;
    wire DDS_MCLK1;
    wire DDS_CS1;
    wire DDS_SCK1;
    wire \RTD.adc_state_3 ;
    wire \RTD.adc_state_1 ;
    wire adc_state_2_adj_1474;
    wire \RTD.n20487 ;
    wire buf_data_iac_22;
    wire DDS_MOSI1;
    wire buf_adcdata_vac_21;
    wire buf_readRTD_8;
    wire n22183_cascade_;
    wire buf_data_iac_2;
    wire buf_readRTD_13;
    wire n22153;
    wire buf_adcdata_iac_2;
    wire n19_adj_1613_cascade_;
    wire n22_adj_1614;
    wire buf_readRTD_15;
    wire buf_adcdata_vac_2;
    wire buf_adcdata_vac_22;
    wire buf_adcdata_vac_14;
    wire buf_adcdata_vac_17;
    wire cmd_rdadctmp_30_adj_1413;
    wire cmd_rdadctmp_31_adj_1412;
    wire buf_adcdata_vac_16;
    wire cmd_rdadctmp_10_adj_1433;
    wire cmd_rdadctmp_11_adj_1432;
    wire cmd_rdadctmp_7_adj_1436;
    wire cmd_rdadctmp_8_adj_1435;
    wire cmd_rdadctmp_9_adj_1434;
    wire VAC_MISO;
    wire n21973;
    wire cmd_rdadctmp_17_adj_1426;
    wire cmd_rdadctmp_16_adj_1427;
    wire cmd_rdadctmp_0_adj_1443;
    wire cmd_rdadctmp_1_adj_1442;
    wire cmd_rdadctmp_2_adj_1441;
    wire cmd_rdadctmp_3_adj_1440;
    wire n20573;
    wire \ADC_VAC.n12556_cascade_ ;
    wire \ADC_VAC.n20667 ;
    wire \ADC_VAC.n20747_cascade_ ;
    wire \ADC_VAC.n20763_cascade_ ;
    wire \ADC_VAC.n21031_cascade_ ;
    wire \ADC_VAC.n20668 ;
    wire VAC_DRDY;
    wire \ADC_VAC.n17_cascade_ ;
    wire \ADC_VAC.n12 ;
    wire \ADC_VAC.bit_cnt_0 ;
    wire bfn_7_17_0_;
    wire \ADC_VAC.bit_cnt_1 ;
    wire \ADC_VAC.n19357 ;
    wire \ADC_VAC.bit_cnt_2 ;
    wire \ADC_VAC.n19358 ;
    wire \ADC_VAC.bit_cnt_3 ;
    wire \ADC_VAC.n19359 ;
    wire \ADC_VAC.bit_cnt_4 ;
    wire \ADC_VAC.n19360 ;
    wire \ADC_VAC.bit_cnt_5 ;
    wire \ADC_VAC.n19361 ;
    wire \ADC_VAC.bit_cnt_6 ;
    wire \ADC_VAC.n19362 ;
    wire \ADC_VAC.n19363 ;
    wire \ADC_VAC.bit_cnt_7 ;
    wire \ADC_VAC.n12556 ;
    wire \ADC_VAC.n14829 ;
    wire \ADC_IAC.n12459_cascade_ ;
    wire bfn_7_19_0_;
    wire \ADC_IAC.n19350 ;
    wire \ADC_IAC.n19351 ;
    wire \ADC_IAC.n19352 ;
    wire \ADC_IAC.n19353 ;
    wire \ADC_IAC.n19354 ;
    wire \ADC_IAC.n19355 ;
    wire \ADC_IAC.n19356 ;
    wire \ADC_IAC.n12459 ;
    wire \ADC_IAC.n14791 ;
    wire bit_cnt_0_adj_1449;
    wire bit_cnt_3;
    wire n21206;
    wire buf_adcdata_vdc_3;
    wire \CLK_DDS.n9_adj_1386 ;
    wire buf_adcdata_vdc_21;
    wire buf_adcdata_vdc_13;
    wire buf_adcdata_vdc_16;
    wire buf_adcdata_vdc_2;
    wire buf_adcdata_vdc_19;
    wire buf_adcdata_vdc_15;
    wire buf_adcdata_vdc_14;
    wire buf_adcdata_vdc_22;
    wire buf_adcdata_vdc_17;
    wire buf_adcdata_vdc_0;
    wire buf_adcdata_vac_0;
    wire buf_adcdata_iac_0;
    wire n19_adj_1477_cascade_;
    wire buf_readRTD_14;
    wire n22141;
    wire buf_readRTD_10;
    wire buf_adcdata_vdc_18;
    wire buf_adcdata_vac_18;
    wire n21931_cascade_;
    wire buf_cfgRTD_2;
    wire buf_cfgRTD_3;
    wire buf_cfgRTD_0;
    wire n14490_cascade_;
    wire buf_cfgRTD_1;
    wire buf_readRTD_9;
    wire n22165;
    wire buf_adcdata_iac_1;
    wire buf_data_iac_1;
    wire n22_adj_1618_cascade_;
    wire buf_data_iac_16;
    wire n20781_cascade_;
    wire buf_adcdata_vdc_1;
    wire buf_adcdata_vac_1;
    wire n19_adj_1617;
    wire n22171_cascade_;
    wire n20775;
    wire n20842;
    wire n20843;
    wire n22051_cascade_;
    wire n20828;
    wire n20814;
    wire cmd_rdadctmp_24_adj_1419;
    wire cmd_rdadctmp_25_adj_1418;
    wire n22039;
    wire n22042;
    wire buf_cfgRTD_7;
    wire cmd_rdadctmp_20_adj_1423;
    wire cmd_rdadctmp_18_adj_1425;
    wire buf_adcdata_vac_12;
    wire buf_adcdata_vdc_10;
    wire buf_adcdata_vac_10;
    wire cmd_rdadctmp_19_adj_1424;
    wire buf_data_iac_23;
    wire n26_adj_1511_cascade_;
    wire n20834_cascade_;
    wire n22057_cascade_;
    wire buf_data_iac_12;
    wire n22135;
    wire buf_adcdata_vac_23;
    wire buf_adcdata_vdc_23;
    wire n20831;
    wire cmd_rdadctmp_7;
    wire n16_adj_1507;
    wire cmd_rdadctmp_6;
    wire data_index_9_N_212_8;
    wire cmd_rdadctmp_22;
    wire n8_adj_1534;
    wire buf_adcdata_iac_8;
    wire cmd_rdadctmp_5;
    wire buf_adcdata_iac_22;
    wire cmd_rdadctmp_1;
    wire n20553;
    wire cmd_rdadctmp_29;
    wire cmd_rdadctmp_27;
    wire IAC_MISO;
    wire cmd_rdadctmp_0;
    wire cmd_rdadctmp_30;
    wire cmd_rdadctmp_4;
    wire cmd_rdadctmp_2;
    wire cmd_rdadctmp_3;
    wire IAC_CS;
    wire n14_adj_1581;
    wire \ADC_IAC.n20669 ;
    wire \ADC_IAC.bit_cnt_4 ;
    wire \ADC_IAC.bit_cnt_3 ;
    wire \ADC_IAC.bit_cnt_1 ;
    wire \ADC_IAC.bit_cnt_2 ;
    wire \ADC_IAC.bit_cnt_6 ;
    wire \ADC_IAC.bit_cnt_0 ;
    wire \ADC_IAC.n20753_cascade_ ;
    wire \ADC_IAC.bit_cnt_7 ;
    wire \ADC_IAC.bit_cnt_5 ;
    wire \ADC_IAC.n20765_cascade_ ;
    wire \ADC_IAC.n21007_cascade_ ;
    wire \ADC_IAC.n20670 ;
    wire IAC_DRDY;
    wire \ADC_IAC.n17_cascade_ ;
    wire \ADC_IAC.n12 ;
    wire \ADC_VDC.n20345 ;
    wire \ADC_VDC.cmd_rdadcbuf_0 ;
    wire bfn_9_5_0_;
    wire \ADC_VDC.cmd_rdadcbuf_1 ;
    wire \ADC_VDC.n19364 ;
    wire \ADC_VDC.cmd_rdadcbuf_2 ;
    wire \ADC_VDC.n19365 ;
    wire \ADC_VDC.cmd_rdadcbuf_3 ;
    wire \ADC_VDC.n19366 ;
    wire \ADC_VDC.cmd_rdadcbuf_4 ;
    wire \ADC_VDC.n19367 ;
    wire cmd_rdadctmp_5_adj_1467;
    wire \ADC_VDC.cmd_rdadcbuf_5 ;
    wire \ADC_VDC.n19368 ;
    wire cmd_rdadctmp_6_adj_1466;
    wire \ADC_VDC.cmd_rdadcbuf_6 ;
    wire \ADC_VDC.n19369 ;
    wire \ADC_VDC.cmd_rdadcbuf_7 ;
    wire \ADC_VDC.n19370 ;
    wire \ADC_VDC.n19371 ;
    wire \ADC_VDC.cmd_rdadcbuf_8 ;
    wire bfn_9_6_0_;
    wire cmd_rdadctmp_9_adj_1463;
    wire \ADC_VDC.cmd_rdadcbuf_9 ;
    wire \ADC_VDC.n19372 ;
    wire \ADC_VDC.cmd_rdadcbuf_10 ;
    wire \ADC_VDC.n19373 ;
    wire cmd_rdadcbuf_11;
    wire \ADC_VDC.n19374 ;
    wire cmd_rdadcbuf_12;
    wire \ADC_VDC.n19375 ;
    wire cmd_rdadctmp_13_adj_1459;
    wire cmd_rdadcbuf_13;
    wire \ADC_VDC.n19376 ;
    wire cmd_rdadctmp_14_adj_1458;
    wire cmd_rdadcbuf_14;
    wire \ADC_VDC.n19377 ;
    wire \ADC_VDC.n19378 ;
    wire \ADC_VDC.n19379 ;
    wire bfn_9_7_0_;
    wire \ADC_VDC.n19380 ;
    wire cmd_rdadctmp_18_adj_1454;
    wire \ADC_VDC.n19381 ;
    wire \ADC_VDC.n19382 ;
    wire \ADC_VDC.n19383 ;
    wire cmd_rdadctmp_21_adj_1451;
    wire cmd_rdadcbuf_21;
    wire \ADC_VDC.n19384 ;
    wire cmd_rdadctmp_22_adj_1450;
    wire \ADC_VDC.n19385 ;
    wire \ADC_VDC.cmd_rdadctmp_23 ;
    wire \ADC_VDC.n19386 ;
    wire \ADC_VDC.n19387 ;
    wire cmd_rdadcbuf_24;
    wire bfn_9_8_0_;
    wire cmd_rdadcbuf_25;
    wire \ADC_VDC.n19388 ;
    wire cmd_rdadcbuf_26;
    wire \ADC_VDC.n19389 ;
    wire cmd_rdadcbuf_27;
    wire \ADC_VDC.n19390 ;
    wire cmd_rdadcbuf_28;
    wire \ADC_VDC.n19391 ;
    wire cmd_rdadcbuf_29;
    wire \ADC_VDC.n19392 ;
    wire cmd_rdadcbuf_30;
    wire \ADC_VDC.n19393 ;
    wire cmd_rdadcbuf_31;
    wire \ADC_VDC.n19394 ;
    wire \ADC_VDC.n19395 ;
    wire cmd_rdadcbuf_32;
    wire bfn_9_9_0_;
    wire cmd_rdadcbuf_33;
    wire \ADC_VDC.n19396 ;
    wire \ADC_VDC.n19397 ;
    wire n20772;
    wire n21943;
    wire n21946_cascade_;
    wire n22060;
    wire n22054;
    wire n22015_cascade_;
    wire buf_data_iac_17;
    wire n20818_cascade_;
    wire n20871;
    wire n20820_cascade_;
    wire n21967;
    wire n21970;
    wire n22003_cascade_;
    wire n20624_cascade_;
    wire \SIG_DDS.n10_cascade_ ;
    wire buf_readRTD_12;
    wire n22006;
    wire n22027_cascade_;
    wire n22030;
    wire buf_adcdata_vac_20;
    wire buf_adcdata_vdc_20;
    wire n22207;
    wire n20801;
    wire buf_adcdata_iac_10;
    wire \SIG_DDS.bit_cnt_1 ;
    wire \SIG_DDS.bit_cnt_2 ;
    wire buf_adcdata_vac_11;
    wire cmd_rdadctmp_23;
    wire n8;
    wire n22117;
    wire buf_adcdata_iac_13;
    wire \SIG_DDS.bit_cnt_3 ;
    wire \SIG_DDS.n21292 ;
    wire VAC_OSR0;
    wire buf_adcdata_iac_19;
    wire n11417;
    wire buf_adcdata_iac_17;
    wire n22201_cascade_;
    wire n20805;
    wire cmd_rdadctmp_24;
    wire cmd_rdadctmp_31;
    wire buf_adcdata_iac_23;
    wire AC_ADC_SYNC;
    wire VAC_FLT1;
    wire IAC_SCLK;
    wire \ADC_VDC.n18394_cascade_ ;
    wire EIS_SYNCCLK;
    wire IAC_CLK;
    wire \ADC_VDC.n31_cascade_ ;
    wire \ADC_VDC.n21925_cascade_ ;
    wire \ADC_VDC.n18397 ;
    wire \ADC_VDC.n21928_cascade_ ;
    wire \ADC_VDC.n20514 ;
    wire \ADC_VDC.n6_cascade_ ;
    wire \ADC_VDC.n10519 ;
    wire n12853_cascade_;
    wire cmd_rdadctmp_0_adj_1472;
    wire cmd_rdadctmp_3_adj_1469;
    wire cmd_rdadctmp_4_adj_1468;
    wire \ADC_VDC.n12885 ;
    wire cmd_rdadctmp_7_adj_1465;
    wire cmd_rdadctmp_8_adj_1464;
    wire cmd_rdadctmp_17_adj_1455;
    wire cmd_rdadctmp_15_adj_1457;
    wire cmd_rdadctmp_16_adj_1456;
    wire cmd_rdadctmp_1_adj_1471;
    wire cmd_rdadctmp_2_adj_1470;
    wire cmd_rdadctmp_12_adj_1460;
    wire cmd_rdadctmp_10_adj_1462;
    wire cmd_rdadctmp_11_adj_1461;
    wire \ADC_VDC.n21673_cascade_ ;
    wire VDC_SCLK;
    wire cmd_rdadctmp_19_adj_1453;
    wire n12853;
    wire cmd_rdadctmp_20_adj_1452;
    wire cmd_rdadcbuf_23;
    wire buf_adcdata_vdc_12;
    wire cmd_rdadcbuf_22;
    wire buf_adcdata_vdc_11;
    wire cmd_rdadcbuf_15;
    wire cmd_rdadcbuf_20;
    wire cmd_rdadcbuf_19;
    wire buf_adcdata_vdc_8;
    wire cmd_rdadcbuf_18;
    wire cmd_rdadcbuf_17;
    wire cmd_rdadcbuf_16;
    wire \ADC_VDC.n18394 ;
    wire \ADC_VDC.cmd_rdadcbuf_35_N_1130_34 ;
    wire \ADC_VDC.n21106_cascade_ ;
    wire cmd_rdadcbuf_34;
    wire \ADC_VDC.n13020 ;
    wire \ADC_VDC.n21 ;
    wire \ADC_VDC.n19 ;
    wire buf_data_vac_16;
    wire buf_data_vac_23;
    wire buf_data_vac_22;
    wire buf_data_vac_21;
    wire buf_data_vac_20;
    wire buf_data_vac_19;
    wire buf_data_vac_18;
    wire buf_data_vac_17;
    wire n21143_cascade_;
    wire n12_cascade_;
    wire n12116;
    wire n12116_cascade_;
    wire n14756;
    wire n25_adj_1592_cascade_;
    wire n11944_cascade_;
    wire n11941_cascade_;
    wire n21919_cascade_;
    wire buf_data_iac_18;
    wire n20794_cascade_;
    wire n21922;
    wire n20796_cascade_;
    wire n21934;
    wire n22213_cascade_;
    wire n22216_cascade_;
    wire n20937;
    wire n20936;
    wire n21907_cascade_;
    wire buf_adcdata_iac_21;
    wire n22033_cascade_;
    wire n22036_cascade_;
    wire n22156;
    wire n21910;
    wire n20823_cascade_;
    wire n30_adj_1514_cascade_;
    wire n11941;
    wire n14735;
    wire \CLK_DDS.tmp_buf_10 ;
    wire \CLK_DDS.tmp_buf_11 ;
    wire \CLK_DDS.tmp_buf_12 ;
    wire \CLK_DDS.tmp_buf_13 ;
    wire \CLK_DDS.tmp_buf_14 ;
    wire \CLK_DDS.tmp_buf_9 ;
    wire \CLK_DDS.tmp_buf_8 ;
    wire buf_dds1_14;
    wire buf_dds1_12;
    wire buf_dds1_9;
    wire tmp_buf_15_adj_1448;
    wire \CLK_DDS.tmp_buf_0 ;
    wire \CLK_DDS.tmp_buf_1 ;
    wire \CLK_DDS.tmp_buf_2 ;
    wire \CLK_DDS.tmp_buf_3 ;
    wire \CLK_DDS.tmp_buf_4 ;
    wire \CLK_DDS.tmp_buf_5 ;
    wire \CLK_DDS.tmp_buf_6 ;
    wire \CLK_DDS.tmp_buf_7 ;
    wire buf_dds1_15;
    wire n22045;
    wire n22048;
    wire VAC_FLT0;
    wire n16_adj_1480;
    wire buf_dds1_0;
    wire buf_adcdata_iac_18;
    wire cmd_rdadctmp_25;
    wire cmd_rdadctmp_26;
    wire n23_adj_1513;
    wire cmd_rdadctmp_28;
    wire buf_adcdata_iac_20;
    wire IAC_FLT1;
    wire IAC_OSR1;
    wire IAC_FLT0;
    wire buf_adcdata_iac_16;
    wire buf_dds1_8;
    wire n22189_cascade_;
    wire n20769;
    wire n16_adj_1489;
    wire IAC_OSR0;
    wire bfn_11_3_0_;
    wire \ADC_VDC.genclk.n19410 ;
    wire \ADC_VDC.genclk.n19411 ;
    wire \ADC_VDC.genclk.n19412 ;
    wire \ADC_VDC.genclk.n19413 ;
    wire \ADC_VDC.genclk.n19414 ;
    wire \ADC_VDC.genclk.n19415 ;
    wire \ADC_VDC.genclk.n19416 ;
    wire \ADC_VDC.genclk.n19417 ;
    wire \INVADC_VDC.genclk.t0off_i0C_net ;
    wire bfn_11_4_0_;
    wire \ADC_VDC.genclk.n19418 ;
    wire \ADC_VDC.genclk.n19419 ;
    wire \ADC_VDC.genclk.n19420 ;
    wire \ADC_VDC.genclk.n19421 ;
    wire \ADC_VDC.genclk.n19422 ;
    wire \ADC_VDC.genclk.n19423 ;
    wire \ADC_VDC.genclk.n19424 ;
    wire \INVADC_VDC.genclk.t0off_i8C_net ;
    wire n13073;
    wire \ADC_VDC.n20618_cascade_ ;
    wire \ADC_VDC.n47 ;
    wire \ADC_VDC.n20702 ;
    wire \ADC_VDC.n20 ;
    wire dds_state_1_adj_1446;
    wire dds_state_2_adj_1445;
    wire trig_dds1;
    wire dds_state_0_adj_1447;
    wire \CLK_DDS.n12722 ;
    wire \ADC_VDC.avg_cnt_0 ;
    wire bfn_11_7_0_;
    wire \ADC_VDC.avg_cnt_1 ;
    wire \ADC_VDC.n19399 ;
    wire \ADC_VDC.avg_cnt_2 ;
    wire \ADC_VDC.n19400 ;
    wire \ADC_VDC.avg_cnt_3 ;
    wire \ADC_VDC.n19401 ;
    wire \ADC_VDC.avg_cnt_4 ;
    wire \ADC_VDC.n19402 ;
    wire \ADC_VDC.avg_cnt_5 ;
    wire \ADC_VDC.n19403 ;
    wire \ADC_VDC.avg_cnt_6 ;
    wire \ADC_VDC.n19404 ;
    wire \ADC_VDC.avg_cnt_7 ;
    wire \ADC_VDC.n19405 ;
    wire \ADC_VDC.n19406 ;
    wire \ADC_VDC.avg_cnt_8 ;
    wire bfn_11_8_0_;
    wire \ADC_VDC.avg_cnt_9 ;
    wire \ADC_VDC.n19407 ;
    wire \ADC_VDC.avg_cnt_10 ;
    wire \ADC_VDC.n19408 ;
    wire \ADC_VDC.n19409 ;
    wire \ADC_VDC.avg_cnt_11 ;
    wire \ADC_VDC.n13060 ;
    wire \ADC_VDC.n14900 ;
    wire n23_adj_1510_cascade_;
    wire n20833;
    wire buf_data_iac_20;
    wire n20810;
    wire THERMOSTAT;
    wire buf_control_7;
    wire n21050_cascade_;
    wire n11905;
    wire buf_cfgRTD_6;
    wire n11882_cascade_;
    wire comm_cmd_4;
    wire comm_cmd_6;
    wire comm_cmd_5;
    wire n8_adj_1522_cascade_;
    wire n12214_cascade_;
    wire buf_dds1_13;
    wire buf_dds1_11;
    wire n22075;
    wire n22078;
    wire buf_dds1_5;
    wire n7;
    wire n12214;
    wire n16539_cascade_;
    wire n17_adj_1601_cascade_;
    wire n16547;
    wire n16547_cascade_;
    wire n13_cascade_;
    wire INVeis_state_i0C_net;
    wire n19_adj_1482;
    wire buf_readRTD_6;
    wire n21937_cascade_;
    wire buf_adcdata_iac_14;
    wire n21940_cascade_;
    wire n30_adj_1490_cascade_;
    wire n26_adj_1495;
    wire n21109;
    wire n22111_cascade_;
    wire n22114;
    wire n8_adj_1536;
    wire AMPV_POW;
    wire DTRIG_N_910;
    wire adc_state_1;
    wire n10503;
    wire DTRIG_N_910_adj_1444;
    wire adc_state_1_adj_1410;
    wire VAC_OSR1;
    wire n4_adj_1473_cascade_;
    wire acadc_skipCount_13;
    wire buf_dds1_10;
    wire n22147;
    wire n22150;
    wire n20690_cascade_;
    wire acadc_trig;
    wire n20529;
    wire eis_end;
    wire INVacadc_trig_300C_net;
    wire eis_start;
    wire n17357;
    wire n11_adj_1620_cascade_;
    wire n11730;
    wire \ADC_VDC.genclk.t0off_6 ;
    wire \ADC_VDC.genclk.t0off_1 ;
    wire \ADC_VDC.genclk.t0off_4 ;
    wire \ADC_VDC.genclk.t0off_0 ;
    wire \ADC_VDC.genclk.n21169_cascade_ ;
    wire \ADC_VDC.genclk.t0off_12 ;
    wire \ADC_VDC.genclk.t0off_2 ;
    wire \ADC_VDC.genclk.t0off_7 ;
    wire \ADC_VDC.genclk.t0off_10 ;
    wire \ADC_VDC.genclk.n27 ;
    wire \ADC_VDC.genclk.t0off_13 ;
    wire \ADC_VDC.genclk.t0off_8 ;
    wire \ADC_VDC.genclk.t0off_5 ;
    wire \ADC_VDC.genclk.t0off_3 ;
    wire \ADC_VDC.genclk.n26 ;
    wire \ADC_VDC.genclk.t0off_14 ;
    wire \ADC_VDC.genclk.t0off_9 ;
    wire \ADC_VDC.genclk.t0off_15 ;
    wire \ADC_VDC.genclk.t0off_11 ;
    wire \ADC_VDC.genclk.n28 ;
    wire \ADC_VDC.genclk.n11721 ;
    wire \ADC_VDC.n10112_cascade_ ;
    wire \ADC_VDC.n12793 ;
    wire \ADC_VDC.n17 ;
    wire \ADC_VDC.n4 ;
    wire \ADC_VDC.n12 ;
    wire \ADC_VDC.n72 ;
    wire \ADC_VDC.n20710 ;
    wire \ADC_VDC.n20490_cascade_ ;
    wire \ADC_VDC.n11251_cascade_ ;
    wire \ADC_VDC.n20523_cascade_ ;
    wire \ADC_VDC.n21178 ;
    wire \ADC_VDC.n20490 ;
    wire \ADC_VDC.n21025 ;
    wire \ADC_VDC.n7_adj_1403 ;
    wire \ADC_VDC.n20712 ;
    wire \ADC_VDC.n11662 ;
    wire \ADC_VDC.n21028 ;
    wire comm_buf_0_7;
    wire \ADC_VDC.n10 ;
    wire \ADC_VDC.n15 ;
    wire \ADC_VDC.n19_adj_1405 ;
    wire wdtick_cnt_0;
    wire wdtick_cnt_1;
    wire wdtick_cnt_2;
    wire n14490;
    wire n11882;
    wire buf_data_iac_0;
    wire n22_adj_1476;
    wire buf_data_vac_8;
    wire buf_data_vac_15;
    wire buf_data_vac_14;
    wire buf_data_vac_13;
    wire buf_data_vac_12;
    wire buf_data_vac_11;
    wire buf_data_vac_10;
    wire buf_data_vac_9;
    wire n14_adj_1516;
    wire bfn_12_12_0_;
    wire n19335;
    wire n19336;
    wire n19337;
    wire n19338;
    wire n19339;
    wire data_idxvec_6;
    wire n19340;
    wire n19341;
    wire n19342;
    wire bfn_12_13_0_;
    wire data_idxvec_9;
    wire n19343;
    wire data_idxvec_10;
    wire n19344;
    wire n19345;
    wire data_idxvec_12;
    wire n19346;
    wire data_idxvec_13;
    wire n19347;
    wire data_idxvec_14;
    wire n19348;
    wire n19349;
    wire data_idxvec_15;
    wire data_idxvec_5;
    wire n26_adj_1486_cascade_;
    wire n22177_cascade_;
    wire n22120;
    wire n22180_cascade_;
    wire n30_adj_1485_cascade_;
    wire buf_data_iac_13;
    wire n21036;
    wire data_index_9_N_212_0;
    wire acadc_skipCount_8;
    wire n20_cascade_;
    wire n14_adj_1498;
    wire n18_adj_1587;
    wire n26_adj_1604_cascade_;
    wire n31;
    wire data_index_9_N_212_3;
    wire acadc_skipCount_5;
    wire n16_adj_1504;
    wire buf_dds1_1;
    wire acadc_skipCount_6;
    wire n17;
    wire acadc_dtrig_v;
    wire acadc_dtrig_i;
    wire iac_raw_buf_N_728_cascade_;
    wire n21997;
    wire buf_dds1_3;
    wire n20624;
    wire n12353_cascade_;
    wire n35;
    wire iac_raw_buf_N_726;
    wire eis_end_N_716;
    wire acadc_rst;
    wire buf_data_iac_15;
    wire buf_dds1_2;
    wire buf_adcdata_iac_15;
    wire n21961;
    wire n16_adj_1621_cascade_;
    wire buf_dds0_10;
    wire \SIG_DDS.tmp_buf_10 ;
    wire buf_dds0_9;
    wire \SIG_DDS.tmp_buf_9 ;
    wire buf_dds0_13;
    wire \SIG_DDS.tmp_buf_13 ;
    wire buf_dds0_14;
    wire buf_dds0_1;
    wire \SIG_DDS.tmp_buf_7 ;
    wire \SIG_DDS.tmp_buf_8 ;
    wire \comm_spi.n22629 ;
    wire \comm_spi.n22629_cascade_ ;
    wire \INVADC_VDC.genclk.t_clk_24C_net ;
    wire \comm_spi.n22632_cascade_ ;
    wire \comm_spi.imosi_cascade_ ;
    wire \comm_spi.imosi ;
    wire \comm_spi.n14599 ;
    wire \comm_spi.DOUT_7__N_738 ;
    wire \ADC_VDC.genclk.n21167 ;
    wire \ADC_VDC.n11_cascade_ ;
    wire \ADC_VDC.n17359 ;
    wire \ADC_VDC.bit_cnt_0 ;
    wire bfn_13_6_0_;
    wire \ADC_VDC.bit_cnt_1 ;
    wire \ADC_VDC.n19469 ;
    wire \ADC_VDC.n19470 ;
    wire \ADC_VDC.n19471 ;
    wire \ADC_VDC.bit_cnt_4 ;
    wire \ADC_VDC.n19472 ;
    wire \ADC_VDC.bit_cnt_5 ;
    wire \ADC_VDC.n19473 ;
    wire \ADC_VDC.bit_cnt_6 ;
    wire \ADC_VDC.n19474 ;
    wire \ADC_VDC.n19475 ;
    wire \ADC_VDC.bit_cnt_7 ;
    wire VDC_CLK;
    wire \ADC_VDC.n18381 ;
    wire \INVcomm_spi.imiso_83_12193_12194_setC_net ;
    wire buf_data_iac_6;
    wire \ADC_VDC.bit_cnt_3 ;
    wire \ADC_VDC.bit_cnt_2 ;
    wire \ADC_VDC.n6_adj_1404 ;
    wire \comm_spi.data_tx_7__N_762 ;
    wire n11727;
    wire \INVcomm_spi.bit_cnt_3767__i1C_net ;
    wire \comm_spi.bit_cnt_1 ;
    wire \comm_spi.bit_cnt_0 ;
    wire \comm_spi.bit_cnt_2 ;
    wire comm_buf_3_1;
    wire n21991_cascade_;
    wire n14763;
    wire comm_buf_3_3;
    wire n21979_cascade_;
    wire comm_buf_4_3;
    wire comm_buf_6_3;
    wire n4_adj_1567_cascade_;
    wire n20783_cascade_;
    wire n21982;
    wire comm_buf_3_5;
    wire n17331_cascade_;
    wire n20903_cascade_;
    wire n1_adj_1561_cascade_;
    wire comm_buf_6_6;
    wire comm_buf_3_6;
    wire n2_adj_1562;
    wire comm_buf_4_6;
    wire n21051;
    wire n4_adj_1563_cascade_;
    wire n22093;
    wire data_idxvec_2;
    wire n26_adj_1506_cascade_;
    wire buf_data_iac_10;
    wire n20816_cascade_;
    wire n20845;
    wire n22087_cascade_;
    wire n22090_cascade_;
    wire n19_adj_1505;
    wire buf_readRTD_2;
    wire n20846;
    wire n20815;
    wire n19;
    wire buf_readRTD_4;
    wire buf_adcdata_iac_12;
    wire n22081_cascade_;
    wire data_idxvec_4;
    wire n21261;
    wire n26_adj_1484_cascade_;
    wire n22159_cascade_;
    wire n22084;
    wire n22162_cascade_;
    wire n30_adj_1493_cascade_;
    wire data_idxvec_3;
    wire n21285;
    wire n26_adj_1502_cascade_;
    wire n22195_cascade_;
    wire acadc_skipCount_3;
    wire n22198_cascade_;
    wire n30_adj_1503_cascade_;
    wire n19_adj_1501;
    wire buf_readRTD_3;
    wire buf_adcdata_iac_11;
    wire n22009_cascade_;
    wire n16_adj_1500;
    wire n22012;
    wire acadc_skipcnt_0;
    wire bfn_13_16_0_;
    wire INVacadc_skipcnt_i0_i0C_net;
    wire n20757;
    wire n19311;
    wire n19311_THRU_CRY_0_THRU_CO;
    wire n19311_THRU_CRY_1_THRU_CO;
    wire n19311_THRU_CRY_2_THRU_CO;
    wire n19311_THRU_CRY_3_THRU_CO;
    wire n19311_THRU_CRY_4_THRU_CO;
    wire GNDG0;
    wire n19311_THRU_CRY_5_THRU_CO;
    wire n19311_THRU_CRY_6_THRU_CO;
    wire acadc_skipcnt_1;
    wire bfn_13_17_0_;
    wire n19312;
    wire acadc_skipcnt_3;
    wire n19313;
    wire acadc_skipcnt_4;
    wire n19314;
    wire acadc_skipcnt_5;
    wire n19315;
    wire acadc_skipcnt_6;
    wire n19316;
    wire n19317;
    wire acadc_skipcnt_8;
    wire n19318;
    wire n19319;
    wire INVacadc_skipcnt_i0_i1C_net;
    wire bfn_13_18_0_;
    wire n19320;
    wire n19321;
    wire n19322;
    wire acadc_skipcnt_13;
    wire n19323;
    wire n19324;
    wire n19325;
    wire INVacadc_skipcnt_i0_i9C_net;
    wire n11538;
    wire n14639;
    wire \SIG_DDS.tmp_buf_11 ;
    wire buf_dds0_12;
    wire \SIG_DDS.tmp_buf_12 ;
    wire \SIG_DDS.tmp_buf_1 ;
    wire \comm_spi.n22632 ;
    wire \comm_spi.n14600 ;
    wire \comm_spi.DOUT_7__N_739 ;
    wire \ADC_VDC.genclk.n21172_cascade_ ;
    wire \ADC_VDC.genclk.n21166 ;
    wire \ADC_VDC.genclk.n28_adj_1400 ;
    wire \ADC_VDC.genclk.n26_adj_1401 ;
    wire \ADC_VDC.genclk.n27_adj_1402 ;
    wire \comm_spi.n14586 ;
    wire \ADC_VDC.genclk.div_state_0 ;
    wire \ADC_VDC.genclk.div_state_1 ;
    wire \INVADC_VDC.genclk.div_state_i1C_net ;
    wire \ADC_VDC.genclk.n6 ;
    wire VDC_SDO;
    wire \ADC_VDC.adc_state_0 ;
    wire \ADC_VDC.n62 ;
    wire adc_state_2;
    wire adc_state_3;
    wire \ADC_VDC.n62_cascade_ ;
    wire \ADC_VDC.adc_state_1 ;
    wire \ADC_VDC.n11736 ;
    wire comm_buf_3_7;
    wire n1;
    wire n2_adj_1559_cascade_;
    wire comm_buf_4_7;
    wire comm_buf_6_7;
    wire n4_adj_1560;
    wire n21276_cascade_;
    wire n22105;
    wire comm_buf_3_2;
    wire n21985_cascade_;
    wire n21988_cascade_;
    wire comm_buf_3_0;
    wire n17304_cascade_;
    wire n20906_cascade_;
    wire comm_buf_4_2;
    wire comm_buf_6_2;
    wire n4_adj_1568_cascade_;
    wire n20786;
    wire n30_adj_1475;
    wire comm_buf_2_7;
    wire n30_adj_1595;
    wire comm_buf_2_6;
    wire n30_adj_1612;
    wire comm_buf_2_3;
    wire n30_adj_1615;
    wire comm_buf_2_2;
    wire n30_adj_1619;
    wire comm_buf_2_1;
    wire buf_data_vac_0;
    wire comm_buf_5_0;
    wire buf_data_vac_7;
    wire comm_buf_5_7;
    wire comm_rx_buf_6;
    wire buf_data_vac_6;
    wire comm_buf_5_6;
    wire buf_data_vac_5;
    wire comm_buf_5_5;
    wire comm_rx_buf_4;
    wire buf_data_vac_4;
    wire comm_rx_buf_3;
    wire buf_data_vac_3;
    wire comm_buf_5_3;
    wire comm_rx_buf_2;
    wire buf_data_vac_2;
    wire comm_buf_5_2;
    wire buf_data_vac_1;
    wire buf_readRTD_1;
    wire buf_adcdata_vdc_9;
    wire buf_adcdata_vac_9;
    wire n19_adj_1508;
    wire n20836;
    wire n22069_cascade_;
    wire n20837;
    wire data_idxvec_1;
    wire n26_adj_1509_cascade_;
    wire buf_data_iac_9;
    wire n20825;
    wire comm_rx_buf_1;
    wire n22072;
    wire data_idxvec_0;
    wire n21001;
    wire n26_cascade_;
    wire acadc_skipCount_0;
    wire n22021_cascade_;
    wire n22024;
    wire n21976;
    wire n30_adj_1478_cascade_;
    wire comm_rx_buf_0;
    wire cmd_rdadctmp_13_adj_1430;
    wire buf_dds1_4;
    wire n16;
    wire buf_dds1_6;
    wire n16_adj_1488;
    wire n20824;
    wire data_index_9_N_212_2;
    wire acadc_skipcnt_14;
    wire acadc_skipcnt_11;
    wire comm_buf_1_3;
    wire n8_adj_1543;
    wire acadc_skipcnt_2;
    wire acadc_skipcnt_7;
    wire acadc_skipCount_2;
    wire n23_adj_1586;
    wire n22_cascade_;
    wire n30_adj_1571;
    wire data_idxvec_7;
    wire acadc_skipCount_14;
    wire n8_adj_1545;
    wire acadc_skipcnt_9;
    wire acadc_skipcnt_15;
    wire acadc_skipCount_15;
    wire n24;
    wire acadc_skipCount_1;
    wire n9_adj_1407;
    wire n20949;
    wire n26_adj_1623;
    wire n21949_cascade_;
    wire acadc_skipCount_7;
    wire n21964;
    wire n21952_cascade_;
    wire acadc_skipCount_4;
    wire acadc_skipCount_9;
    wire comm_rx_buf_7;
    wire n30_adj_1624;
    wire n14742;
    wire buf_dds0_3;
    wire \SIG_DDS.tmp_buf_2 ;
    wire \SIG_DDS.tmp_buf_3 ;
    wire \SIG_DDS.tmp_buf_4 ;
    wire \SIG_DDS.tmp_buf_5 ;
    wire \SIG_DDS.tmp_buf_6 ;
    wire \ADC_VDC.genclk.t0on_0 ;
    wire bfn_15_3_0_;
    wire \ADC_VDC.genclk.t0on_1 ;
    wire \ADC_VDC.genclk.n19425 ;
    wire \ADC_VDC.genclk.t0on_2 ;
    wire \ADC_VDC.genclk.n19426 ;
    wire \ADC_VDC.genclk.t0on_3 ;
    wire \ADC_VDC.genclk.n19427 ;
    wire \ADC_VDC.genclk.t0on_4 ;
    wire \ADC_VDC.genclk.n19428 ;
    wire \ADC_VDC.genclk.t0on_5 ;
    wire \ADC_VDC.genclk.n19429 ;
    wire \ADC_VDC.genclk.t0on_6 ;
    wire \ADC_VDC.genclk.n19430 ;
    wire \ADC_VDC.genclk.t0on_7 ;
    wire \ADC_VDC.genclk.n19431 ;
    wire \ADC_VDC.genclk.n19432 ;
    wire \INVADC_VDC.genclk.t0on_i0C_net ;
    wire \ADC_VDC.genclk.t0on_8 ;
    wire bfn_15_4_0_;
    wire \ADC_VDC.genclk.t0on_9 ;
    wire \ADC_VDC.genclk.n19433 ;
    wire \ADC_VDC.genclk.t0on_10 ;
    wire \ADC_VDC.genclk.n19434 ;
    wire \ADC_VDC.genclk.t0on_11 ;
    wire \ADC_VDC.genclk.n19435 ;
    wire \ADC_VDC.genclk.t0on_12 ;
    wire \ADC_VDC.genclk.n19436 ;
    wire \ADC_VDC.genclk.t0on_13 ;
    wire \ADC_VDC.genclk.n19437 ;
    wire \ADC_VDC.genclk.t0on_14 ;
    wire \ADC_VDC.genclk.n19438 ;
    wire \ADC_VDC.genclk.n19439 ;
    wire \ADC_VDC.genclk.t0on_15 ;
    wire \INVADC_VDC.genclk.t0on_i8C_net ;
    wire \ADC_VDC.genclk.div_state_1__N_1266 ;
    wire \ADC_VDC.genclk.n14695 ;
    wire \comm_spi.n14585 ;
    wire \INVcomm_spi.MISO_48_12187_12188_setC_net ;
    wire comm_tx_buf_7;
    wire comm_tx_buf_2;
    wire \comm_spi.imosi_N_744 ;
    wire ICE_SPI_MOSI;
    wire \comm_spi.imosi_N_745 ;
    wire \comm_spi.n22644 ;
    wire \comm_spi.data_tx_7__N_778 ;
    wire \comm_spi.n14608 ;
    wire \comm_spi.data_tx_7__N_781 ;
    wire \comm_spi.n14607 ;
    wire \comm_spi.data_tx_7__N_763 ;
    wire comm_tx_buf_3;
    wire eis_state_0;
    wire n21067;
    wire n10508;
    wire n11839_cascade_;
    wire n9222;
    wire n9222_cascade_;
    wire n24_adj_1579_cascade_;
    wire n21079_cascade_;
    wire n12643;
    wire n16_adj_1570;
    wire n12080_cascade_;
    wire comm_buf_4_0;
    wire n22132;
    wire n12206;
    wire n12206_cascade_;
    wire n14770;
    wire comm_buf_6_0;
    wire comm_buf_2_0;
    wire n22129;
    wire buf_data_iac_5;
    wire n22_adj_1599_cascade_;
    wire n30_adj_1600_cascade_;
    wire comm_rx_buf_5;
    wire n12080;
    wire n14749;
    wire buf_adcdata_vdc_5;
    wire buf_adcdata_vac_5;
    wire n19_adj_1598;
    wire comm_buf_2_5;
    wire comm_buf_6_5;
    wire comm_buf_4_5;
    wire n22123_cascade_;
    wire n22126;
    wire n20602;
    wire SELIRNG0;
    wire n14_adj_1552;
    wire n14_adj_1552_cascade_;
    wire n14_adj_1550;
    wire n12254;
    wire n12007;
    wire n14_adj_1527;
    wire n14_adj_1529;
    wire req_data_cnt_5;
    wire req_data_cnt_4;
    wire req_data_cnt_1;
    wire n20_adj_1496;
    wire n18_adj_1553_cascade_;
    wire eis_stop;
    wire n29_cascade_;
    wire n16_adj_1609;
    wire n14_adj_1558;
    wire req_data_cnt_3;
    wire acadc_skipcnt_12;
    wire acadc_skipcnt_10;
    wire n21;
    wire n9_adj_1408_cascade_;
    wire cmd_rdadctmp_14_adj_1429;
    wire comm_buf_0_2;
    wire acadc_skipCount_10;
    wire n12391;
    wire n12367;
    wire n11324;
    wire n8780_cascade_;
    wire eis_state_1;
    wire buf_dds0_7;
    wire n8_adj_1541;
    wire n8_adj_1541_cascade_;
    wire data_index_9_N_212_4;
    wire data_count_0;
    wire bfn_15_17_0_;
    wire data_count_1;
    wire n19287;
    wire data_count_2;
    wire n19288;
    wire data_count_3;
    wire n19289;
    wire data_count_4;
    wire n19290;
    wire data_count_5;
    wire n19291;
    wire data_count_6;
    wire n19292;
    wire data_count_7;
    wire n19293;
    wire n19294;
    wire INVdata_count_i0_i0C_net;
    wire data_count_8;
    wire bfn_15_18_0_;
    wire n19295;
    wire data_count_9;
    wire INVdata_count_i0_i8C_net;
    wire \SIG_DDS.tmp_buf_14 ;
    wire buf_dds0_0;
    wire \SIG_DDS.tmp_buf_0 ;
    wire \SIG_DDS.n12700 ;
    wire comm_tx_buf_6;
    wire \comm_spi.data_tx_7__N_758 ;
    wire \comm_spi.n22623 ;
    wire \comm_spi.n14592 ;
    wire \comm_spi.n14593 ;
    wire \INVcomm_spi.imiso_83_12193_12194_resetC_net ;
    wire n17393;
    wire n30;
    wire comm_state_3_N_412_3_cascade_;
    wire n20700_cascade_;
    wire flagcntwd;
    wire n11411;
    wire n20081;
    wire n11333;
    wire comm_buf_0_6;
    wire n28;
    wire n27;
    wire n26_adj_1625_cascade_;
    wire n25_adj_1616;
    wire n19553_cascade_;
    wire n22_adj_1594;
    wire n10_adj_1582;
    wire clk_cnt_1;
    wire clk_cnt_0;
    wire clk_RTD;
    wire TEST_LED;
    wire buf_adcdata_vdc_6;
    wire buf_adcdata_vac_6;
    wire n19_adj_1593;
    wire n21071;
    wire n20_adj_1607;
    wire comm_buf_5_4;
    wire comm_buf_4_4;
    wire data_idxvec_8;
    wire n20779;
    wire n12415_cascade_;
    wire buf_cfgRTD_5;
    wire comm_buf_1_0;
    wire n14_adj_1528;
    wire n14_adj_1525;
    wire n20850;
    wire n30_adj_1520;
    wire n14_adj_1524;
    wire req_data_cnt_0;
    wire req_data_cnt_6;
    wire n17_adj_1554;
    wire req_data_cnt_15;
    wire req_data_cnt_9;
    wire n20613;
    wire req_data_cnt_2;
    wire req_data_cnt_7;
    wire n14_adj_1548;
    wire n22_adj_1492;
    wire n21_adj_1494_cascade_;
    wire n24_adj_1530;
    wire n30_adj_1597;
    wire n14_adj_1549;
    wire buf_cfgRTD_4;
    wire n12415;
    wire n14_adj_1551;
    wire req_data_cnt_10;
    wire req_data_cnt_8;
    wire n19_adj_1499;
    wire bfn_16_15_0_;
    wire n19326;
    wire data_index_2;
    wire n7_adj_1544;
    wire n19327;
    wire data_index_3;
    wire n7_adj_1542;
    wire n19328;
    wire data_index_4;
    wire n7_adj_1540;
    wire n19329;
    wire n19330;
    wire n19331;
    wire data_index_7;
    wire n7_adj_1535;
    wire n19332;
    wire n19333;
    wire data_index_8;
    wire n7_adj_1533;
    wire bfn_16_16_0_;
    wire n10579;
    wire n19334;
    wire n17338_cascade_;
    wire data_index_9_N_212_5;
    wire n7_adj_1515;
    wire n17314;
    wire data_index_0;
    wire comm_buf_1_2;
    wire buf_dds0_2;
    wire data_index_9;
    wire buf_dds0_4;
    wire n8_adj_1538_cascade_;
    wire data_index_6;
    wire buf_dds0_6;
    wire comm_buf_1_7;
    wire buf_dds1_7;
    wire comm_buf_0_0;
    wire buf_dds0_8;
    wire comm_buf_1_1;
    wire data_index_1;
    wire n8780;
    wire n8_adj_1547;
    wire n8_adj_1547_cascade_;
    wire n7_adj_1546;
    wire data_index_9_N_212_1;
    wire buf_dds0_11;
    wire buf_dds0_5;
    wire n8_adj_1532;
    wire n7_adj_1531;
    wire data_index_9_N_212_9;
    wire tmp_buf_15;
    wire DDS_MOSI;
    wire comm_buf_0_1;
    wire DDS_RNG_0;
    wire n8_adj_1538;
    wire n7_adj_1537;
    wire data_index_9_N_212_6;
    wire n11901;
    wire comm_buf_0_3;
    wire n14869;
    wire bit_cnt_0;
    wire \comm_spi.n14624 ;
    wire \comm_spi.data_tx_7__N_769 ;
    wire \comm_spi.n22626 ;
    wire \comm_spi.n22626_cascade_ ;
    wire \comm_spi.n14589 ;
    wire ICE_SPI_MISO;
    wire \comm_spi.n22635 ;
    wire \comm_spi.n14623 ;
    wire \comm_spi.data_tx_7__N_759 ;
    wire \comm_spi.n14596 ;
    wire \comm_spi.n14595 ;
    wire \comm_spi.n14588 ;
    wire \comm_spi.n14590 ;
    wire \INVcomm_spi.MISO_48_12187_12188_resetC_net ;
    wire \comm_spi.data_tx_7__N_766 ;
    wire n20931;
    wire n21913_cascade_;
    wire n21916;
    wire n1252_cascade_;
    wire n2;
    wire n21088_cascade_;
    wire n14_adj_1497;
    wire comm_state_3_N_412_3;
    wire n1252;
    wire n8_adj_1555;
    wire n2342_cascade_;
    wire comm_state_3_N_428_2;
    wire n15_adj_1602_cascade_;
    wire n20571;
    wire n20641_cascade_;
    wire n12_adj_1603;
    wire n7_adj_1588;
    wire secclk_cnt_0;
    wire bfn_17_9_0_;
    wire secclk_cnt_1;
    wire n19447;
    wire secclk_cnt_2;
    wire n19448;
    wire secclk_cnt_3;
    wire n19449;
    wire secclk_cnt_4;
    wire n19450;
    wire secclk_cnt_5;
    wire n19451;
    wire secclk_cnt_6;
    wire n19452;
    wire secclk_cnt_7;
    wire n19453;
    wire n19454;
    wire secclk_cnt_8;
    wire bfn_17_10_0_;
    wire secclk_cnt_9;
    wire n19455;
    wire secclk_cnt_10;
    wire n19456;
    wire secclk_cnt_11;
    wire n19457;
    wire n19458;
    wire secclk_cnt_13;
    wire n19459;
    wire secclk_cnt_14;
    wire n19460;
    wire secclk_cnt_15;
    wire n19461;
    wire n19462;
    wire secclk_cnt_16;
    wire bfn_17_11_0_;
    wire secclk_cnt_17;
    wire n19463;
    wire secclk_cnt_18;
    wire n19464;
    wire n19465;
    wire secclk_cnt_20;
    wire n19466;
    wire n19467;
    wire n19468;
    wire n14700;
    wire comm_buf_0_5;
    wire n14_adj_1556;
    wire VDC_RNG0;
    wire acadc_skipCount_12;
    wire req_data_cnt_13;
    wire n21022;
    wire n21049;
    wire comm_length_2;
    wire n21955_cascade_;
    wire n21958;
    wire n21024;
    wire buf_data_iac_19;
    wire n20950;
    wire data_idxvec_11;
    wire n26_adj_1519;
    wire SELIRNG1;
    wire acadc_skipCount_11;
    wire n23_adj_1518;
    wire comm_length_0;
    wire n11846;
    wire n14652;
    wire n10553;
    wire n20622;
    wire n12381;
    wire req_data_cnt_11;
    wire req_data_cnt_14;
    wire n23_adj_1491;
    wire cmd_rdadctmp_15_adj_1428;
    wire cmd_rdadctmp_15;
    wire cmd_rdadctmp_16;
    wire n17338;
    wire n17336;
    wire data_index_5;
    wire n16708;
    wire n20626;
    wire n11805;
    wire n14_adj_1523;
    wire n12353;
    wire buf_dds0_15;
    wire n9;
    wire \SIG_DDS.n9 ;
    wire \comm_spi.n14620 ;
    wire \comm_spi.data_tx_7__N_772 ;
    wire \comm_spi.n22638 ;
    wire \comm_spi.n14619 ;
    wire \comm_spi.n14615 ;
    wire \comm_spi.data_tx_7__N_761 ;
    wire \comm_spi.n22641 ;
    wire \comm_spi.n14611 ;
    wire \comm_spi.n14612 ;
    wire \comm_spi.n14616 ;
    wire n20641;
    wire n17656;
    wire n21162;
    wire n17658_cascade_;
    wire n20653;
    wire n12220_cascade_;
    wire n4_adj_1483_cascade_;
    wire n12205;
    wire n4;
    wire n20510_cascade_;
    wire n3;
    wire n20534;
    wire n11810;
    wire n11810_cascade_;
    wire n20650;
    wire n20672_cascade_;
    wire n20510;
    wire n20585;
    wire n11824;
    wire \comm_spi.bit_cnt_3 ;
    wire \comm_spi.n16858 ;
    wire \INVcomm_spi.data_valid_85C_net ;
    wire n21087;
    wire n4_adj_1566;
    wire n22063_cascade_;
    wire comm_buf_6_4;
    wire n21081;
    wire comm_buf_0_4;
    wire comm_buf_1_4;
    wire n1_adj_1564;
    wire n18824_cascade_;
    wire n20507;
    wire comm_buf_2_4;
    wire comm_buf_3_4;
    wire n2_adj_1565;
    wire comm_buf_5_1;
    wire comm_buf_4_1;
    wire n4_adj_1569_cascade_;
    wire comm_buf_6_1;
    wire n20792_cascade_;
    wire n21994;
    wire n12322;
    wire n14784;
    wire n21069;
    wire iac_raw_buf_N_728;
    wire data_cntvec_0;
    wire bfn_18_12_0_;
    wire data_cntvec_1;
    wire n19296;
    wire data_cntvec_2;
    wire n19297;
    wire data_cntvec_3;
    wire n19298;
    wire data_cntvec_4;
    wire n19299;
    wire data_cntvec_5;
    wire n19300;
    wire data_cntvec_6;
    wire n19301;
    wire data_cntvec_7;
    wire n19302;
    wire n19303;
    wire INVdata_cntvec_i0_i0C_net;
    wire data_cntvec_8;
    wire bfn_18_13_0_;
    wire data_cntvec_9;
    wire n19304;
    wire data_cntvec_10;
    wire n19305;
    wire data_cntvec_11;
    wire n19306;
    wire data_cntvec_12;
    wire n19307;
    wire data_cntvec_13;
    wire n19308;
    wire data_cntvec_14;
    wire n19309;
    wire n19310;
    wire data_cntvec_15;
    wire INVdata_cntvec_i0_i8C_net;
    wire n13443;
    wire n14632;
    wire buf_adcdata_iac_6;
    wire n20540;
    wire adc_state_0_adj_1411;
    wire cmd_rdadctmp_12_adj_1431;
    wire buf_adcdata_vac_7;
    wire buf_adcdata_vdc_7;
    wire buf_adcdata_iac_7;
    wire n19_adj_1589_cascade_;
    wire comm_cmd_2;
    wire buf_data_iac_7;
    wire n22_adj_1590_cascade_;
    wire n30_adj_1591;
    wire buf_adcdata_iac_5;
    wire cmd_rdadctmp_11;
    wire n20543;
    wire buf_adcdata_iac_4;
    wire cmd_rdadctmp_14;
    wire \comm_spi.n14581 ;
    wire \comm_spi.iclk_N_754 ;
    wire comm_tx_buf_5;
    wire \comm_spi.data_tx_7__N_760 ;
    wire ICE_GPMI_0;
    wire n11406;
    wire n12220;
    wire n10_adj_1572_cascade_;
    wire n20643;
    wire n4_adj_1596;
    wire n2342;
    wire n11836;
    wire n14722;
    wire \comm_spi.n22647 ;
    wire comm_buf_1_5;
    wire n14_adj_1557;
    wire comm_index_2;
    wire n18824;
    wire n20563_cascade_;
    wire n20627;
    wire n12_adj_1539_cascade_;
    wire n20556;
    wire n12164;
    wire ICE_SPI_CE0;
    wire comm_data_vld;
    wire n23_adj_1574;
    wire n21_adj_1573_cascade_;
    wire n18;
    wire comm_index_1;
    wire comm_length_1;
    wire n4_adj_1576;
    wire comm_cmd_7;
    wire n5_cascade_;
    wire n20863;
    wire n14514;
    wire n21658_cascade_;
    wire n9273;
    wire n20865_cascade_;
    wire n20536;
    wire n10540;
    wire comm_index_0;
    wire n20563;
    wire n12_adj_1585;
    wire comm_buf_1_6;
    wire n14_adj_1526;
    wire buf_adcdata_vdc_4;
    wire buf_adcdata_vac_4;
    wire n19_adj_1605;
    wire comm_state_2;
    wire n20734;
    wire adc_state_0;
    wire cmd_rdadctmp_12;
    wire n12542;
    wire cmd_rdadctmp_13;
    wire buf_control_0;
    wire wdtick_flag;
    wire CONT_SD;
    wire trig_dds0;
    wire \comm_spi.n14582 ;
    wire ICE_SPI_SCLK;
    wire \comm_spi.iclk_N_755 ;
    wire \comm_spi.data_tx_7__N_765 ;
    wire CONSTANT_ONE_NET;
    wire \comm_spi.data_tx_7__N_787 ;
    wire \comm_spi.n14604 ;
    wire \comm_spi.n14578 ;
    wire \comm_spi.n14577 ;
    wire \comm_spi.n14603 ;
    wire \comm_spi.iclk ;
    wire comm_tx_buf_0;
    wire \comm_spi.n22650 ;
    wire \comm_spi.data_tx_7__N_764 ;
    wire comm_tx_buf_1;
    wire \comm_spi.data_tx_7__N_784 ;
    wire comm_tx_buf_4;
    wire \comm_spi.data_tx_7__N_775 ;
    wire n20502_cascade_;
    wire n12_adj_1583;
    wire n20502;
    wire INVdds0_mclk_294C_net;
    wire secclk_cnt_19;
    wire secclk_cnt_21;
    wire secclk_cnt_12;
    wire secclk_cnt_22;
    wire n14_adj_1578;
    wire comm_cmd_1;
    wire comm_cmd_0;
    wire n23_adj_1517;
    wire req_data_cnt_12;
    wire n20809;
    wire n17415;
    wire buf_data_iac_4;
    wire comm_cmd_3;
    wire n22_adj_1606;
    wire n30_adj_1608;
    wire clk_16MHz;
    wire dds0_mclk;
    wire buf_control_6;
    wire DDS_MCLK;
    wire DDS_SCK;
    wire dds_state_2;
    wire dds_state_0;
    wire dds_state_1;
    wire DDS_CS;
    wire \SIG_DDS.n9_adj_1385 ;
    wire comm_clear;
    wire clk_32MHz;
    wire comm_state_3;
    wire comm_state_1;
    wire comm_state_0;
    wire n11347;
    wire dds0_mclkcnt_0;
    wire bfn_22_11_0_;
    wire dds0_mclkcnt_1;
    wire n19440;
    wire dds0_mclkcnt_2;
    wire n19441;
    wire dds0_mclkcnt_3;
    wire n19442;
    wire dds0_mclkcnt_4;
    wire n19443;
    wire dds0_mclkcnt_5;
    wire n19444;
    wire n10;
    wire dds0_mclkcnt_6;
    wire n19445;
    wire n19446;
    wire dds0_mclkcnt_7;
    wire INVdds0_mclkcnt_i7_3772__i0C_net;
    wire _gnd_net_;

    defparam \pll_main.zim_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \pll_main.zim_pll_inst .TEST_MODE=1'b0;
    defparam \pll_main.zim_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \pll_main.zim_pll_inst .PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam \pll_main.zim_pll_inst .PLLOUT_SELECT_PORTA="GENCLK";
    defparam \pll_main.zim_pll_inst .FILTER_RANGE=3'b011;
    defparam \pll_main.zim_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \pll_main.zim_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \pll_main.zim_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \pll_main.zim_pll_inst .ENABLE_ICEGATE_PORTB=1'b0;
    defparam \pll_main.zim_pll_inst .ENABLE_ICEGATE_PORTA=1'b0;
    defparam \pll_main.zim_pll_inst .DIVR=4'b0000;
    defparam \pll_main.zim_pll_inst .DIVQ=3'b101;
    defparam \pll_main.zim_pll_inst .DIVF=7'b0011111;
    defparam \pll_main.zim_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE \pll_main.zim_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(),
            .REFERENCECLK(N__19018),
            .RESETB(N__52877),
            .BYPASS(GNDG0),
            .PLLOUTCOREA(),
            .SDI(GNDG0),
            .PLLOUTGLOBALB(clk_16MHz),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(GNDG0),
            .PLLOUTGLOBALA(clk_32MHz),
            .SCLK(GNDG0));
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged2_physical (
            .RDATA({dangling_wire_0,dangling_wire_1,buf_data_iac_19,dangling_wire_2,dangling_wire_3,dangling_wire_4,buf_data_vac_19,dangling_wire_5,dangling_wire_6,dangling_wire_7,buf_data_iac_18,dangling_wire_8,dangling_wire_9,dangling_wire_10,buf_data_vac_18,dangling_wire_11}),
            .RADDR({dangling_wire_12,N__42985,N__24526,N__20374,N__43942,N__42238,N__39010,N__31453,N__36502,N__43183,N__31612}),
            .WADDR({dangling_wire_13,N__40471,N__40579,N__39409,N__39514,N__39622,N__39730,N__39832,N__39940,N__40045,N__40150}),
            .MASK({dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29}),
            .WDATA({dangling_wire_30,dangling_wire_31,N__26077,dangling_wire_32,dangling_wire_33,dangling_wire_34,N__21073,dangling_wire_35,dangling_wire_36,dangling_wire_37,N__27811,dangling_wire_38,dangling_wire_39,dangling_wire_40,N__23856,dangling_wire_41}),
            .RCLKE(),
            .RCLK(N__55158),
            .RE(N__52860),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged2WCLKN_net),
            .WE(N__31753));
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged7_physical (
            .RDATA({dangling_wire_42,dangling_wire_43,buf_data_iac_9,dangling_wire_44,dangling_wire_45,dangling_wire_46,buf_data_vac_9,dangling_wire_47,dangling_wire_48,dangling_wire_49,buf_data_iac_8,dangling_wire_50,dangling_wire_51,dangling_wire_52,buf_data_vac_8,dangling_wire_53}),
            .RADDR({dangling_wire_54,N__42945,N__24480,N__20322,N__43902,N__42201,N__38970,N__31413,N__36468,N__43149,N__31578}),
            .WADDR({dangling_wire_55,N__40437,N__40548,N__39369,N__39477,N__39588,N__39696,N__39792,N__39906,N__40011,N__40116}),
            .MASK({dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71}),
            .WDATA({dangling_wire_72,dangling_wire_73,N__21676,dangling_wire_74,dangling_wire_75,dangling_wire_76,N__35284,dangling_wire_77,dangling_wire_78,dangling_wire_79,N__24424,dangling_wire_80,dangling_wire_81,dangling_wire_82,N__21397,dangling_wire_83}),
            .RCLKE(),
            .RCLK(N__55245),
            .RE(N__52888),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged7WCLKN_net),
            .WE(N__31751));
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged1_physical (
            .RDATA({dangling_wire_84,dangling_wire_85,buf_data_iac_21,dangling_wire_86,dangling_wire_87,dangling_wire_88,buf_data_vac_21,dangling_wire_89,dangling_wire_90,dangling_wire_91,buf_data_iac_20,dangling_wire_92,dangling_wire_93,dangling_wire_94,buf_data_vac_20,dangling_wire_95}),
            .RADDR({dangling_wire_96,N__43003,N__24544,N__20392,N__43960,N__42256,N__39028,N__31471,N__36520,N__43201,N__31630}),
            .WADDR({dangling_wire_97,N__40489,N__40597,N__39427,N__39532,N__39640,N__39748,N__39850,N__39958,N__40063,N__40168}),
            .MASK({dangling_wire_98,dangling_wire_99,dangling_wire_100,dangling_wire_101,dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,dangling_wire_109,dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113}),
            .WDATA({dangling_wire_114,dangling_wire_115,N__27301,dangling_wire_116,dangling_wire_117,dangling_wire_118,N__21856,dangling_wire_119,dangling_wire_120,dangling_wire_121,N__28138,dangling_wire_122,dangling_wire_123,dangling_wire_124,N__25711,dangling_wire_125}),
            .RCLKE(),
            .RCLK(N__55093),
            .RE(N__52873),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged1WCLKN_net),
            .WE(N__31776));
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged6_physical (
            .RDATA({dangling_wire_126,dangling_wire_127,buf_data_iac_11,dangling_wire_128,dangling_wire_129,dangling_wire_130,buf_data_vac_11,dangling_wire_131,dangling_wire_132,dangling_wire_133,buf_data_iac_10,dangling_wire_134,dangling_wire_135,dangling_wire_136,buf_data_vac_10,dangling_wire_137}),
            .RADDR({dangling_wire_138,N__42957,N__24492,N__20334,N__43914,N__42213,N__38982,N__31425,N__36478,N__43159,N__31588}),
            .WADDR({dangling_wire_139,N__40447,N__40555,N__39381,N__39489,N__39598,N__39706,N__39804,N__39916,N__40021,N__40126}),
            .MASK({dangling_wire_140,dangling_wire_141,dangling_wire_142,dangling_wire_143,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,dangling_wire_151,dangling_wire_152,dangling_wire_153,dangling_wire_154,dangling_wire_155}),
            .WDATA({dangling_wire_156,dangling_wire_157,N__33533,dangling_wire_158,dangling_wire_159,dangling_wire_160,N__25897,dangling_wire_161,dangling_wire_162,dangling_wire_163,N__25969,dangling_wire_164,dangling_wire_165,dangling_wire_166,N__24055,dangling_wire_167}),
            .RCLKE(),
            .RCLK(N__55242),
            .RE(N__52887),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged6WCLKN_net),
            .WE(N__31719));
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged0_physical (
            .RDATA({dangling_wire_168,dangling_wire_169,buf_data_iac_23,dangling_wire_170,dangling_wire_171,dangling_wire_172,buf_data_vac_23,dangling_wire_173,dangling_wire_174,dangling_wire_175,buf_data_iac_22,dangling_wire_176,dangling_wire_177,dangling_wire_178,buf_data_vac_22,dangling_wire_179}),
            .RADDR({dangling_wire_180,N__43009,N__24550,N__20398,N__43966,N__42262,N__39034,N__31477,N__36526,N__43207,N__31636}),
            .WADDR({dangling_wire_181,N__40495,N__40603,N__39433,N__39538,N__39646,N__39754,N__39856,N__39964,N__40069,N__40174}),
            .MASK({dangling_wire_182,dangling_wire_183,dangling_wire_184,dangling_wire_185,dangling_wire_186,dangling_wire_187,dangling_wire_188,dangling_wire_189,dangling_wire_190,dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197}),
            .WDATA({dangling_wire_198,dangling_wire_199,N__26275,dangling_wire_200,dangling_wire_201,dangling_wire_202,N__24346,dangling_wire_203,dangling_wire_204,dangling_wire_205,N__24700,dangling_wire_206,dangling_wire_207,dangling_wire_208,N__22711,dangling_wire_209}),
            .RCLKE(),
            .RCLK(N__55079),
            .RE(N__52886),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged0WCLKN_net),
            .WE(N__31777));
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged5_physical (
            .RDATA({dangling_wire_210,dangling_wire_211,buf_data_iac_13,dangling_wire_212,dangling_wire_213,dangling_wire_214,buf_data_vac_13,dangling_wire_215,dangling_wire_216,dangling_wire_217,buf_data_iac_12,dangling_wire_218,dangling_wire_219,dangling_wire_220,buf_data_vac_12,dangling_wire_221}),
            .RADDR({dangling_wire_222,N__42967,N__24504,N__20346,N__43924,N__42220,N__38992,N__31435,N__36484,N__43165,N__31594}),
            .WADDR({dangling_wire_223,N__40453,N__40561,N__39391,N__39496,N__39604,N__39712,N__39814,N__39922,N__40027,N__40132}),
            .MASK({dangling_wire_224,dangling_wire_225,dangling_wire_226,dangling_wire_227,dangling_wire_228,dangling_wire_229,dangling_wire_230,dangling_wire_231,dangling_wire_232,dangling_wire_233,dangling_wire_234,dangling_wire_235,dangling_wire_236,dangling_wire_237,dangling_wire_238,dangling_wire_239}),
            .WDATA({dangling_wire_240,dangling_wire_241,N__25812,dangling_wire_242,dangling_wire_243,dangling_wire_244,N__21540,dangling_wire_245,dangling_wire_246,dangling_wire_247,N__33461,dangling_wire_248,dangling_wire_249,dangling_wire_250,N__24097,dangling_wire_251}),
            .RCLKE(),
            .RCLK(N__55235),
            .RE(N__52879),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged5WCLKN_net),
            .WE(N__31750));
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged9_physical (
            .RDATA({dangling_wire_252,dangling_wire_253,buf_data_iac_5,dangling_wire_254,dangling_wire_255,dangling_wire_256,buf_data_vac_5,dangling_wire_257,dangling_wire_258,dangling_wire_259,buf_data_iac_4,dangling_wire_260,dangling_wire_261,dangling_wire_262,buf_data_vac_4,dangling_wire_263}),
            .RADDR({dangling_wire_264,N__42954,N__24501,N__20355,N__43911,N__42204,N__38979,N__31422,N__36465,N__43146,N__31575}),
            .WADDR({dangling_wire_265,N__40434,N__40539,N__39378,N__39480,N__39585,N__39693,N__39801,N__39903,N__40008,N__40113}),
            .MASK({dangling_wire_266,dangling_wire_267,dangling_wire_268,dangling_wire_269,dangling_wire_270,dangling_wire_271,dangling_wire_272,dangling_wire_273,dangling_wire_274,dangling_wire_275,dangling_wire_276,dangling_wire_277,dangling_wire_278,dangling_wire_279,dangling_wire_280,dangling_wire_281}),
            .WDATA({dangling_wire_282,dangling_wire_283,N__49078,dangling_wire_284,dangling_wire_285,dangling_wire_286,N__38308,dangling_wire_287,dangling_wire_288,dangling_wire_289,N__48829,dangling_wire_290,dangling_wire_291,dangling_wire_292,N__51331,dangling_wire_293}),
            .RCLKE(),
            .RCLK(N__55225),
            .RE(N__52836),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged9WCLKN_net),
            .WE(N__31766));
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged4_physical (
            .RDATA({dangling_wire_294,dangling_wire_295,buf_data_iac_15,dangling_wire_296,dangling_wire_297,dangling_wire_298,buf_data_vac_15,dangling_wire_299,dangling_wire_300,dangling_wire_301,buf_data_iac_14,dangling_wire_302,dangling_wire_303,dangling_wire_304,buf_data_vac_14,dangling_wire_305}),
            .RADDR({dangling_wire_306,N__42973,N__24514,N__20358,N__43930,N__42226,N__38998,N__31441,N__36490,N__43171,N__31600}),
            .WADDR({dangling_wire_307,N__40459,N__40567,N__39397,N__39502,N__39610,N__39718,N__39820,N__39928,N__40033,N__40138}),
            .MASK({dangling_wire_308,dangling_wire_309,dangling_wire_310,dangling_wire_311,dangling_wire_312,dangling_wire_313,dangling_wire_314,dangling_wire_315,dangling_wire_316,dangling_wire_317,dangling_wire_318,dangling_wire_319,dangling_wire_320,dangling_wire_321,dangling_wire_322,dangling_wire_323}),
            .WDATA({dangling_wire_324,dangling_wire_325,N__31990,dangling_wire_326,dangling_wire_327,dangling_wire_328,N__20197,dangling_wire_329,dangling_wire_330,dangling_wire_331,N__29586,dangling_wire_332,dangling_wire_333,dangling_wire_334,N__22681,dangling_wire_335}),
            .RCLKE(),
            .RCLK(N__55214),
            .RE(N__52878),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged4WCLKN_net),
            .WE(N__31726));
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged8_physical (
            .RDATA({dangling_wire_336,dangling_wire_337,buf_data_iac_7,dangling_wire_338,dangling_wire_339,dangling_wire_340,buf_data_vac_7,dangling_wire_341,dangling_wire_342,dangling_wire_343,buf_data_iac_6,dangling_wire_344,dangling_wire_345,dangling_wire_346,buf_data_vac_6,dangling_wire_347}),
            .RADDR({dangling_wire_348,N__42966,N__24513,N__20367,N__43923,N__42216,N__38991,N__31434,N__36477,N__43158,N__31587}),
            .WADDR({dangling_wire_349,N__40446,N__40551,N__39390,N__39492,N__39597,N__39705,N__39813,N__39915,N__40020,N__40125}),
            .MASK({dangling_wire_350,dangling_wire_351,dangling_wire_352,dangling_wire_353,dangling_wire_354,dangling_wire_355,dangling_wire_356,dangling_wire_357,dangling_wire_358,dangling_wire_359,dangling_wire_360,dangling_wire_361,dangling_wire_362,dangling_wire_363,dangling_wire_364,dangling_wire_365}),
            .WDATA({dangling_wire_366,dangling_wire_367,N__47881,dangling_wire_368,dangling_wire_369,dangling_wire_370,N__47932,dangling_wire_371,dangling_wire_372,dangling_wire_373,N__48565,dangling_wire_374,dangling_wire_375,dangling_wire_376,N__40864,dangling_wire_377}),
            .RCLKE(),
            .RCLK(N__55202),
            .RE(N__52835),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged8WCLKN_net),
            .WE(N__31767));
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged10_physical (
            .RDATA({dangling_wire_378,dangling_wire_379,buf_data_iac_3,dangling_wire_380,dangling_wire_381,dangling_wire_382,buf_data_vac_3,dangling_wire_383,dangling_wire_384,dangling_wire_385,buf_data_iac_2,dangling_wire_386,dangling_wire_387,dangling_wire_388,buf_data_vac_2,dangling_wire_389}),
            .RADDR({dangling_wire_390,N__42997,N__24538,N__20386,N__43954,N__42250,N__39022,N__31465,N__36514,N__43195,N__31624}),
            .WADDR({dangling_wire_391,N__40483,N__40591,N__39421,N__39526,N__39634,N__39742,N__39844,N__39952,N__40057,N__40162}),
            .MASK({dangling_wire_392,dangling_wire_393,dangling_wire_394,dangling_wire_395,dangling_wire_396,dangling_wire_397,dangling_wire_398,dangling_wire_399,dangling_wire_400,dangling_wire_401,dangling_wire_402,dangling_wire_403,dangling_wire_404,dangling_wire_405,dangling_wire_406,dangling_wire_407}),
            .WDATA({dangling_wire_408,dangling_wire_409,N__21046,dangling_wire_410,dangling_wire_411,dangling_wire_412,N__21481,dangling_wire_413,dangling_wire_414,dangling_wire_415,N__22495,dangling_wire_416,dangling_wire_417,dangling_wire_418,N__22435,dangling_wire_419}),
            .RCLKE(),
            .RCLK(N__55110),
            .RE(N__52837),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged10WCLKN_net),
            .WE(N__31769));
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged3_physical (
            .RDATA({dangling_wire_420,dangling_wire_421,buf_data_iac_17,dangling_wire_422,dangling_wire_423,dangling_wire_424,buf_data_vac_17,dangling_wire_425,dangling_wire_426,dangling_wire_427,buf_data_iac_16,dangling_wire_428,dangling_wire_429,dangling_wire_430,buf_data_vac_16,dangling_wire_431}),
            .RADDR({dangling_wire_432,N__42979,N__24520,N__20368,N__43936,N__42232,N__39004,N__31447,N__36496,N__43177,N__31606}),
            .WADDR({dangling_wire_433,N__40465,N__40573,N__39403,N__39508,N__39616,N__39724,N__39826,N__39934,N__40039,N__40144}),
            .MASK({dangling_wire_434,dangling_wire_435,dangling_wire_436,dangling_wire_437,dangling_wire_438,dangling_wire_439,dangling_wire_440,dangling_wire_441,dangling_wire_442,dangling_wire_443,dangling_wire_444,dangling_wire_445,dangling_wire_446,dangling_wire_447,dangling_wire_448,dangling_wire_449}),
            .WDATA({dangling_wire_450,dangling_wire_451,N__26038,dangling_wire_452,dangling_wire_453,dangling_wire_454,N__22657,dangling_wire_455,dangling_wire_456,dangling_wire_457,N__27997,dangling_wire_458,dangling_wire_459,dangling_wire_460,N__22595,dangling_wire_461}),
            .RCLKE(),
            .RCLK(N__55188),
            .RE(N__52861),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged3WCLKN_net),
            .WE(N__31752));
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged11_physical (
            .RDATA({dangling_wire_462,dangling_wire_463,buf_data_iac_1,dangling_wire_464,dangling_wire_465,dangling_wire_466,buf_data_vac_1,dangling_wire_467,dangling_wire_468,dangling_wire_469,buf_data_iac_0,dangling_wire_470,dangling_wire_471,dangling_wire_472,buf_data_vac_0,dangling_wire_473}),
            .RADDR({dangling_wire_474,N__42991,N__24532,N__20380,N__43948,N__42244,N__39016,N__31459,N__36508,N__43189,N__31618}),
            .WADDR({dangling_wire_475,N__40477,N__40585,N__39415,N__39520,N__39628,N__39736,N__39838,N__39946,N__40051,N__40156}),
            .MASK({dangling_wire_476,dangling_wire_477,dangling_wire_478,dangling_wire_479,dangling_wire_480,dangling_wire_481,dangling_wire_482,dangling_wire_483,dangling_wire_484,dangling_wire_485,dangling_wire_486,dangling_wire_487,dangling_wire_488,dangling_wire_489,dangling_wire_490,dangling_wire_491}),
            .WDATA({dangling_wire_492,dangling_wire_493,N__23628,dangling_wire_494,dangling_wire_495,dangling_wire_496,N__23968,dangling_wire_497,dangling_wire_498,dangling_wire_499,N__23458,dangling_wire_500,dangling_wire_501,dangling_wire_502,N__23482,dangling_wire_503}),
            .RCLKE(),
            .RCLK(N__55131),
            .RE(N__52723),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged11WCLKN_net),
            .WE(N__31768));
    IO_PAD ipInertedIOPad_VAC_DRDY_iopad (
            .OE(N__58652),
            .DIN(N__58651),
            .DOUT(N__58650),
            .PACKAGEPIN(VAC_DRDY));
    defparam ipInertedIOPad_VAC_DRDY_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VAC_DRDY_preio (
            .PADOEN(N__58652),
            .PADOUT(N__58651),
            .PADIN(N__58650),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(VAC_DRDY),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_FLT1_iopad (
            .OE(N__58643),
            .DIN(N__58642),
            .DOUT(N__58641),
            .PACKAGEPIN(IAC_FLT1));
    defparam ipInertedIOPad_IAC_FLT1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_FLT1_preio (
            .PADOEN(N__58643),
            .PADOUT(N__58642),
            .PADIN(N__58641),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__28099),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_SCK_iopad (
            .OE(N__58634),
            .DIN(N__58633),
            .DOUT(N__58632),
            .PACKAGEPIN(DDS_SCK));
    defparam ipInertedIOPad_DDS_SCK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_SCK_preio (
            .PADOEN(N__58634),
            .PADOUT(N__58633),
            .PADIN(N__58632),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__55915),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_166_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_166_iopad (
            .OE(N__58625),
            .DIN(N__58624),
            .DOUT(N__58623),
            .PACKAGEPIN(ICE_IOR_166));
    defparam ipInertedIOPad_ICE_IOR_166_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_166_preio (
            .PADOEN(N__58625),
            .PADOUT(N__58624),
            .PADIN(N__58623),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_119_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_119_iopad (
            .OE(N__58616),
            .DIN(N__58615),
            .DOUT(N__58614),
            .PACKAGEPIN(ICE_IOR_119));
    defparam ipInertedIOPad_ICE_IOR_119_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_119_preio (
            .PADOEN(N__58616),
            .PADOUT(N__58615),
            .PADIN(N__58614),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_MOSI_iopad (
            .OE(N__58607),
            .DIN(N__58606),
            .DOUT(N__58605),
            .PACKAGEPIN(DDS_MOSI));
    defparam ipInertedIOPad_DDS_MOSI_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_MOSI_preio (
            .PADOEN(N__58607),
            .PADOUT(N__58606),
            .PADIN(N__58605),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__42901),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_MISO_iopad (
            .OE(N__58598),
            .DIN(N__58597),
            .DOUT(N__58596),
            .PACKAGEPIN(VAC_MISO));
    defparam ipInertedIOPad_VAC_MISO_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VAC_MISO_preio (
            .PADOEN(N__58598),
            .PADOUT(N__58597),
            .PADIN(N__58596),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(VAC_MISO),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_MOSI1_iopad (
            .OE(N__58589),
            .DIN(N__58588),
            .DOUT(N__58587),
            .PACKAGEPIN(DDS_MOSI1));
    defparam ipInertedIOPad_DDS_MOSI1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_MOSI1_preio (
            .PADOEN(N__58589),
            .PADOUT(N__58588),
            .PADIN(N__58587),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__21874),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_146_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_146_iopad (
            .OE(N__58580),
            .DIN(N__58579),
            .DOUT(N__58578),
            .PACKAGEPIN(ICE_IOR_146));
    defparam ipInertedIOPad_ICE_IOR_146_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_146_preio (
            .PADOEN(N__58580),
            .PADOUT(N__58579),
            .PADIN(N__58578),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VDC_CLK_iopad (
            .OE(N__58571),
            .DIN(N__58570),
            .DOUT(N__58569),
            .PACKAGEPIN(VDC_CLK));
    defparam ipInertedIOPad_VDC_CLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VDC_CLK_preio (
            .PADOEN(N__58571),
            .PADOUT(N__58570),
            .PADIN(N__58569),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__32914),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_222_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_222_iopad (
            .OE(N__58562),
            .DIN(N__58561),
            .DOUT(N__58560),
            .PACKAGEPIN(ICE_IOT_222));
    defparam ipInertedIOPad_ICE_IOT_222_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_222_preio (
            .PADOEN(N__58562),
            .PADOUT(N__58561),
            .PADIN(N__58560),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_CS_iopad (
            .OE(N__58553),
            .DIN(N__58552),
            .DOUT(N__58551),
            .PACKAGEPIN(IAC_CS));
    defparam ipInertedIOPad_IAC_CS_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_CS_preio (
            .PADOEN(N__58553),
            .PADOUT(N__58552),
            .PADIN(N__58551),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__24847),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_18B_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_18B_iopad (
            .OE(N__58544),
            .DIN(N__58543),
            .DOUT(N__58542),
            .PACKAGEPIN(ICE_IOL_18B));
    defparam ipInertedIOPad_ICE_IOL_18B_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_18B_preio (
            .PADOEN(N__58544),
            .PADOUT(N__58543),
            .PADIN(N__58542),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_13A_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_13A_iopad (
            .OE(N__58535),
            .DIN(N__58534),
            .DOUT(N__58533),
            .PACKAGEPIN(ICE_IOL_13A));
    defparam ipInertedIOPad_ICE_IOL_13A_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_13A_preio (
            .PADOEN(N__58535),
            .PADOUT(N__58534),
            .PADIN(N__58533),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_ICE_IOB_81_iopad (
            .OE(N__58526),
            .DIN(N__58525),
            .DOUT(N__58524),
            .PACKAGEPIN(ICE_IOB_81));
    defparam ipInertedIOPad_ICE_IOB_81_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_81_preio (
            .PADOEN(N__58526),
            .PADOUT(N__58525),
            .PADIN(N__58524),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_OSR1_iopad (
            .OE(N__58517),
            .DIN(N__58516),
            .DOUT(N__58515),
            .PACKAGEPIN(VAC_OSR1));
    defparam ipInertedIOPad_VAC_OSR1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_OSR1_preio (
            .PADOEN(N__58517),
            .PADOUT(N__58516),
            .PADIN(N__58515),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__29725),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_MOSI_iopad (
            .OE(N__58508),
            .DIN(N__58507),
            .DOUT(N__58506),
            .PACKAGEPIN(IAC_MOSI));
    defparam ipInertedIOPad_IAC_MOSI_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_MOSI_preio (
            .PADOEN(N__58508),
            .PADOUT(N__58507),
            .PADIN(N__58506),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_CS1_iopad (
            .OE(N__58499),
            .DIN(N__58498),
            .DOUT(N__58497),
            .PACKAGEPIN(DDS_CS1));
    defparam ipInertedIOPad_DDS_CS1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_CS1_preio (
            .PADOEN(N__58499),
            .PADOUT(N__58498),
            .PADIN(N__58497),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__21631),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_4B_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_4B_iopad (
            .OE(N__58490),
            .DIN(N__58489),
            .DOUT(N__58488),
            .PACKAGEPIN(ICE_IOL_4B));
    defparam ipInertedIOPad_ICE_IOL_4B_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_4B_preio (
            .PADOEN(N__58490),
            .PADOUT(N__58489),
            .PADIN(N__58488),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOB_94_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOB_94_iopad (
            .OE(N__58481),
            .DIN(N__58480),
            .DOUT(N__58479),
            .PACKAGEPIN(ICE_IOB_94));
    defparam ipInertedIOPad_ICE_IOB_94_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_94_preio (
            .PADOEN(N__58481),
            .PADOUT(N__58480),
            .PADIN(N__58479),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_CS_iopad (
            .OE(N__58472),
            .DIN(N__58471),
            .DOUT(N__58470),
            .PACKAGEPIN(VAC_CS));
    defparam ipInertedIOPad_VAC_CS_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_CS_preio (
            .PADOEN(N__58472),
            .PADOUT(N__58471),
            .PADIN(N__58470),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__20254),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_CLK_iopad (
            .OE(N__58463),
            .DIN(N__58462),
            .DOUT(N__58461),
            .PACKAGEPIN(VAC_CLK));
    defparam ipInertedIOPad_VAC_CLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_CLK_preio (
            .PADOEN(N__58463),
            .PADOUT(N__58462),
            .PADIN(N__58461),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__26148),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_SPI_CE0_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_SPI_CE0_iopad (
            .OE(N__58454),
            .DIN(N__58453),
            .DOUT(N__58452),
            .PACKAGEPIN(ICE_SPI_CE0));
    defparam ipInertedIOPad_ICE_SPI_CE0_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_SPI_CE0_preio (
            .PADOEN(N__58454),
            .PADOUT(N__58453),
            .PADIN(N__58452),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(ICE_SPI_CE0),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_167_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_167_iopad (
            .OE(N__58445),
            .DIN(N__58444),
            .DOUT(N__58443),
            .PACKAGEPIN(ICE_IOR_167));
    defparam ipInertedIOPad_ICE_IOR_167_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_167_preio (
            .PADOEN(N__58445),
            .PADOUT(N__58444),
            .PADIN(N__58443),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_118_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_118_iopad (
            .OE(N__58436),
            .DIN(N__58435),
            .DOUT(N__58434),
            .PACKAGEPIN(ICE_IOR_118));
    defparam ipInertedIOPad_ICE_IOR_118_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_118_preio (
            .PADOEN(N__58436),
            .PADOUT(N__58435),
            .PADIN(N__58434),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_RTD_SDO_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_RTD_SDO_iopad (
            .OE(N__58427),
            .DIN(N__58426),
            .DOUT(N__58425),
            .PACKAGEPIN(RTD_SDO));
    defparam ipInertedIOPad_RTD_SDO_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_RTD_SDO_preio (
            .PADOEN(N__58427),
            .PADOUT(N__58426),
            .PADIN(N__58425),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(RTD_SDO),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_OSR0_iopad (
            .OE(N__58418),
            .DIN(N__58417),
            .DOUT(N__58416),
            .PACKAGEPIN(IAC_OSR0));
    defparam ipInertedIOPad_IAC_OSR0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_OSR0_preio (
            .PADOEN(N__58418),
            .PADOUT(N__58417),
            .PADIN(N__58416),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__28225),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VDC_SCLK_iopad (
            .OE(N__58409),
            .DIN(N__58408),
            .DOUT(N__58407),
            .PACKAGEPIN(VDC_SCLK));
    defparam ipInertedIOPad_VDC_SCLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VDC_SCLK_preio (
            .PADOEN(N__58409),
            .PADOUT(N__58408),
            .PADIN(N__58407),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__26938),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_FLT1_iopad (
            .OE(N__58400),
            .DIN(N__58399),
            .DOUT(N__58398),
            .PACKAGEPIN(VAC_FLT1));
    defparam ipInertedIOPad_VAC_FLT1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_FLT1_preio (
            .PADOEN(N__58400),
            .PADOUT(N__58399),
            .PADIN(N__58398),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__26221),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_SPI_MOSI_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_SPI_MOSI_iopad (
            .OE(N__58391),
            .DIN(N__58390),
            .DOUT(N__58389),
            .PACKAGEPIN(ICE_SPI_MOSI));
    defparam ipInertedIOPad_ICE_SPI_MOSI_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_SPI_MOSI_preio (
            .PADOEN(N__58391),
            .PADOUT(N__58390),
            .PADIN(N__58389),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(ICE_SPI_MOSI),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_165_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_165_iopad (
            .OE(N__58382),
            .DIN(N__58381),
            .DOUT(N__58380),
            .PACKAGEPIN(ICE_IOR_165));
    defparam ipInertedIOPad_ICE_IOR_165_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_165_preio (
            .PADOEN(N__58382),
            .PADOUT(N__58381),
            .PADIN(N__58380),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_147_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_147_iopad (
            .OE(N__58373),
            .DIN(N__58372),
            .DOUT(N__58371),
            .PACKAGEPIN(ICE_IOR_147));
    defparam ipInertedIOPad_ICE_IOR_147_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_147_preio (
            .PADOEN(N__58373),
            .PADOUT(N__58372),
            .PADIN(N__58371),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_14A_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_14A_iopad (
            .OE(N__58364),
            .DIN(N__58363),
            .DOUT(N__58362),
            .PACKAGEPIN(ICE_IOL_14A));
    defparam ipInertedIOPad_ICE_IOL_14A_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_14A_preio (
            .PADOEN(N__58364),
            .PADOUT(N__58363),
            .PADIN(N__58362),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_13B_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_13B_iopad (
            .OE(N__58355),
            .DIN(N__58354),
            .DOUT(N__58353),
            .PACKAGEPIN(ICE_IOL_13B));
    defparam ipInertedIOPad_ICE_IOL_13B_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_13B_preio (
            .PADOEN(N__58355),
            .PADOUT(N__58354),
            .PADIN(N__58353),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOB_91_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOB_91_iopad (
            .OE(N__58346),
            .DIN(N__58345),
            .DOUT(N__58344),
            .PACKAGEPIN(ICE_IOB_91));
    defparam ipInertedIOPad_ICE_IOB_91_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_91_preio (
            .PADOEN(N__58346),
            .PADOUT(N__58345),
            .PADIN(N__58344),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_GPMO_0_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_GPMO_0_iopad (
            .OE(N__58337),
            .DIN(N__58336),
            .DOUT(N__58335),
            .PACKAGEPIN(ICE_GPMO_0));
    defparam ipInertedIOPad_ICE_GPMO_0_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_GPMO_0_preio (
            .PADOEN(N__58337),
            .PADOUT(N__58336),
            .PADIN(N__58335),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_RNG_0_iopad (
            .OE(N__58328),
            .DIN(N__58327),
            .DOUT(N__58326),
            .PACKAGEPIN(DDS_RNG_0));
    defparam ipInertedIOPad_DDS_RNG_0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_RNG_0_preio (
            .PADOEN(N__58328),
            .PADOUT(N__58327),
            .PADIN(N__58326),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__44035),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VDC_RNG0_iopad (
            .OE(N__58319),
            .DIN(N__58318),
            .DOUT(N__58317),
            .PACKAGEPIN(VDC_RNG0));
    defparam ipInertedIOPad_VDC_RNG0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VDC_RNG0_preio (
            .PADOEN(N__58319),
            .PADOUT(N__58318),
            .PADIN(N__58317),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__44767),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_SPI_SCLK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_SPI_SCLK_iopad (
            .OE(N__58310),
            .DIN(N__58309),
            .DOUT(N__58308),
            .PACKAGEPIN(ICE_SPI_SCLK));
    defparam ipInertedIOPad_ICE_SPI_SCLK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_SPI_SCLK_preio (
            .PADOEN(N__58310),
            .PADOUT(N__58309),
            .PADIN(N__58308),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(ICE_SPI_SCLK),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_152_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_152_iopad (
            .OE(N__58301),
            .DIN(N__58300),
            .DOUT(N__58299),
            .PACKAGEPIN(ICE_IOR_152));
    defparam ipInertedIOPad_ICE_IOR_152_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_152_preio (
            .PADOEN(N__58301),
            .PADOUT(N__58300),
            .PADIN(N__58299),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_12A_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_12A_iopad (
            .OE(N__58292),
            .DIN(N__58291),
            .DOUT(N__58290),
            .PACKAGEPIN(ICE_IOL_12A));
    defparam ipInertedIOPad_ICE_IOL_12A_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_12A_preio (
            .PADOEN(N__58292),
            .PADOUT(N__58291),
            .PADIN(N__58290),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_RTD_DRDY_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_RTD_DRDY_iopad (
            .OE(N__58283),
            .DIN(N__58282),
            .DOUT(N__58281),
            .PACKAGEPIN(RTD_DRDY));
    defparam ipInertedIOPad_RTD_DRDY_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_RTD_DRDY_preio (
            .PADOEN(N__58283),
            .PADOUT(N__58282),
            .PADIN(N__58281),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(RTD_DRDY),
            .DIN1());
    IO_PAD ipInertedIOPad_ICE_SPI_MISO_iopad (
            .OE(N__58274),
            .DIN(N__58273),
            .DOUT(N__58272),
            .PACKAGEPIN(ICE_SPI_MISO));
    defparam ipInertedIOPad_ICE_SPI_MISO_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_ICE_SPI_MISO_preio (
            .PADOEN(N__58274),
            .PADOUT(N__58273),
            .PADIN(N__58272),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__43591),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_177_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_177_iopad (
            .OE(N__58265),
            .DIN(N__58264),
            .DOUT(N__58263),
            .PACKAGEPIN(ICE_IOT_177));
    defparam ipInertedIOPad_ICE_IOT_177_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_177_preio (
            .PADOEN(N__58265),
            .PADOUT(N__58264),
            .PADIN(N__58263),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_141_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_141_iopad (
            .OE(N__58256),
            .DIN(N__58255),
            .DOUT(N__58254),
            .PACKAGEPIN(ICE_IOR_141));
    defparam ipInertedIOPad_ICE_IOR_141_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_141_preio (
            .PADOEN(N__58256),
            .PADOUT(N__58255),
            .PADIN(N__58254),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOB_80_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOB_80_iopad (
            .OE(N__58247),
            .DIN(N__58246),
            .DOUT(N__58245),
            .PACKAGEPIN(ICE_IOB_80));
    defparam ipInertedIOPad_ICE_IOB_80_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_80_preio (
            .PADOEN(N__58247),
            .PADOUT(N__58246),
            .PADIN(N__58245),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOB_102_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOB_102_iopad (
            .OE(N__58238),
            .DIN(N__58237),
            .DOUT(N__58236),
            .PACKAGEPIN(ICE_IOB_102));
    defparam ipInertedIOPad_ICE_IOB_102_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_102_preio (
            .PADOEN(N__58238),
            .PADOUT(N__58237),
            .PADIN(N__58236),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_GPMO_2_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_GPMO_2_iopad (
            .OE(N__58229),
            .DIN(N__58228),
            .DOUT(N__58227),
            .PACKAGEPIN(ICE_GPMO_2));
    defparam ipInertedIOPad_ICE_GPMO_2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_GPMO_2_preio (
            .PADOEN(N__58229),
            .PADOUT(N__58228),
            .PADIN(N__58227),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(ICE_GPMO_2),
            .DIN1());
    IO_PAD ipInertedIOPad_ICE_GPMI_0_iopad (
            .OE(N__58220),
            .DIN(N__58219),
            .DOUT(N__58218),
            .PACKAGEPIN(ICE_GPMI_0));
    defparam ipInertedIOPad_ICE_GPMI_0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_ICE_GPMI_0_preio (
            .PADOEN(N__58220),
            .PADOUT(N__58219),
            .PADIN(N__58218),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__49267),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_MISO_iopad (
            .OE(N__58211),
            .DIN(N__58210),
            .DOUT(N__58209),
            .PACKAGEPIN(IAC_MISO));
    defparam ipInertedIOPad_IAC_MISO_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_IAC_MISO_preio (
            .PADOEN(N__58211),
            .PADOUT(N__58210),
            .PADIN(N__58209),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(IAC_MISO),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_OSR0_iopad (
            .OE(N__58202),
            .DIN(N__58201),
            .DOUT(N__58200),
            .PACKAGEPIN(VAC_OSR0));
    defparam ipInertedIOPad_VAC_OSR0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_OSR0_preio (
            .PADOEN(N__58202),
            .PADOUT(N__58201),
            .PADIN(N__58200),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__26113),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_MOSI_iopad (
            .OE(N__58193),
            .DIN(N__58192),
            .DOUT(N__58191),
            .PACKAGEPIN(VAC_MOSI));
    defparam ipInertedIOPad_VAC_MOSI_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_MOSI_preio (
            .PADOEN(N__58193),
            .PADOUT(N__58192),
            .PADIN(N__58191),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_TEST_LED_iopad (
            .OE(N__58184),
            .DIN(N__58183),
            .DOUT(N__58182),
            .PACKAGEPIN(TEST_LED));
    defparam ipInertedIOPad_TEST_LED_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_TEST_LED_preio (
            .PADOEN(N__58184),
            .PADOUT(N__58183),
            .PADIN(N__58182),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__40945),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_148_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_148_iopad (
            .OE(N__58175),
            .DIN(N__58174),
            .DOUT(N__58173),
            .PACKAGEPIN(ICE_IOR_148));
    defparam ipInertedIOPad_ICE_IOR_148_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_148_preio (
            .PADOEN(N__58175),
            .PADOUT(N__58174),
            .PADIN(N__58173),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_STAT_COMM_iopad (
            .OE(N__58166),
            .DIN(N__58165),
            .DOUT(N__58164),
            .PACKAGEPIN(STAT_COMM));
    defparam ipInertedIOPad_STAT_COMM_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_STAT_COMM_preio (
            .PADOEN(N__58166),
            .PADOUT(N__58165),
            .PADIN(N__58164),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__19003),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_SYSCLK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_SYSCLK_iopad (
            .OE(N__58157),
            .DIN(N__58156),
            .DOUT(N__58155),
            .PACKAGEPIN(ICE_SYSCLK));
    defparam ipInertedIOPad_ICE_SYSCLK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_SYSCLK_preio (
            .PADOEN(N__58157),
            .PADOUT(N__58156),
            .PADIN(N__58155),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(ICE_SYSCLK),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_161_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_161_iopad (
            .OE(N__58148),
            .DIN(N__58147),
            .DOUT(N__58146),
            .PACKAGEPIN(ICE_IOR_161));
    defparam ipInertedIOPad_ICE_IOR_161_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_161_preio (
            .PADOEN(N__58148),
            .PADOUT(N__58147),
            .PADIN(N__58146),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOB_95_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOB_95_iopad (
            .OE(N__58139),
            .DIN(N__58138),
            .DOUT(N__58137),
            .PACKAGEPIN(ICE_IOB_95));
    defparam ipInertedIOPad_ICE_IOB_95_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_95_preio (
            .PADOEN(N__58139),
            .PADOUT(N__58138),
            .PADIN(N__58137),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_ICE_IOB_82_iopad (
            .OE(N__58130),
            .DIN(N__58129),
            .DOUT(N__58128),
            .PACKAGEPIN(ICE_IOB_82));
    defparam ipInertedIOPad_ICE_IOB_82_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_82_preio (
            .PADOEN(N__58130),
            .PADOUT(N__58129),
            .PADIN(N__58128),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_ICE_IOB_104_iopad (
            .OE(N__58121),
            .DIN(N__58120),
            .DOUT(N__58119),
            .PACKAGEPIN(ICE_IOB_104));
    defparam ipInertedIOPad_ICE_IOB_104_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_104_preio (
            .PADOEN(N__58121),
            .PADOUT(N__58120),
            .PADIN(N__58119),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_CLK_iopad (
            .OE(N__58112),
            .DIN(N__58111),
            .DOUT(N__58110),
            .PACKAGEPIN(IAC_CLK));
    defparam ipInertedIOPad_IAC_CLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_CLK_preio (
            .PADOEN(N__58112),
            .PADOUT(N__58111),
            .PADIN(N__58110),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__26152),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_CS_iopad (
            .OE(N__58103),
            .DIN(N__58102),
            .DOUT(N__58101),
            .PACKAGEPIN(DDS_CS));
    defparam ipInertedIOPad_DDS_CS_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_CS_preio (
            .PADOEN(N__58103),
            .PADOUT(N__58102),
            .PADIN(N__58101),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__55504),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SELIRNG0_iopad (
            .OE(N__58094),
            .DIN(N__58093),
            .DOUT(N__58092),
            .PACKAGEPIN(SELIRNG0));
    defparam ipInertedIOPad_SELIRNG0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_SELIRNG0_preio (
            .PADOEN(N__58094),
            .PADOUT(N__58093),
            .PADIN(N__58092),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__38185),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_RTD_SDI_iopad (
            .OE(N__58085),
            .DIN(N__58084),
            .DOUT(N__58083),
            .PACKAGEPIN(RTD_SDI));
    defparam ipInertedIOPad_RTD_SDI_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_RTD_SDI_preio (
            .PADOEN(N__58085),
            .PADOUT(N__58084),
            .PADIN(N__58083),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__19798),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_221_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_221_iopad (
            .OE(N__58076),
            .DIN(N__58075),
            .DOUT(N__58074),
            .PACKAGEPIN(ICE_IOT_221));
    defparam ipInertedIOPad_ICE_IOT_221_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_221_preio (
            .PADOEN(N__58076),
            .PADOUT(N__58075),
            .PADIN(N__58074),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_197_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_197_iopad (
            .OE(N__58067),
            .DIN(N__58066),
            .DOUT(N__58065),
            .PACKAGEPIN(ICE_IOT_197));
    defparam ipInertedIOPad_ICE_IOT_197_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_197_preio (
            .PADOEN(N__58067),
            .PADOUT(N__58066),
            .PADIN(N__58065),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_MCLK_iopad (
            .OE(N__58058),
            .DIN(N__58057),
            .DOUT(N__58056),
            .PACKAGEPIN(DDS_MCLK));
    defparam ipInertedIOPad_DDS_MCLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_MCLK_preio (
            .PADOEN(N__58058),
            .PADOUT(N__58057),
            .PADIN(N__58056),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__55933),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_RTD_SCLK_iopad (
            .OE(N__58049),
            .DIN(N__58048),
            .DOUT(N__58047),
            .PACKAGEPIN(RTD_SCLK));
    defparam ipInertedIOPad_RTD_SCLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_RTD_SCLK_preio (
            .PADOEN(N__58049),
            .PADOUT(N__58048),
            .PADIN(N__58047),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__19045),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_RTD_CS_iopad (
            .OE(N__58040),
            .DIN(N__58039),
            .DOUT(N__58038),
            .PACKAGEPIN(RTD_CS));
    defparam ipInertedIOPad_RTD_CS_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_RTD_CS_preio (
            .PADOEN(N__58040),
            .PADOUT(N__58039),
            .PADIN(N__58038),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__19099),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_137_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_137_iopad (
            .OE(N__58031),
            .DIN(N__58030),
            .DOUT(N__58029),
            .PACKAGEPIN(ICE_IOR_137));
    defparam ipInertedIOPad_ICE_IOR_137_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_137_preio (
            .PADOEN(N__58031),
            .PADOUT(N__58030),
            .PADIN(N__58029),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_OSR1_iopad (
            .OE(N__58022),
            .DIN(N__58021),
            .DOUT(N__58020),
            .PACKAGEPIN(IAC_OSR1));
    defparam ipInertedIOPad_IAC_OSR1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_OSR1_preio (
            .PADOEN(N__58022),
            .PADOUT(N__58021),
            .PADIN(N__58020),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__28060),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_FLT0_iopad (
            .OE(N__58013),
            .DIN(N__58012),
            .DOUT(N__58011),
            .PACKAGEPIN(VAC_FLT0));
    defparam ipInertedIOPad_VAC_FLT0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_FLT0_preio (
            .PADOEN(N__58013),
            .PADOUT(N__58012),
            .PADIN(N__58011),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__27880),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_144_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_144_iopad (
            .OE(N__58004),
            .DIN(N__58003),
            .DOUT(N__58002),
            .PACKAGEPIN(ICE_IOR_144));
    defparam ipInertedIOPad_ICE_IOR_144_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_144_preio (
            .PADOEN(N__58004),
            .PADOUT(N__58003),
            .PADIN(N__58002),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_128_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_128_iopad (
            .OE(N__57995),
            .DIN(N__57994),
            .DOUT(N__57993),
            .PACKAGEPIN(ICE_IOR_128));
    defparam ipInertedIOPad_ICE_IOR_128_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_128_preio (
            .PADOEN(N__57995),
            .PADOUT(N__57994),
            .PADIN(N__57993),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_GPMO_1_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_GPMO_1_iopad (
            .OE(N__57986),
            .DIN(N__57985),
            .DOUT(N__57984),
            .PACKAGEPIN(ICE_GPMO_1));
    defparam ipInertedIOPad_ICE_GPMO_1_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_GPMO_1_preio (
            .PADOEN(N__57986),
            .PADOUT(N__57985),
            .PADIN(N__57984),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_SCLK_iopad (
            .OE(N__57977),
            .DIN(N__57976),
            .DOUT(N__57975),
            .PACKAGEPIN(IAC_SCLK));
    defparam ipInertedIOPad_IAC_SCLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_SCLK_preio (
            .PADOEN(N__57977),
            .PADOUT(N__57976),
            .PADIN(N__57975),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__26194),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_EIS_SYNCCLK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_EIS_SYNCCLK_iopad (
            .OE(N__57968),
            .DIN(N__57967),
            .DOUT(N__57966),
            .PACKAGEPIN(EIS_SYNCCLK));
    defparam ipInertedIOPad_EIS_SYNCCLK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_EIS_SYNCCLK_preio (
            .PADOEN(N__57968),
            .PADOUT(N__57967),
            .PADIN(N__57966),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(EIS_SYNCCLK),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_139_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_139_iopad (
            .OE(N__57959),
            .DIN(N__57958),
            .DOUT(N__57957),
            .PACKAGEPIN(ICE_IOR_139));
    defparam ipInertedIOPad_ICE_IOR_139_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_139_preio (
            .PADOEN(N__57959),
            .PADOUT(N__57958),
            .PADIN(N__57957),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_4A_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_4A_iopad (
            .OE(N__57950),
            .DIN(N__57949),
            .DOUT(N__57948),
            .PACKAGEPIN(ICE_IOL_4A));
    defparam ipInertedIOPad_ICE_IOL_4A_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_4A_preio (
            .PADOEN(N__57950),
            .PADOUT(N__57949),
            .PADIN(N__57948),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_SCLK_iopad (
            .OE(N__57941),
            .DIN(N__57940),
            .DOUT(N__57939),
            .PACKAGEPIN(VAC_SCLK));
    defparam ipInertedIOPad_VAC_SCLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_SCLK_preio (
            .PADOEN(N__57941),
            .PADOUT(N__57940),
            .PADIN(N__57939),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__20227),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_THERMOSTAT_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_THERMOSTAT_iopad (
            .OE(N__57932),
            .DIN(N__57931),
            .DOUT(N__57930),
            .PACKAGEPIN(THERMOSTAT));
    defparam ipInertedIOPad_THERMOSTAT_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_THERMOSTAT_preio (
            .PADOEN(N__57932),
            .PADOUT(N__57931),
            .PADIN(N__57930),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(THERMOSTAT),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_164_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_164_iopad (
            .OE(N__57923),
            .DIN(N__57922),
            .DOUT(N__57921),
            .PACKAGEPIN(ICE_IOR_164));
    defparam ipInertedIOPad_ICE_IOR_164_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_164_preio (
            .PADOEN(N__57923),
            .PADOUT(N__57922),
            .PADIN(N__57921),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_ICE_IOB_103_iopad (
            .OE(N__57914),
            .DIN(N__57913),
            .DOUT(N__57912),
            .PACKAGEPIN(ICE_IOB_103));
    defparam ipInertedIOPad_ICE_IOB_103_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_103_preio (
            .PADOEN(N__57914),
            .PADOUT(N__57913),
            .PADIN(N__57912),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_AMPV_POW_iopad (
            .OE(N__57905),
            .DIN(N__57904),
            .DOUT(N__57903),
            .PACKAGEPIN(AMPV_POW));
    defparam ipInertedIOPad_AMPV_POW_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_AMPV_POW_preio (
            .PADOEN(N__57905),
            .PADOUT(N__57904),
            .PADIN(N__57903),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__30058),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VDC_SDO_iopad (
            .OE(N__57896),
            .DIN(N__57895),
            .DOUT(N__57894),
            .PACKAGEPIN(VDC_SDO));
    defparam ipInertedIOPad_VDC_SDO_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VDC_SDO_preio (
            .PADOEN(N__57896),
            .PADOUT(N__57895),
            .PADIN(N__57894),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(VDC_SDO),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_174_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_174_iopad (
            .OE(N__57887),
            .DIN(N__57886),
            .DOUT(N__57885),
            .PACKAGEPIN(ICE_IOT_174));
    defparam ipInertedIOPad_ICE_IOT_174_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_174_preio (
            .PADOEN(N__57887),
            .PADOUT(N__57886),
            .PADIN(N__57885),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_140_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_140_iopad (
            .OE(N__57878),
            .DIN(N__57877),
            .DOUT(N__57876),
            .PACKAGEPIN(ICE_IOR_140));
    defparam ipInertedIOPad_ICE_IOR_140_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_140_preio (
            .PADOEN(N__57878),
            .PADOUT(N__57877),
            .PADIN(N__57876),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOB_96_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOB_96_iopad (
            .OE(N__57869),
            .DIN(N__57868),
            .DOUT(N__57867),
            .PACKAGEPIN(ICE_IOB_96));
    defparam ipInertedIOPad_ICE_IOB_96_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_96_preio (
            .PADOEN(N__57869),
            .PADOUT(N__57868),
            .PADIN(N__57867),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_CONT_SD_iopad (
            .OE(N__57860),
            .DIN(N__57859),
            .DOUT(N__57858),
            .PACKAGEPIN(CONT_SD));
    defparam ipInertedIOPad_CONT_SD_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_CONT_SD_preio (
            .PADOEN(N__57860),
            .PADOUT(N__57859),
            .PADIN(N__57858),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__50239),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_AC_ADC_SYNC_iopad (
            .OE(N__57851),
            .DIN(N__57850),
            .DOUT(N__57849),
            .PACKAGEPIN(AC_ADC_SYNC));
    defparam ipInertedIOPad_AC_ADC_SYNC_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_AC_ADC_SYNC_preio (
            .PADOEN(N__57851),
            .PADOUT(N__57850),
            .PADIN(N__57849),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__26242),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SELIRNG1_iopad (
            .OE(N__57842),
            .DIN(N__57841),
            .DOUT(N__57840),
            .PACKAGEPIN(SELIRNG1));
    defparam ipInertedIOPad_SELIRNG1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_SELIRNG1_preio (
            .PADOEN(N__57842),
            .PADOUT(N__57841),
            .PADIN(N__57840),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__45511),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_12B_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_12B_iopad (
            .OE(N__57833),
            .DIN(N__57832),
            .DOUT(N__57831),
            .PACKAGEPIN(ICE_IOL_12B));
    defparam ipInertedIOPad_ICE_IOL_12B_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_12B_preio (
            .PADOEN(N__57833),
            .PADOUT(N__57832),
            .PADIN(N__57831),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_160_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_160_iopad (
            .OE(N__57824),
            .DIN(N__57823),
            .DOUT(N__57822),
            .PACKAGEPIN(ICE_IOR_160));
    defparam ipInertedIOPad_ICE_IOR_160_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_160_preio (
            .PADOEN(N__57824),
            .PADOUT(N__57823),
            .PADIN(N__57822),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_136_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_136_iopad (
            .OE(N__57815),
            .DIN(N__57814),
            .DOUT(N__57813),
            .PACKAGEPIN(ICE_IOR_136));
    defparam ipInertedIOPad_ICE_IOR_136_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_136_preio (
            .PADOEN(N__57815),
            .PADOUT(N__57814),
            .PADIN(N__57813),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_MCLK1_iopad (
            .OE(N__57806),
            .DIN(N__57805),
            .DOUT(N__57804),
            .PACKAGEPIN(DDS_MCLK1));
    defparam ipInertedIOPad_DDS_MCLK1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_MCLK1_preio (
            .PADOEN(N__57806),
            .PADOUT(N__57805),
            .PADIN(N__57804),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__21649),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_198_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_198_iopad (
            .OE(N__57797),
            .DIN(N__57796),
            .DOUT(N__57795),
            .PACKAGEPIN(ICE_IOT_198));
    defparam ipInertedIOPad_ICE_IOT_198_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_198_preio (
            .PADOEN(N__57797),
            .PADOUT(N__57796),
            .PADIN(N__57795),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_173_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_173_iopad (
            .OE(N__57788),
            .DIN(N__57787),
            .DOUT(N__57786),
            .PACKAGEPIN(ICE_IOT_173));
    defparam ipInertedIOPad_ICE_IOT_173_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_173_preio (
            .PADOEN(N__57788),
            .PADOUT(N__57787),
            .PADIN(N__57786),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_DRDY_iopad (
            .OE(N__57779),
            .DIN(N__57778),
            .DOUT(N__57777),
            .PACKAGEPIN(IAC_DRDY));
    defparam ipInertedIOPad_IAC_DRDY_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_IAC_DRDY_preio (
            .PADOEN(N__57779),
            .PADOUT(N__57778),
            .PADIN(N__57777),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(IAC_DRDY),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_178_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_178_iopad (
            .OE(N__57770),
            .DIN(N__57769),
            .DOUT(N__57768),
            .PACKAGEPIN(ICE_IOT_178));
    defparam ipInertedIOPad_ICE_IOT_178_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_178_preio (
            .PADOEN(N__57770),
            .PADOUT(N__57769),
            .PADIN(N__57768),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_138_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_138_iopad (
            .OE(N__57761),
            .DIN(N__57760),
            .DOUT(N__57759),
            .PACKAGEPIN(ICE_IOR_138));
    defparam ipInertedIOPad_ICE_IOR_138_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_138_preio (
            .PADOEN(N__57761),
            .PADOUT(N__57760),
            .PADIN(N__57759),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_120_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_120_iopad (
            .OE(N__57752),
            .DIN(N__57751),
            .DOUT(N__57750),
            .PACKAGEPIN(ICE_IOR_120));
    defparam ipInertedIOPad_ICE_IOR_120_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_120_preio (
            .PADOEN(N__57752),
            .PADOUT(N__57751),
            .PADIN(N__57750),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_FLT0_iopad (
            .OE(N__57743),
            .DIN(N__57742),
            .DOUT(N__57741),
            .PACKAGEPIN(IAC_FLT0));
    defparam ipInertedIOPad_IAC_FLT0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_FLT0_preio (
            .PADOEN(N__57743),
            .PADOUT(N__57742),
            .PADIN(N__57741),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__28027),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_SCK1_iopad (
            .OE(N__57734),
            .DIN(N__57733),
            .DOUT(N__57732),
            .PACKAGEPIN(DDS_SCK1));
    defparam ipInertedIOPad_DDS_SCK1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_SCK1_preio (
            .PADOEN(N__57734),
            .PADOUT(N__57733),
            .PADIN(N__57732),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__21613),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    InMux I__14461 (
            .O(N__57715),
            .I(N__57711));
    InMux I__14460 (
            .O(N__57714),
            .I(N__57708));
    LocalMux I__14459 (
            .O(N__57711),
            .I(N__57705));
    LocalMux I__14458 (
            .O(N__57708),
            .I(dds0_mclkcnt_0));
    Odrv4 I__14457 (
            .O(N__57705),
            .I(dds0_mclkcnt_0));
    InMux I__14456 (
            .O(N__57700),
            .I(bfn_22_11_0_));
    CascadeMux I__14455 (
            .O(N__57697),
            .I(N__57694));
    InMux I__14454 (
            .O(N__57694),
            .I(N__57690));
    InMux I__14453 (
            .O(N__57693),
            .I(N__57687));
    LocalMux I__14452 (
            .O(N__57690),
            .I(N__57684));
    LocalMux I__14451 (
            .O(N__57687),
            .I(N__57679));
    Span4Mux_h I__14450 (
            .O(N__57684),
            .I(N__57679));
    Odrv4 I__14449 (
            .O(N__57679),
            .I(dds0_mclkcnt_1));
    InMux I__14448 (
            .O(N__57676),
            .I(n19440));
    CascadeMux I__14447 (
            .O(N__57673),
            .I(N__57670));
    InMux I__14446 (
            .O(N__57670),
            .I(N__57666));
    InMux I__14445 (
            .O(N__57669),
            .I(N__57663));
    LocalMux I__14444 (
            .O(N__57666),
            .I(N__57660));
    LocalMux I__14443 (
            .O(N__57663),
            .I(dds0_mclkcnt_2));
    Odrv4 I__14442 (
            .O(N__57660),
            .I(dds0_mclkcnt_2));
    InMux I__14441 (
            .O(N__57655),
            .I(n19441));
    InMux I__14440 (
            .O(N__57652),
            .I(N__57648));
    InMux I__14439 (
            .O(N__57651),
            .I(N__57645));
    LocalMux I__14438 (
            .O(N__57648),
            .I(N__57642));
    LocalMux I__14437 (
            .O(N__57645),
            .I(dds0_mclkcnt_3));
    Odrv12 I__14436 (
            .O(N__57642),
            .I(dds0_mclkcnt_3));
    InMux I__14435 (
            .O(N__57637),
            .I(n19442));
    InMux I__14434 (
            .O(N__57634),
            .I(N__57630));
    InMux I__14433 (
            .O(N__57633),
            .I(N__57627));
    LocalMux I__14432 (
            .O(N__57630),
            .I(N__57624));
    LocalMux I__14431 (
            .O(N__57627),
            .I(dds0_mclkcnt_4));
    Odrv4 I__14430 (
            .O(N__57624),
            .I(dds0_mclkcnt_4));
    InMux I__14429 (
            .O(N__57619),
            .I(n19443));
    InMux I__14428 (
            .O(N__57616),
            .I(N__57612));
    InMux I__14427 (
            .O(N__57615),
            .I(N__57609));
    LocalMux I__14426 (
            .O(N__57612),
            .I(N__57606));
    LocalMux I__14425 (
            .O(N__57609),
            .I(dds0_mclkcnt_5));
    Odrv4 I__14424 (
            .O(N__57606),
            .I(dds0_mclkcnt_5));
    InMux I__14423 (
            .O(N__57601),
            .I(n19444));
    InMux I__14422 (
            .O(N__57598),
            .I(N__57595));
    LocalMux I__14421 (
            .O(N__57595),
            .I(N__57592));
    Odrv4 I__14420 (
            .O(N__57592),
            .I(n10));
    InMux I__14419 (
            .O(N__57589),
            .I(N__57583));
    InMux I__14418 (
            .O(N__57588),
            .I(N__57583));
    LocalMux I__14417 (
            .O(N__57583),
            .I(N__57580));
    Span4Mux_h I__14416 (
            .O(N__57580),
            .I(N__57577));
    Odrv4 I__14415 (
            .O(N__57577),
            .I(dds0_mclkcnt_6));
    InMux I__14414 (
            .O(N__57574),
            .I(n19445));
    InMux I__14413 (
            .O(N__57571),
            .I(n19446));
    InMux I__14412 (
            .O(N__57568),
            .I(N__57564));
    InMux I__14411 (
            .O(N__57567),
            .I(N__57561));
    LocalMux I__14410 (
            .O(N__57564),
            .I(N__57558));
    LocalMux I__14409 (
            .O(N__57561),
            .I(dds0_mclkcnt_7));
    Odrv4 I__14408 (
            .O(N__57558),
            .I(dds0_mclkcnt_7));
    InMux I__14407 (
            .O(N__57553),
            .I(N__57544));
    InMux I__14406 (
            .O(N__57552),
            .I(N__57526));
    InMux I__14405 (
            .O(N__57551),
            .I(N__57526));
    InMux I__14404 (
            .O(N__57550),
            .I(N__57516));
    InMux I__14403 (
            .O(N__57549),
            .I(N__57516));
    InMux I__14402 (
            .O(N__57548),
            .I(N__57513));
    InMux I__14401 (
            .O(N__57547),
            .I(N__57510));
    LocalMux I__14400 (
            .O(N__57544),
            .I(N__57507));
    InMux I__14399 (
            .O(N__57543),
            .I(N__57504));
    InMux I__14398 (
            .O(N__57542),
            .I(N__57497));
    InMux I__14397 (
            .O(N__57541),
            .I(N__57497));
    InMux I__14396 (
            .O(N__57540),
            .I(N__57494));
    InMux I__14395 (
            .O(N__57539),
            .I(N__57490));
    CascadeMux I__14394 (
            .O(N__57538),
            .I(N__57486));
    InMux I__14393 (
            .O(N__57537),
            .I(N__57472));
    InMux I__14392 (
            .O(N__57536),
            .I(N__57472));
    InMux I__14391 (
            .O(N__57535),
            .I(N__57472));
    InMux I__14390 (
            .O(N__57534),
            .I(N__57469));
    CascadeMux I__14389 (
            .O(N__57533),
            .I(N__57466));
    InMux I__14388 (
            .O(N__57532),
            .I(N__57459));
    InMux I__14387 (
            .O(N__57531),
            .I(N__57456));
    LocalMux I__14386 (
            .O(N__57526),
            .I(N__57453));
    InMux I__14385 (
            .O(N__57525),
            .I(N__57450));
    CascadeMux I__14384 (
            .O(N__57524),
            .I(N__57437));
    InMux I__14383 (
            .O(N__57523),
            .I(N__57433));
    InMux I__14382 (
            .O(N__57522),
            .I(N__57430));
    InMux I__14381 (
            .O(N__57521),
            .I(N__57427));
    LocalMux I__14380 (
            .O(N__57516),
            .I(N__57422));
    LocalMux I__14379 (
            .O(N__57513),
            .I(N__57422));
    LocalMux I__14378 (
            .O(N__57510),
            .I(N__57419));
    Span4Mux_h I__14377 (
            .O(N__57507),
            .I(N__57414));
    LocalMux I__14376 (
            .O(N__57504),
            .I(N__57414));
    InMux I__14375 (
            .O(N__57503),
            .I(N__57411));
    InMux I__14374 (
            .O(N__57502),
            .I(N__57404));
    LocalMux I__14373 (
            .O(N__57497),
            .I(N__57399));
    LocalMux I__14372 (
            .O(N__57494),
            .I(N__57399));
    InMux I__14371 (
            .O(N__57493),
            .I(N__57396));
    LocalMux I__14370 (
            .O(N__57490),
            .I(N__57383));
    InMux I__14369 (
            .O(N__57489),
            .I(N__57380));
    InMux I__14368 (
            .O(N__57486),
            .I(N__57377));
    InMux I__14367 (
            .O(N__57485),
            .I(N__57374));
    InMux I__14366 (
            .O(N__57484),
            .I(N__57371));
    InMux I__14365 (
            .O(N__57483),
            .I(N__57367));
    InMux I__14364 (
            .O(N__57482),
            .I(N__57364));
    InMux I__14363 (
            .O(N__57481),
            .I(N__57359));
    InMux I__14362 (
            .O(N__57480),
            .I(N__57359));
    InMux I__14361 (
            .O(N__57479),
            .I(N__57356));
    LocalMux I__14360 (
            .O(N__57472),
            .I(N__57353));
    LocalMux I__14359 (
            .O(N__57469),
            .I(N__57350));
    InMux I__14358 (
            .O(N__57466),
            .I(N__57347));
    CascadeMux I__14357 (
            .O(N__57465),
            .I(N__57342));
    InMux I__14356 (
            .O(N__57464),
            .I(N__57334));
    InMux I__14355 (
            .O(N__57463),
            .I(N__57334));
    InMux I__14354 (
            .O(N__57462),
            .I(N__57334));
    LocalMux I__14353 (
            .O(N__57459),
            .I(N__57331));
    LocalMux I__14352 (
            .O(N__57456),
            .I(N__57328));
    Span4Mux_v I__14351 (
            .O(N__57453),
            .I(N__57323));
    LocalMux I__14350 (
            .O(N__57450),
            .I(N__57323));
    InMux I__14349 (
            .O(N__57449),
            .I(N__57318));
    InMux I__14348 (
            .O(N__57448),
            .I(N__57318));
    CascadeMux I__14347 (
            .O(N__57447),
            .I(N__57315));
    InMux I__14346 (
            .O(N__57446),
            .I(N__57312));
    InMux I__14345 (
            .O(N__57445),
            .I(N__57305));
    InMux I__14344 (
            .O(N__57444),
            .I(N__57305));
    InMux I__14343 (
            .O(N__57443),
            .I(N__57300));
    InMux I__14342 (
            .O(N__57442),
            .I(N__57300));
    InMux I__14341 (
            .O(N__57441),
            .I(N__57297));
    InMux I__14340 (
            .O(N__57440),
            .I(N__57294));
    InMux I__14339 (
            .O(N__57437),
            .I(N__57291));
    InMux I__14338 (
            .O(N__57436),
            .I(N__57288));
    LocalMux I__14337 (
            .O(N__57433),
            .I(N__57279));
    LocalMux I__14336 (
            .O(N__57430),
            .I(N__57279));
    LocalMux I__14335 (
            .O(N__57427),
            .I(N__57279));
    Span4Mux_h I__14334 (
            .O(N__57422),
            .I(N__57279));
    Span4Mux_v I__14333 (
            .O(N__57419),
            .I(N__57274));
    Span4Mux_h I__14332 (
            .O(N__57414),
            .I(N__57274));
    LocalMux I__14331 (
            .O(N__57411),
            .I(N__57271));
    InMux I__14330 (
            .O(N__57410),
            .I(N__57262));
    InMux I__14329 (
            .O(N__57409),
            .I(N__57262));
    InMux I__14328 (
            .O(N__57408),
            .I(N__57262));
    InMux I__14327 (
            .O(N__57407),
            .I(N__57262));
    LocalMux I__14326 (
            .O(N__57404),
            .I(N__57259));
    Span4Mux_v I__14325 (
            .O(N__57399),
            .I(N__57254));
    LocalMux I__14324 (
            .O(N__57396),
            .I(N__57254));
    InMux I__14323 (
            .O(N__57395),
            .I(N__57251));
    InMux I__14322 (
            .O(N__57394),
            .I(N__57243));
    InMux I__14321 (
            .O(N__57393),
            .I(N__57243));
    InMux I__14320 (
            .O(N__57392),
            .I(N__57243));
    InMux I__14319 (
            .O(N__57391),
            .I(N__57238));
    InMux I__14318 (
            .O(N__57390),
            .I(N__57233));
    InMux I__14317 (
            .O(N__57389),
            .I(N__57233));
    InMux I__14316 (
            .O(N__57388),
            .I(N__57230));
    InMux I__14315 (
            .O(N__57387),
            .I(N__57225));
    InMux I__14314 (
            .O(N__57386),
            .I(N__57225));
    Span4Mux_h I__14313 (
            .O(N__57383),
            .I(N__57220));
    LocalMux I__14312 (
            .O(N__57380),
            .I(N__57220));
    LocalMux I__14311 (
            .O(N__57377),
            .I(N__57215));
    LocalMux I__14310 (
            .O(N__57374),
            .I(N__57215));
    LocalMux I__14309 (
            .O(N__57371),
            .I(N__57212));
    InMux I__14308 (
            .O(N__57370),
            .I(N__57209));
    LocalMux I__14307 (
            .O(N__57367),
            .I(N__57206));
    LocalMux I__14306 (
            .O(N__57364),
            .I(N__57193));
    LocalMux I__14305 (
            .O(N__57359),
            .I(N__57193));
    LocalMux I__14304 (
            .O(N__57356),
            .I(N__57193));
    Span4Mux_h I__14303 (
            .O(N__57353),
            .I(N__57193));
    Span4Mux_v I__14302 (
            .O(N__57350),
            .I(N__57193));
    LocalMux I__14301 (
            .O(N__57347),
            .I(N__57193));
    InMux I__14300 (
            .O(N__57346),
            .I(N__57172));
    InMux I__14299 (
            .O(N__57345),
            .I(N__57172));
    InMux I__14298 (
            .O(N__57342),
            .I(N__57172));
    InMux I__14297 (
            .O(N__57341),
            .I(N__57172));
    LocalMux I__14296 (
            .O(N__57334),
            .I(N__57163));
    Span4Mux_h I__14295 (
            .O(N__57331),
            .I(N__57163));
    Span4Mux_v I__14294 (
            .O(N__57328),
            .I(N__57163));
    Span4Mux_h I__14293 (
            .O(N__57323),
            .I(N__57163));
    LocalMux I__14292 (
            .O(N__57318),
            .I(N__57160));
    InMux I__14291 (
            .O(N__57315),
            .I(N__57157));
    LocalMux I__14290 (
            .O(N__57312),
            .I(N__57154));
    InMux I__14289 (
            .O(N__57311),
            .I(N__57149));
    InMux I__14288 (
            .O(N__57310),
            .I(N__57149));
    LocalMux I__14287 (
            .O(N__57305),
            .I(N__57142));
    LocalMux I__14286 (
            .O(N__57300),
            .I(N__57142));
    LocalMux I__14285 (
            .O(N__57297),
            .I(N__57142));
    LocalMux I__14284 (
            .O(N__57294),
            .I(N__57135));
    LocalMux I__14283 (
            .O(N__57291),
            .I(N__57135));
    LocalMux I__14282 (
            .O(N__57288),
            .I(N__57135));
    Span4Mux_v I__14281 (
            .O(N__57279),
            .I(N__57126));
    Span4Mux_h I__14280 (
            .O(N__57274),
            .I(N__57126));
    Span4Mux_h I__14279 (
            .O(N__57271),
            .I(N__57126));
    LocalMux I__14278 (
            .O(N__57262),
            .I(N__57126));
    Sp12to4 I__14277 (
            .O(N__57259),
            .I(N__57119));
    Sp12to4 I__14276 (
            .O(N__57254),
            .I(N__57119));
    LocalMux I__14275 (
            .O(N__57251),
            .I(N__57119));
    InMux I__14274 (
            .O(N__57250),
            .I(N__57116));
    LocalMux I__14273 (
            .O(N__57243),
            .I(N__57113));
    InMux I__14272 (
            .O(N__57242),
            .I(N__57108));
    InMux I__14271 (
            .O(N__57241),
            .I(N__57108));
    LocalMux I__14270 (
            .O(N__57238),
            .I(N__57091));
    LocalMux I__14269 (
            .O(N__57233),
            .I(N__57091));
    LocalMux I__14268 (
            .O(N__57230),
            .I(N__57091));
    LocalMux I__14267 (
            .O(N__57225),
            .I(N__57091));
    Span4Mux_h I__14266 (
            .O(N__57220),
            .I(N__57091));
    Span4Mux_h I__14265 (
            .O(N__57215),
            .I(N__57091));
    Span4Mux_v I__14264 (
            .O(N__57212),
            .I(N__57091));
    LocalMux I__14263 (
            .O(N__57209),
            .I(N__57091));
    Span4Mux_v I__14262 (
            .O(N__57206),
            .I(N__57086));
    Span4Mux_h I__14261 (
            .O(N__57193),
            .I(N__57086));
    InMux I__14260 (
            .O(N__57192),
            .I(N__57081));
    InMux I__14259 (
            .O(N__57191),
            .I(N__57081));
    InMux I__14258 (
            .O(N__57190),
            .I(N__57074));
    InMux I__14257 (
            .O(N__57189),
            .I(N__57074));
    InMux I__14256 (
            .O(N__57188),
            .I(N__57074));
    InMux I__14255 (
            .O(N__57187),
            .I(N__57071));
    InMux I__14254 (
            .O(N__57186),
            .I(N__57064));
    InMux I__14253 (
            .O(N__57185),
            .I(N__57064));
    InMux I__14252 (
            .O(N__57184),
            .I(N__57064));
    InMux I__14251 (
            .O(N__57183),
            .I(N__57061));
    InMux I__14250 (
            .O(N__57182),
            .I(N__57058));
    InMux I__14249 (
            .O(N__57181),
            .I(N__57055));
    LocalMux I__14248 (
            .O(N__57172),
            .I(N__57050));
    Span4Mux_v I__14247 (
            .O(N__57163),
            .I(N__57050));
    Span12Mux_v I__14246 (
            .O(N__57160),
            .I(N__57045));
    LocalMux I__14245 (
            .O(N__57157),
            .I(N__57045));
    Span4Mux_v I__14244 (
            .O(N__57154),
            .I(N__57040));
    LocalMux I__14243 (
            .O(N__57149),
            .I(N__57040));
    Span4Mux_h I__14242 (
            .O(N__57142),
            .I(N__57037));
    Span4Mux_v I__14241 (
            .O(N__57135),
            .I(N__57032));
    Span4Mux_h I__14240 (
            .O(N__57126),
            .I(N__57032));
    Span12Mux_h I__14239 (
            .O(N__57119),
            .I(N__57029));
    LocalMux I__14238 (
            .O(N__57116),
            .I(N__57018));
    Span4Mux_h I__14237 (
            .O(N__57113),
            .I(N__57018));
    LocalMux I__14236 (
            .O(N__57108),
            .I(N__57018));
    Span4Mux_v I__14235 (
            .O(N__57091),
            .I(N__57018));
    Span4Mux_h I__14234 (
            .O(N__57086),
            .I(N__57018));
    LocalMux I__14233 (
            .O(N__57081),
            .I(comm_cmd_1));
    LocalMux I__14232 (
            .O(N__57074),
            .I(comm_cmd_1));
    LocalMux I__14231 (
            .O(N__57071),
            .I(comm_cmd_1));
    LocalMux I__14230 (
            .O(N__57064),
            .I(comm_cmd_1));
    LocalMux I__14229 (
            .O(N__57061),
            .I(comm_cmd_1));
    LocalMux I__14228 (
            .O(N__57058),
            .I(comm_cmd_1));
    LocalMux I__14227 (
            .O(N__57055),
            .I(comm_cmd_1));
    Odrv4 I__14226 (
            .O(N__57050),
            .I(comm_cmd_1));
    Odrv12 I__14225 (
            .O(N__57045),
            .I(comm_cmd_1));
    Odrv4 I__14224 (
            .O(N__57040),
            .I(comm_cmd_1));
    Odrv4 I__14223 (
            .O(N__57037),
            .I(comm_cmd_1));
    Odrv4 I__14222 (
            .O(N__57032),
            .I(comm_cmd_1));
    Odrv12 I__14221 (
            .O(N__57029),
            .I(comm_cmd_1));
    Odrv4 I__14220 (
            .O(N__57018),
            .I(comm_cmd_1));
    InMux I__14219 (
            .O(N__56989),
            .I(N__56985));
    InMux I__14218 (
            .O(N__56988),
            .I(N__56979));
    LocalMux I__14217 (
            .O(N__56985),
            .I(N__56974));
    InMux I__14216 (
            .O(N__56984),
            .I(N__56969));
    InMux I__14215 (
            .O(N__56983),
            .I(N__56969));
    InMux I__14214 (
            .O(N__56982),
            .I(N__56961));
    LocalMux I__14213 (
            .O(N__56979),
            .I(N__56946));
    InMux I__14212 (
            .O(N__56978),
            .I(N__56942));
    CascadeMux I__14211 (
            .O(N__56977),
            .I(N__56935));
    Span4Mux_h I__14210 (
            .O(N__56974),
            .I(N__56922));
    LocalMux I__14209 (
            .O(N__56969),
            .I(N__56922));
    InMux I__14208 (
            .O(N__56968),
            .I(N__56918));
    InMux I__14207 (
            .O(N__56967),
            .I(N__56915));
    InMux I__14206 (
            .O(N__56966),
            .I(N__56898));
    InMux I__14205 (
            .O(N__56965),
            .I(N__56894));
    InMux I__14204 (
            .O(N__56964),
            .I(N__56891));
    LocalMux I__14203 (
            .O(N__56961),
            .I(N__56880));
    InMux I__14202 (
            .O(N__56960),
            .I(N__56875));
    InMux I__14201 (
            .O(N__56959),
            .I(N__56875));
    InMux I__14200 (
            .O(N__56958),
            .I(N__56868));
    InMux I__14199 (
            .O(N__56957),
            .I(N__56868));
    InMux I__14198 (
            .O(N__56956),
            .I(N__56868));
    InMux I__14197 (
            .O(N__56955),
            .I(N__56860));
    InMux I__14196 (
            .O(N__56954),
            .I(N__56860));
    InMux I__14195 (
            .O(N__56953),
            .I(N__56855));
    InMux I__14194 (
            .O(N__56952),
            .I(N__56855));
    InMux I__14193 (
            .O(N__56951),
            .I(N__56848));
    InMux I__14192 (
            .O(N__56950),
            .I(N__56848));
    InMux I__14191 (
            .O(N__56949),
            .I(N__56848));
    Span4Mux_h I__14190 (
            .O(N__56946),
            .I(N__56845));
    InMux I__14189 (
            .O(N__56945),
            .I(N__56842));
    LocalMux I__14188 (
            .O(N__56942),
            .I(N__56837));
    InMux I__14187 (
            .O(N__56941),
            .I(N__56834));
    InMux I__14186 (
            .O(N__56940),
            .I(N__56824));
    InMux I__14185 (
            .O(N__56939),
            .I(N__56824));
    InMux I__14184 (
            .O(N__56938),
            .I(N__56824));
    InMux I__14183 (
            .O(N__56935),
            .I(N__56811));
    InMux I__14182 (
            .O(N__56934),
            .I(N__56811));
    InMux I__14181 (
            .O(N__56933),
            .I(N__56811));
    InMux I__14180 (
            .O(N__56932),
            .I(N__56811));
    InMux I__14179 (
            .O(N__56931),
            .I(N__56811));
    InMux I__14178 (
            .O(N__56930),
            .I(N__56811));
    InMux I__14177 (
            .O(N__56929),
            .I(N__56804));
    InMux I__14176 (
            .O(N__56928),
            .I(N__56804));
    InMux I__14175 (
            .O(N__56927),
            .I(N__56804));
    Span4Mux_v I__14174 (
            .O(N__56922),
            .I(N__56794));
    InMux I__14173 (
            .O(N__56921),
            .I(N__56791));
    LocalMux I__14172 (
            .O(N__56918),
            .I(N__56786));
    LocalMux I__14171 (
            .O(N__56915),
            .I(N__56786));
    InMux I__14170 (
            .O(N__56914),
            .I(N__56781));
    InMux I__14169 (
            .O(N__56913),
            .I(N__56781));
    InMux I__14168 (
            .O(N__56912),
            .I(N__56778));
    InMux I__14167 (
            .O(N__56911),
            .I(N__56775));
    InMux I__14166 (
            .O(N__56910),
            .I(N__56772));
    InMux I__14165 (
            .O(N__56909),
            .I(N__56763));
    InMux I__14164 (
            .O(N__56908),
            .I(N__56763));
    InMux I__14163 (
            .O(N__56907),
            .I(N__56763));
    InMux I__14162 (
            .O(N__56906),
            .I(N__56763));
    InMux I__14161 (
            .O(N__56905),
            .I(N__56760));
    InMux I__14160 (
            .O(N__56904),
            .I(N__56757));
    InMux I__14159 (
            .O(N__56903),
            .I(N__56754));
    InMux I__14158 (
            .O(N__56902),
            .I(N__56749));
    InMux I__14157 (
            .O(N__56901),
            .I(N__56749));
    LocalMux I__14156 (
            .O(N__56898),
            .I(N__56746));
    InMux I__14155 (
            .O(N__56897),
            .I(N__56743));
    LocalMux I__14154 (
            .O(N__56894),
            .I(N__56738));
    LocalMux I__14153 (
            .O(N__56891),
            .I(N__56738));
    InMux I__14152 (
            .O(N__56890),
            .I(N__56733));
    InMux I__14151 (
            .O(N__56889),
            .I(N__56733));
    InMux I__14150 (
            .O(N__56888),
            .I(N__56730));
    InMux I__14149 (
            .O(N__56887),
            .I(N__56727));
    InMux I__14148 (
            .O(N__56886),
            .I(N__56722));
    InMux I__14147 (
            .O(N__56885),
            .I(N__56717));
    InMux I__14146 (
            .O(N__56884),
            .I(N__56717));
    InMux I__14145 (
            .O(N__56883),
            .I(N__56714));
    Span4Mux_h I__14144 (
            .O(N__56880),
            .I(N__56707));
    LocalMux I__14143 (
            .O(N__56875),
            .I(N__56707));
    LocalMux I__14142 (
            .O(N__56868),
            .I(N__56707));
    InMux I__14141 (
            .O(N__56867),
            .I(N__56700));
    InMux I__14140 (
            .O(N__56866),
            .I(N__56700));
    InMux I__14139 (
            .O(N__56865),
            .I(N__56700));
    LocalMux I__14138 (
            .O(N__56860),
            .I(N__56695));
    LocalMux I__14137 (
            .O(N__56855),
            .I(N__56690));
    LocalMux I__14136 (
            .O(N__56848),
            .I(N__56687));
    Span4Mux_v I__14135 (
            .O(N__56845),
            .I(N__56678));
    LocalMux I__14134 (
            .O(N__56842),
            .I(N__56678));
    InMux I__14133 (
            .O(N__56841),
            .I(N__56675));
    InMux I__14132 (
            .O(N__56840),
            .I(N__56672));
    Span4Mux_v I__14131 (
            .O(N__56837),
            .I(N__56667));
    LocalMux I__14130 (
            .O(N__56834),
            .I(N__56667));
    InMux I__14129 (
            .O(N__56833),
            .I(N__56662));
    InMux I__14128 (
            .O(N__56832),
            .I(N__56662));
    InMux I__14127 (
            .O(N__56831),
            .I(N__56659));
    LocalMux I__14126 (
            .O(N__56824),
            .I(N__56652));
    LocalMux I__14125 (
            .O(N__56811),
            .I(N__56652));
    LocalMux I__14124 (
            .O(N__56804),
            .I(N__56652));
    InMux I__14123 (
            .O(N__56803),
            .I(N__56649));
    InMux I__14122 (
            .O(N__56802),
            .I(N__56646));
    InMux I__14121 (
            .O(N__56801),
            .I(N__56643));
    InMux I__14120 (
            .O(N__56800),
            .I(N__56625));
    InMux I__14119 (
            .O(N__56799),
            .I(N__56625));
    InMux I__14118 (
            .O(N__56798),
            .I(N__56625));
    InMux I__14117 (
            .O(N__56797),
            .I(N__56625));
    Span4Mux_h I__14116 (
            .O(N__56794),
            .I(N__56616));
    LocalMux I__14115 (
            .O(N__56791),
            .I(N__56616));
    Span4Mux_v I__14114 (
            .O(N__56786),
            .I(N__56616));
    LocalMux I__14113 (
            .O(N__56781),
            .I(N__56616));
    LocalMux I__14112 (
            .O(N__56778),
            .I(N__56607));
    LocalMux I__14111 (
            .O(N__56775),
            .I(N__56607));
    LocalMux I__14110 (
            .O(N__56772),
            .I(N__56607));
    LocalMux I__14109 (
            .O(N__56763),
            .I(N__56607));
    LocalMux I__14108 (
            .O(N__56760),
            .I(N__56598));
    LocalMux I__14107 (
            .O(N__56757),
            .I(N__56598));
    LocalMux I__14106 (
            .O(N__56754),
            .I(N__56598));
    LocalMux I__14105 (
            .O(N__56749),
            .I(N__56598));
    Span4Mux_v I__14104 (
            .O(N__56746),
            .I(N__56595));
    LocalMux I__14103 (
            .O(N__56743),
            .I(N__56584));
    Span4Mux_v I__14102 (
            .O(N__56738),
            .I(N__56584));
    LocalMux I__14101 (
            .O(N__56733),
            .I(N__56584));
    LocalMux I__14100 (
            .O(N__56730),
            .I(N__56584));
    LocalMux I__14099 (
            .O(N__56727),
            .I(N__56584));
    InMux I__14098 (
            .O(N__56726),
            .I(N__56579));
    InMux I__14097 (
            .O(N__56725),
            .I(N__56579));
    LocalMux I__14096 (
            .O(N__56722),
            .I(N__56568));
    LocalMux I__14095 (
            .O(N__56717),
            .I(N__56568));
    LocalMux I__14094 (
            .O(N__56714),
            .I(N__56568));
    Span4Mux_h I__14093 (
            .O(N__56707),
            .I(N__56568));
    LocalMux I__14092 (
            .O(N__56700),
            .I(N__56568));
    CascadeMux I__14091 (
            .O(N__56699),
            .I(N__56564));
    InMux I__14090 (
            .O(N__56698),
            .I(N__56559));
    Span4Mux_h I__14089 (
            .O(N__56695),
            .I(N__56556));
    InMux I__14088 (
            .O(N__56694),
            .I(N__56551));
    InMux I__14087 (
            .O(N__56693),
            .I(N__56551));
    Span4Mux_h I__14086 (
            .O(N__56690),
            .I(N__56546));
    Span4Mux_h I__14085 (
            .O(N__56687),
            .I(N__56546));
    InMux I__14084 (
            .O(N__56686),
            .I(N__56543));
    InMux I__14083 (
            .O(N__56685),
            .I(N__56536));
    InMux I__14082 (
            .O(N__56684),
            .I(N__56536));
    InMux I__14081 (
            .O(N__56683),
            .I(N__56536));
    Span4Mux_h I__14080 (
            .O(N__56678),
            .I(N__56533));
    LocalMux I__14079 (
            .O(N__56675),
            .I(N__56528));
    LocalMux I__14078 (
            .O(N__56672),
            .I(N__56528));
    Span4Mux_h I__14077 (
            .O(N__56667),
            .I(N__56517));
    LocalMux I__14076 (
            .O(N__56662),
            .I(N__56517));
    LocalMux I__14075 (
            .O(N__56659),
            .I(N__56517));
    Span4Mux_v I__14074 (
            .O(N__56652),
            .I(N__56517));
    LocalMux I__14073 (
            .O(N__56649),
            .I(N__56517));
    LocalMux I__14072 (
            .O(N__56646),
            .I(N__56512));
    LocalMux I__14071 (
            .O(N__56643),
            .I(N__56512));
    InMux I__14070 (
            .O(N__56642),
            .I(N__56509));
    InMux I__14069 (
            .O(N__56641),
            .I(N__56502));
    InMux I__14068 (
            .O(N__56640),
            .I(N__56502));
    InMux I__14067 (
            .O(N__56639),
            .I(N__56502));
    InMux I__14066 (
            .O(N__56638),
            .I(N__56499));
    InMux I__14065 (
            .O(N__56637),
            .I(N__56490));
    InMux I__14064 (
            .O(N__56636),
            .I(N__56490));
    InMux I__14063 (
            .O(N__56635),
            .I(N__56490));
    InMux I__14062 (
            .O(N__56634),
            .I(N__56490));
    LocalMux I__14061 (
            .O(N__56625),
            .I(N__56487));
    Span4Mux_v I__14060 (
            .O(N__56616),
            .I(N__56480));
    Span4Mux_v I__14059 (
            .O(N__56607),
            .I(N__56480));
    Span4Mux_v I__14058 (
            .O(N__56598),
            .I(N__56480));
    Span4Mux_h I__14057 (
            .O(N__56595),
            .I(N__56471));
    Span4Mux_v I__14056 (
            .O(N__56584),
            .I(N__56471));
    LocalMux I__14055 (
            .O(N__56579),
            .I(N__56471));
    Span4Mux_v I__14054 (
            .O(N__56568),
            .I(N__56471));
    InMux I__14053 (
            .O(N__56567),
            .I(N__56462));
    InMux I__14052 (
            .O(N__56564),
            .I(N__56462));
    InMux I__14051 (
            .O(N__56563),
            .I(N__56462));
    InMux I__14050 (
            .O(N__56562),
            .I(N__56462));
    LocalMux I__14049 (
            .O(N__56559),
            .I(N__56451));
    Span4Mux_h I__14048 (
            .O(N__56556),
            .I(N__56451));
    LocalMux I__14047 (
            .O(N__56551),
            .I(N__56451));
    Span4Mux_h I__14046 (
            .O(N__56546),
            .I(N__56451));
    LocalMux I__14045 (
            .O(N__56543),
            .I(N__56451));
    LocalMux I__14044 (
            .O(N__56536),
            .I(N__56446));
    Span4Mux_h I__14043 (
            .O(N__56533),
            .I(N__56446));
    Span4Mux_v I__14042 (
            .O(N__56528),
            .I(N__56441));
    Span4Mux_h I__14041 (
            .O(N__56517),
            .I(N__56441));
    Odrv12 I__14040 (
            .O(N__56512),
            .I(comm_cmd_0));
    LocalMux I__14039 (
            .O(N__56509),
            .I(comm_cmd_0));
    LocalMux I__14038 (
            .O(N__56502),
            .I(comm_cmd_0));
    LocalMux I__14037 (
            .O(N__56499),
            .I(comm_cmd_0));
    LocalMux I__14036 (
            .O(N__56490),
            .I(comm_cmd_0));
    Odrv4 I__14035 (
            .O(N__56487),
            .I(comm_cmd_0));
    Odrv4 I__14034 (
            .O(N__56480),
            .I(comm_cmd_0));
    Odrv4 I__14033 (
            .O(N__56471),
            .I(comm_cmd_0));
    LocalMux I__14032 (
            .O(N__56462),
            .I(comm_cmd_0));
    Odrv4 I__14031 (
            .O(N__56451),
            .I(comm_cmd_0));
    Odrv4 I__14030 (
            .O(N__56446),
            .I(comm_cmd_0));
    Odrv4 I__14029 (
            .O(N__56441),
            .I(comm_cmd_0));
    CascadeMux I__14028 (
            .O(N__56416),
            .I(N__56413));
    InMux I__14027 (
            .O(N__56413),
            .I(N__56410));
    LocalMux I__14026 (
            .O(N__56410),
            .I(N__56407));
    Span4Mux_v I__14025 (
            .O(N__56407),
            .I(N__56404));
    Odrv4 I__14024 (
            .O(N__56404),
            .I(n23_adj_1517));
    InMux I__14023 (
            .O(N__56401),
            .I(N__56398));
    LocalMux I__14022 (
            .O(N__56398),
            .I(N__56394));
    InMux I__14021 (
            .O(N__56397),
            .I(N__56391));
    Span4Mux_h I__14020 (
            .O(N__56394),
            .I(N__56388));
    LocalMux I__14019 (
            .O(N__56391),
            .I(N__56382));
    Span4Mux_v I__14018 (
            .O(N__56388),
            .I(N__56382));
    InMux I__14017 (
            .O(N__56387),
            .I(N__56379));
    Odrv4 I__14016 (
            .O(N__56382),
            .I(req_data_cnt_12));
    LocalMux I__14015 (
            .O(N__56379),
            .I(req_data_cnt_12));
    InMux I__14014 (
            .O(N__56374),
            .I(N__56371));
    LocalMux I__14013 (
            .O(N__56371),
            .I(N__56368));
    Span12Mux_v I__14012 (
            .O(N__56368),
            .I(N__56365));
    Odrv12 I__14011 (
            .O(N__56365),
            .I(n20809));
    InMux I__14010 (
            .O(N__56362),
            .I(N__56359));
    LocalMux I__14009 (
            .O(N__56359),
            .I(N__56356));
    Odrv4 I__14008 (
            .O(N__56356),
            .I(n17415));
    InMux I__14007 (
            .O(N__56353),
            .I(N__56350));
    LocalMux I__14006 (
            .O(N__56350),
            .I(buf_data_iac_4));
    InMux I__14005 (
            .O(N__56347),
            .I(N__56331));
    InMux I__14004 (
            .O(N__56346),
            .I(N__56326));
    InMux I__14003 (
            .O(N__56345),
            .I(N__56326));
    InMux I__14002 (
            .O(N__56344),
            .I(N__56321));
    InMux I__14001 (
            .O(N__56343),
            .I(N__56321));
    CascadeMux I__14000 (
            .O(N__56342),
            .I(N__56318));
    CascadeMux I__13999 (
            .O(N__56341),
            .I(N__56312));
    InMux I__13998 (
            .O(N__56340),
            .I(N__56301));
    InMux I__13997 (
            .O(N__56339),
            .I(N__56301));
    InMux I__13996 (
            .O(N__56338),
            .I(N__56301));
    InMux I__13995 (
            .O(N__56337),
            .I(N__56296));
    InMux I__13994 (
            .O(N__56336),
            .I(N__56296));
    InMux I__13993 (
            .O(N__56335),
            .I(N__56291));
    InMux I__13992 (
            .O(N__56334),
            .I(N__56291));
    LocalMux I__13991 (
            .O(N__56331),
            .I(N__56284));
    LocalMux I__13990 (
            .O(N__56326),
            .I(N__56281));
    LocalMux I__13989 (
            .O(N__56321),
            .I(N__56278));
    InMux I__13988 (
            .O(N__56318),
            .I(N__56275));
    InMux I__13987 (
            .O(N__56317),
            .I(N__56266));
    InMux I__13986 (
            .O(N__56316),
            .I(N__56261));
    InMux I__13985 (
            .O(N__56315),
            .I(N__56253));
    InMux I__13984 (
            .O(N__56312),
            .I(N__56248));
    InMux I__13983 (
            .O(N__56311),
            .I(N__56248));
    InMux I__13982 (
            .O(N__56310),
            .I(N__56245));
    InMux I__13981 (
            .O(N__56309),
            .I(N__56240));
    InMux I__13980 (
            .O(N__56308),
            .I(N__56240));
    LocalMux I__13979 (
            .O(N__56301),
            .I(N__56233));
    LocalMux I__13978 (
            .O(N__56296),
            .I(N__56233));
    LocalMux I__13977 (
            .O(N__56291),
            .I(N__56233));
    InMux I__13976 (
            .O(N__56290),
            .I(N__56228));
    InMux I__13975 (
            .O(N__56289),
            .I(N__56228));
    InMux I__13974 (
            .O(N__56288),
            .I(N__56225));
    InMux I__13973 (
            .O(N__56287),
            .I(N__56222));
    Span4Mux_h I__13972 (
            .O(N__56284),
            .I(N__56213));
    Span4Mux_h I__13971 (
            .O(N__56281),
            .I(N__56213));
    Span4Mux_v I__13970 (
            .O(N__56278),
            .I(N__56213));
    LocalMux I__13969 (
            .O(N__56275),
            .I(N__56213));
    InMux I__13968 (
            .O(N__56274),
            .I(N__56210));
    InMux I__13967 (
            .O(N__56273),
            .I(N__56207));
    InMux I__13966 (
            .O(N__56272),
            .I(N__56204));
    InMux I__13965 (
            .O(N__56271),
            .I(N__56201));
    InMux I__13964 (
            .O(N__56270),
            .I(N__56198));
    InMux I__13963 (
            .O(N__56269),
            .I(N__56195));
    LocalMux I__13962 (
            .O(N__56266),
            .I(N__56192));
    InMux I__13961 (
            .O(N__56265),
            .I(N__56187));
    InMux I__13960 (
            .O(N__56264),
            .I(N__56187));
    LocalMux I__13959 (
            .O(N__56261),
            .I(N__56184));
    InMux I__13958 (
            .O(N__56260),
            .I(N__56181));
    InMux I__13957 (
            .O(N__56259),
            .I(N__56176));
    InMux I__13956 (
            .O(N__56258),
            .I(N__56176));
    InMux I__13955 (
            .O(N__56257),
            .I(N__56173));
    InMux I__13954 (
            .O(N__56256),
            .I(N__56170));
    LocalMux I__13953 (
            .O(N__56253),
            .I(N__56166));
    LocalMux I__13952 (
            .O(N__56248),
            .I(N__56161));
    LocalMux I__13951 (
            .O(N__56245),
            .I(N__56161));
    LocalMux I__13950 (
            .O(N__56240),
            .I(N__56156));
    Span4Mux_v I__13949 (
            .O(N__56233),
            .I(N__56156));
    LocalMux I__13948 (
            .O(N__56228),
            .I(N__56147));
    LocalMux I__13947 (
            .O(N__56225),
            .I(N__56147));
    LocalMux I__13946 (
            .O(N__56222),
            .I(N__56147));
    Span4Mux_h I__13945 (
            .O(N__56213),
            .I(N__56147));
    LocalMux I__13944 (
            .O(N__56210),
            .I(N__56139));
    LocalMux I__13943 (
            .O(N__56207),
            .I(N__56139));
    LocalMux I__13942 (
            .O(N__56204),
            .I(N__56134));
    LocalMux I__13941 (
            .O(N__56201),
            .I(N__56134));
    LocalMux I__13940 (
            .O(N__56198),
            .I(N__56131));
    LocalMux I__13939 (
            .O(N__56195),
            .I(N__56118));
    Span4Mux_v I__13938 (
            .O(N__56192),
            .I(N__56118));
    LocalMux I__13937 (
            .O(N__56187),
            .I(N__56118));
    Span4Mux_h I__13936 (
            .O(N__56184),
            .I(N__56118));
    LocalMux I__13935 (
            .O(N__56181),
            .I(N__56118));
    LocalMux I__13934 (
            .O(N__56176),
            .I(N__56118));
    LocalMux I__13933 (
            .O(N__56173),
            .I(N__56115));
    LocalMux I__13932 (
            .O(N__56170),
            .I(N__56112));
    InMux I__13931 (
            .O(N__56169),
            .I(N__56109));
    Span4Mux_v I__13930 (
            .O(N__56166),
            .I(N__56106));
    Span12Mux_h I__13929 (
            .O(N__56161),
            .I(N__56103));
    Span4Mux_h I__13928 (
            .O(N__56156),
            .I(N__56098));
    Span4Mux_v I__13927 (
            .O(N__56147),
            .I(N__56098));
    InMux I__13926 (
            .O(N__56146),
            .I(N__56091));
    InMux I__13925 (
            .O(N__56145),
            .I(N__56091));
    InMux I__13924 (
            .O(N__56144),
            .I(N__56091));
    Span4Mux_v I__13923 (
            .O(N__56139),
            .I(N__56082));
    Span4Mux_h I__13922 (
            .O(N__56134),
            .I(N__56082));
    Span4Mux_v I__13921 (
            .O(N__56131),
            .I(N__56082));
    Span4Mux_v I__13920 (
            .O(N__56118),
            .I(N__56082));
    Odrv12 I__13919 (
            .O(N__56115),
            .I(comm_cmd_3));
    Odrv4 I__13918 (
            .O(N__56112),
            .I(comm_cmd_3));
    LocalMux I__13917 (
            .O(N__56109),
            .I(comm_cmd_3));
    Odrv4 I__13916 (
            .O(N__56106),
            .I(comm_cmd_3));
    Odrv12 I__13915 (
            .O(N__56103),
            .I(comm_cmd_3));
    Odrv4 I__13914 (
            .O(N__56098),
            .I(comm_cmd_3));
    LocalMux I__13913 (
            .O(N__56091),
            .I(comm_cmd_3));
    Odrv4 I__13912 (
            .O(N__56082),
            .I(comm_cmd_3));
    InMux I__13911 (
            .O(N__56065),
            .I(N__56062));
    LocalMux I__13910 (
            .O(N__56062),
            .I(N__56059));
    Span4Mux_h I__13909 (
            .O(N__56059),
            .I(N__56056));
    Odrv4 I__13908 (
            .O(N__56056),
            .I(n22_adj_1606));
    InMux I__13907 (
            .O(N__56053),
            .I(N__56050));
    LocalMux I__13906 (
            .O(N__56050),
            .I(N__56047));
    Span12Mux_v I__13905 (
            .O(N__56047),
            .I(N__56044));
    Odrv12 I__13904 (
            .O(N__56044),
            .I(n30_adj_1608));
    InMux I__13903 (
            .O(N__56041),
            .I(N__56037));
    InMux I__13902 (
            .O(N__56040),
            .I(N__56034));
    LocalMux I__13901 (
            .O(N__56037),
            .I(N__56031));
    LocalMux I__13900 (
            .O(N__56034),
            .I(N__56019));
    Glb2LocalMux I__13899 (
            .O(N__56031),
            .I(N__55984));
    ClkMux I__13898 (
            .O(N__56030),
            .I(N__55984));
    ClkMux I__13897 (
            .O(N__56029),
            .I(N__55984));
    ClkMux I__13896 (
            .O(N__56028),
            .I(N__55984));
    ClkMux I__13895 (
            .O(N__56027),
            .I(N__55984));
    ClkMux I__13894 (
            .O(N__56026),
            .I(N__55984));
    ClkMux I__13893 (
            .O(N__56025),
            .I(N__55984));
    ClkMux I__13892 (
            .O(N__56024),
            .I(N__55984));
    ClkMux I__13891 (
            .O(N__56023),
            .I(N__55984));
    ClkMux I__13890 (
            .O(N__56022),
            .I(N__55984));
    Glb2LocalMux I__13889 (
            .O(N__56019),
            .I(N__55984));
    ClkMux I__13888 (
            .O(N__56018),
            .I(N__55984));
    ClkMux I__13887 (
            .O(N__56017),
            .I(N__55984));
    ClkMux I__13886 (
            .O(N__56016),
            .I(N__55984));
    ClkMux I__13885 (
            .O(N__56015),
            .I(N__55984));
    GlobalMux I__13884 (
            .O(N__55984),
            .I(clk_16MHz));
    InMux I__13883 (
            .O(N__55981),
            .I(N__55978));
    LocalMux I__13882 (
            .O(N__55978),
            .I(N__55974));
    InMux I__13881 (
            .O(N__55977),
            .I(N__55971));
    Odrv12 I__13880 (
            .O(N__55974),
            .I(dds0_mclk));
    LocalMux I__13879 (
            .O(N__55971),
            .I(dds0_mclk));
    InMux I__13878 (
            .O(N__55966),
            .I(N__55963));
    LocalMux I__13877 (
            .O(N__55963),
            .I(N__55959));
    InMux I__13876 (
            .O(N__55962),
            .I(N__55956));
    Span4Mux_h I__13875 (
            .O(N__55959),
            .I(N__55953));
    LocalMux I__13874 (
            .O(N__55956),
            .I(N__55950));
    Span4Mux_h I__13873 (
            .O(N__55953),
            .I(N__55944));
    Span4Mux_h I__13872 (
            .O(N__55950),
            .I(N__55944));
    InMux I__13871 (
            .O(N__55949),
            .I(N__55941));
    Span4Mux_h I__13870 (
            .O(N__55944),
            .I(N__55938));
    LocalMux I__13869 (
            .O(N__55941),
            .I(buf_control_6));
    Odrv4 I__13868 (
            .O(N__55938),
            .I(buf_control_6));
    IoInMux I__13867 (
            .O(N__55933),
            .I(N__55930));
    LocalMux I__13866 (
            .O(N__55930),
            .I(N__55927));
    Span4Mux_s3_v I__13865 (
            .O(N__55927),
            .I(N__55924));
    Sp12to4 I__13864 (
            .O(N__55924),
            .I(N__55921));
    Span12Mux_s8_h I__13863 (
            .O(N__55921),
            .I(N__55918));
    Odrv12 I__13862 (
            .O(N__55918),
            .I(DDS_MCLK));
    IoInMux I__13861 (
            .O(N__55915),
            .I(N__55912));
    LocalMux I__13860 (
            .O(N__55912),
            .I(N__55909));
    Span4Mux_s1_v I__13859 (
            .O(N__55909),
            .I(N__55906));
    Sp12to4 I__13858 (
            .O(N__55906),
            .I(N__55902));
    CascadeMux I__13857 (
            .O(N__55905),
            .I(N__55899));
    Span12Mux_s8_h I__13856 (
            .O(N__55902),
            .I(N__55896));
    InMux I__13855 (
            .O(N__55899),
            .I(N__55893));
    Odrv12 I__13854 (
            .O(N__55896),
            .I(DDS_SCK));
    LocalMux I__13853 (
            .O(N__55893),
            .I(DDS_SCK));
    CascadeMux I__13852 (
            .O(N__55888),
            .I(N__55875));
    InMux I__13851 (
            .O(N__55887),
            .I(N__55863));
    InMux I__13850 (
            .O(N__55886),
            .I(N__55845));
    InMux I__13849 (
            .O(N__55885),
            .I(N__55845));
    InMux I__13848 (
            .O(N__55884),
            .I(N__55845));
    InMux I__13847 (
            .O(N__55883),
            .I(N__55845));
    InMux I__13846 (
            .O(N__55882),
            .I(N__55845));
    InMux I__13845 (
            .O(N__55881),
            .I(N__55845));
    InMux I__13844 (
            .O(N__55880),
            .I(N__55845));
    InMux I__13843 (
            .O(N__55879),
            .I(N__55840));
    InMux I__13842 (
            .O(N__55878),
            .I(N__55840));
    InMux I__13841 (
            .O(N__55875),
            .I(N__55833));
    InMux I__13840 (
            .O(N__55874),
            .I(N__55833));
    InMux I__13839 (
            .O(N__55873),
            .I(N__55833));
    InMux I__13838 (
            .O(N__55872),
            .I(N__55827));
    InMux I__13837 (
            .O(N__55871),
            .I(N__55827));
    InMux I__13836 (
            .O(N__55870),
            .I(N__55816));
    InMux I__13835 (
            .O(N__55869),
            .I(N__55816));
    InMux I__13834 (
            .O(N__55868),
            .I(N__55816));
    InMux I__13833 (
            .O(N__55867),
            .I(N__55816));
    InMux I__13832 (
            .O(N__55866),
            .I(N__55816));
    LocalMux I__13831 (
            .O(N__55863),
            .I(N__55813));
    InMux I__13830 (
            .O(N__55862),
            .I(N__55810));
    InMux I__13829 (
            .O(N__55861),
            .I(N__55807));
    InMux I__13828 (
            .O(N__55860),
            .I(N__55804));
    LocalMux I__13827 (
            .O(N__55845),
            .I(N__55801));
    LocalMux I__13826 (
            .O(N__55840),
            .I(N__55796));
    LocalMux I__13825 (
            .O(N__55833),
            .I(N__55796));
    InMux I__13824 (
            .O(N__55832),
            .I(N__55792));
    LocalMux I__13823 (
            .O(N__55827),
            .I(N__55787));
    LocalMux I__13822 (
            .O(N__55816),
            .I(N__55787));
    Span4Mux_h I__13821 (
            .O(N__55813),
            .I(N__55784));
    LocalMux I__13820 (
            .O(N__55810),
            .I(N__55781));
    LocalMux I__13819 (
            .O(N__55807),
            .I(N__55776));
    LocalMux I__13818 (
            .O(N__55804),
            .I(N__55776));
    Span4Mux_v I__13817 (
            .O(N__55801),
            .I(N__55771));
    Span4Mux_v I__13816 (
            .O(N__55796),
            .I(N__55771));
    InMux I__13815 (
            .O(N__55795),
            .I(N__55768));
    LocalMux I__13814 (
            .O(N__55792),
            .I(N__55765));
    Span4Mux_v I__13813 (
            .O(N__55787),
            .I(N__55760));
    Span4Mux_h I__13812 (
            .O(N__55784),
            .I(N__55760));
    Span4Mux_v I__13811 (
            .O(N__55781),
            .I(N__55753));
    Span4Mux_v I__13810 (
            .O(N__55776),
            .I(N__55753));
    Span4Mux_h I__13809 (
            .O(N__55771),
            .I(N__55753));
    LocalMux I__13808 (
            .O(N__55768),
            .I(dds_state_2));
    Odrv4 I__13807 (
            .O(N__55765),
            .I(dds_state_2));
    Odrv4 I__13806 (
            .O(N__55760),
            .I(dds_state_2));
    Odrv4 I__13805 (
            .O(N__55753),
            .I(dds_state_2));
    InMux I__13804 (
            .O(N__55744),
            .I(N__55741));
    LocalMux I__13803 (
            .O(N__55741),
            .I(N__55734));
    InMux I__13802 (
            .O(N__55740),
            .I(N__55731));
    InMux I__13801 (
            .O(N__55739),
            .I(N__55728));
    InMux I__13800 (
            .O(N__55738),
            .I(N__55725));
    InMux I__13799 (
            .O(N__55737),
            .I(N__55722));
    Span4Mux_v I__13798 (
            .O(N__55734),
            .I(N__55713));
    LocalMux I__13797 (
            .O(N__55731),
            .I(N__55713));
    LocalMux I__13796 (
            .O(N__55728),
            .I(N__55713));
    LocalMux I__13795 (
            .O(N__55725),
            .I(N__55713));
    LocalMux I__13794 (
            .O(N__55722),
            .I(N__55708));
    Span4Mux_h I__13793 (
            .O(N__55713),
            .I(N__55705));
    InMux I__13792 (
            .O(N__55712),
            .I(N__55700));
    InMux I__13791 (
            .O(N__55711),
            .I(N__55700));
    Span4Mux_v I__13790 (
            .O(N__55708),
            .I(N__55697));
    Span4Mux_h I__13789 (
            .O(N__55705),
            .I(N__55690));
    LocalMux I__13788 (
            .O(N__55700),
            .I(N__55690));
    Span4Mux_h I__13787 (
            .O(N__55697),
            .I(N__55687));
    InMux I__13786 (
            .O(N__55696),
            .I(N__55682));
    InMux I__13785 (
            .O(N__55695),
            .I(N__55682));
    Span4Mux_v I__13784 (
            .O(N__55690),
            .I(N__55679));
    Odrv4 I__13783 (
            .O(N__55687),
            .I(dds_state_0));
    LocalMux I__13782 (
            .O(N__55682),
            .I(dds_state_0));
    Odrv4 I__13781 (
            .O(N__55679),
            .I(dds_state_0));
    CEMux I__13780 (
            .O(N__55672),
            .I(N__55669));
    LocalMux I__13779 (
            .O(N__55669),
            .I(N__55656));
    InMux I__13778 (
            .O(N__55668),
            .I(N__55640));
    InMux I__13777 (
            .O(N__55667),
            .I(N__55640));
    InMux I__13776 (
            .O(N__55666),
            .I(N__55640));
    InMux I__13775 (
            .O(N__55665),
            .I(N__55640));
    InMux I__13774 (
            .O(N__55664),
            .I(N__55640));
    InMux I__13773 (
            .O(N__55663),
            .I(N__55640));
    InMux I__13772 (
            .O(N__55662),
            .I(N__55640));
    InMux I__13771 (
            .O(N__55661),
            .I(N__55635));
    InMux I__13770 (
            .O(N__55660),
            .I(N__55635));
    SRMux I__13769 (
            .O(N__55659),
            .I(N__55623));
    Span4Mux_v I__13768 (
            .O(N__55656),
            .I(N__55617));
    InMux I__13767 (
            .O(N__55655),
            .I(N__55614));
    LocalMux I__13766 (
            .O(N__55640),
            .I(N__55608));
    LocalMux I__13765 (
            .O(N__55635),
            .I(N__55608));
    InMux I__13764 (
            .O(N__55634),
            .I(N__55603));
    InMux I__13763 (
            .O(N__55633),
            .I(N__55603));
    InMux I__13762 (
            .O(N__55632),
            .I(N__55592));
    InMux I__13761 (
            .O(N__55631),
            .I(N__55592));
    InMux I__13760 (
            .O(N__55630),
            .I(N__55592));
    InMux I__13759 (
            .O(N__55629),
            .I(N__55592));
    InMux I__13758 (
            .O(N__55628),
            .I(N__55592));
    InMux I__13757 (
            .O(N__55627),
            .I(N__55589));
    InMux I__13756 (
            .O(N__55626),
            .I(N__55586));
    LocalMux I__13755 (
            .O(N__55623),
            .I(N__55582));
    InMux I__13754 (
            .O(N__55622),
            .I(N__55579));
    InMux I__13753 (
            .O(N__55621),
            .I(N__55574));
    InMux I__13752 (
            .O(N__55620),
            .I(N__55574));
    Span4Mux_h I__13751 (
            .O(N__55617),
            .I(N__55571));
    LocalMux I__13750 (
            .O(N__55614),
            .I(N__55568));
    InMux I__13749 (
            .O(N__55613),
            .I(N__55563));
    Span4Mux_h I__13748 (
            .O(N__55608),
            .I(N__55556));
    LocalMux I__13747 (
            .O(N__55603),
            .I(N__55556));
    LocalMux I__13746 (
            .O(N__55592),
            .I(N__55556));
    LocalMux I__13745 (
            .O(N__55589),
            .I(N__55553));
    LocalMux I__13744 (
            .O(N__55586),
            .I(N__55550));
    InMux I__13743 (
            .O(N__55585),
            .I(N__55547));
    Span4Mux_h I__13742 (
            .O(N__55582),
            .I(N__55540));
    LocalMux I__13741 (
            .O(N__55579),
            .I(N__55540));
    LocalMux I__13740 (
            .O(N__55574),
            .I(N__55540));
    Span4Mux_h I__13739 (
            .O(N__55571),
            .I(N__55537));
    Span12Mux_h I__13738 (
            .O(N__55568),
            .I(N__55534));
    InMux I__13737 (
            .O(N__55567),
            .I(N__55529));
    InMux I__13736 (
            .O(N__55566),
            .I(N__55529));
    LocalMux I__13735 (
            .O(N__55563),
            .I(N__55524));
    Span4Mux_h I__13734 (
            .O(N__55556),
            .I(N__55524));
    Span4Mux_v I__13733 (
            .O(N__55553),
            .I(N__55515));
    Span4Mux_h I__13732 (
            .O(N__55550),
            .I(N__55515));
    LocalMux I__13731 (
            .O(N__55547),
            .I(N__55515));
    Span4Mux_h I__13730 (
            .O(N__55540),
            .I(N__55515));
    Odrv4 I__13729 (
            .O(N__55537),
            .I(dds_state_1));
    Odrv12 I__13728 (
            .O(N__55534),
            .I(dds_state_1));
    LocalMux I__13727 (
            .O(N__55529),
            .I(dds_state_1));
    Odrv4 I__13726 (
            .O(N__55524),
            .I(dds_state_1));
    Odrv4 I__13725 (
            .O(N__55515),
            .I(dds_state_1));
    IoInMux I__13724 (
            .O(N__55504),
            .I(N__55501));
    LocalMux I__13723 (
            .O(N__55501),
            .I(N__55498));
    Span4Mux_s0_v I__13722 (
            .O(N__55498),
            .I(N__55495));
    Span4Mux_h I__13721 (
            .O(N__55495),
            .I(N__55492));
    Span4Mux_v I__13720 (
            .O(N__55492),
            .I(N__55489));
    Span4Mux_v I__13719 (
            .O(N__55489),
            .I(N__55486));
    Odrv4 I__13718 (
            .O(N__55486),
            .I(DDS_CS));
    CEMux I__13717 (
            .O(N__55483),
            .I(N__55480));
    LocalMux I__13716 (
            .O(N__55480),
            .I(N__55477));
    Odrv4 I__13715 (
            .O(N__55477),
            .I(\SIG_DDS.n9_adj_1385 ));
    InMux I__13714 (
            .O(N__55474),
            .I(N__55469));
    CascadeMux I__13713 (
            .O(N__55473),
            .I(N__55466));
    InMux I__13712 (
            .O(N__55472),
            .I(N__55455));
    LocalMux I__13711 (
            .O(N__55469),
            .I(N__55452));
    InMux I__13710 (
            .O(N__55466),
            .I(N__55443));
    InMux I__13709 (
            .O(N__55465),
            .I(N__55443));
    InMux I__13708 (
            .O(N__55464),
            .I(N__55443));
    InMux I__13707 (
            .O(N__55463),
            .I(N__55443));
    InMux I__13706 (
            .O(N__55462),
            .I(N__55438));
    InMux I__13705 (
            .O(N__55461),
            .I(N__55438));
    InMux I__13704 (
            .O(N__55460),
            .I(N__55432));
    InMux I__13703 (
            .O(N__55459),
            .I(N__55432));
    InMux I__13702 (
            .O(N__55458),
            .I(N__55418));
    LocalMux I__13701 (
            .O(N__55455),
            .I(N__55415));
    Span4Mux_v I__13700 (
            .O(N__55452),
            .I(N__55410));
    LocalMux I__13699 (
            .O(N__55443),
            .I(N__55410));
    LocalMux I__13698 (
            .O(N__55438),
            .I(N__55398));
    SRMux I__13697 (
            .O(N__55437),
            .I(N__55395));
    LocalMux I__13696 (
            .O(N__55432),
            .I(N__55392));
    SRMux I__13695 (
            .O(N__55431),
            .I(N__55389));
    InMux I__13694 (
            .O(N__55430),
            .I(N__55384));
    InMux I__13693 (
            .O(N__55429),
            .I(N__55384));
    InMux I__13692 (
            .O(N__55428),
            .I(N__55379));
    InMux I__13691 (
            .O(N__55427),
            .I(N__55362));
    InMux I__13690 (
            .O(N__55426),
            .I(N__55362));
    InMux I__13689 (
            .O(N__55425),
            .I(N__55362));
    InMux I__13688 (
            .O(N__55424),
            .I(N__55362));
    InMux I__13687 (
            .O(N__55423),
            .I(N__55362));
    InMux I__13686 (
            .O(N__55422),
            .I(N__55362));
    InMux I__13685 (
            .O(N__55421),
            .I(N__55362));
    LocalMux I__13684 (
            .O(N__55418),
            .I(N__55355));
    Span4Mux_h I__13683 (
            .O(N__55415),
            .I(N__55355));
    Span4Mux_h I__13682 (
            .O(N__55410),
            .I(N__55355));
    InMux I__13681 (
            .O(N__55409),
            .I(N__55350));
    InMux I__13680 (
            .O(N__55408),
            .I(N__55350));
    InMux I__13679 (
            .O(N__55407),
            .I(N__55347));
    InMux I__13678 (
            .O(N__55406),
            .I(N__55342));
    InMux I__13677 (
            .O(N__55405),
            .I(N__55342));
    InMux I__13676 (
            .O(N__55404),
            .I(N__55333));
    InMux I__13675 (
            .O(N__55403),
            .I(N__55333));
    InMux I__13674 (
            .O(N__55402),
            .I(N__55333));
    InMux I__13673 (
            .O(N__55401),
            .I(N__55333));
    Span4Mux_v I__13672 (
            .O(N__55398),
            .I(N__55328));
    LocalMux I__13671 (
            .O(N__55395),
            .I(N__55328));
    Span4Mux_v I__13670 (
            .O(N__55392),
            .I(N__55321));
    LocalMux I__13669 (
            .O(N__55389),
            .I(N__55321));
    LocalMux I__13668 (
            .O(N__55384),
            .I(N__55321));
    SRMux I__13667 (
            .O(N__55383),
            .I(N__55318));
    InMux I__13666 (
            .O(N__55382),
            .I(N__55315));
    LocalMux I__13665 (
            .O(N__55379),
            .I(N__55312));
    InMux I__13664 (
            .O(N__55378),
            .I(N__55307));
    InMux I__13663 (
            .O(N__55377),
            .I(N__55307));
    LocalMux I__13662 (
            .O(N__55362),
            .I(N__55304));
    Span4Mux_v I__13661 (
            .O(N__55355),
            .I(N__55299));
    LocalMux I__13660 (
            .O(N__55350),
            .I(N__55299));
    LocalMux I__13659 (
            .O(N__55347),
            .I(N__55294));
    LocalMux I__13658 (
            .O(N__55342),
            .I(N__55294));
    LocalMux I__13657 (
            .O(N__55333),
            .I(N__55291));
    Span4Mux_h I__13656 (
            .O(N__55328),
            .I(N__55284));
    Span4Mux_h I__13655 (
            .O(N__55321),
            .I(N__55284));
    LocalMux I__13654 (
            .O(N__55318),
            .I(N__55284));
    LocalMux I__13653 (
            .O(N__55315),
            .I(N__55281));
    Span4Mux_v I__13652 (
            .O(N__55312),
            .I(N__55274));
    LocalMux I__13651 (
            .O(N__55307),
            .I(N__55274));
    Span4Mux_h I__13650 (
            .O(N__55304),
            .I(N__55274));
    Span4Mux_h I__13649 (
            .O(N__55299),
            .I(N__55271));
    Span4Mux_h I__13648 (
            .O(N__55294),
            .I(N__55268));
    Span4Mux_v I__13647 (
            .O(N__55291),
            .I(N__55263));
    Span4Mux_h I__13646 (
            .O(N__55284),
            .I(N__55263));
    Span4Mux_h I__13645 (
            .O(N__55281),
            .I(N__55258));
    Span4Mux_h I__13644 (
            .O(N__55274),
            .I(N__55258));
    Span4Mux_h I__13643 (
            .O(N__55271),
            .I(N__55255));
    Odrv4 I__13642 (
            .O(N__55268),
            .I(comm_clear));
    Odrv4 I__13641 (
            .O(N__55263),
            .I(comm_clear));
    Odrv4 I__13640 (
            .O(N__55258),
            .I(comm_clear));
    Odrv4 I__13639 (
            .O(N__55255),
            .I(comm_clear));
    ClkMux I__13638 (
            .O(N__55246),
            .I(N__54727));
    ClkMux I__13637 (
            .O(N__55245),
            .I(N__54727));
    ClkMux I__13636 (
            .O(N__55244),
            .I(N__54727));
    ClkMux I__13635 (
            .O(N__55243),
            .I(N__54727));
    ClkMux I__13634 (
            .O(N__55242),
            .I(N__54727));
    ClkMux I__13633 (
            .O(N__55241),
            .I(N__54727));
    ClkMux I__13632 (
            .O(N__55240),
            .I(N__54727));
    ClkMux I__13631 (
            .O(N__55239),
            .I(N__54727));
    ClkMux I__13630 (
            .O(N__55238),
            .I(N__54727));
    ClkMux I__13629 (
            .O(N__55237),
            .I(N__54727));
    ClkMux I__13628 (
            .O(N__55236),
            .I(N__54727));
    ClkMux I__13627 (
            .O(N__55235),
            .I(N__54727));
    ClkMux I__13626 (
            .O(N__55234),
            .I(N__54727));
    ClkMux I__13625 (
            .O(N__55233),
            .I(N__54727));
    ClkMux I__13624 (
            .O(N__55232),
            .I(N__54727));
    ClkMux I__13623 (
            .O(N__55231),
            .I(N__54727));
    ClkMux I__13622 (
            .O(N__55230),
            .I(N__54727));
    ClkMux I__13621 (
            .O(N__55229),
            .I(N__54727));
    ClkMux I__13620 (
            .O(N__55228),
            .I(N__54727));
    ClkMux I__13619 (
            .O(N__55227),
            .I(N__54727));
    ClkMux I__13618 (
            .O(N__55226),
            .I(N__54727));
    ClkMux I__13617 (
            .O(N__55225),
            .I(N__54727));
    ClkMux I__13616 (
            .O(N__55224),
            .I(N__54727));
    ClkMux I__13615 (
            .O(N__55223),
            .I(N__54727));
    ClkMux I__13614 (
            .O(N__55222),
            .I(N__54727));
    ClkMux I__13613 (
            .O(N__55221),
            .I(N__54727));
    ClkMux I__13612 (
            .O(N__55220),
            .I(N__54727));
    ClkMux I__13611 (
            .O(N__55219),
            .I(N__54727));
    ClkMux I__13610 (
            .O(N__55218),
            .I(N__54727));
    ClkMux I__13609 (
            .O(N__55217),
            .I(N__54727));
    ClkMux I__13608 (
            .O(N__55216),
            .I(N__54727));
    ClkMux I__13607 (
            .O(N__55215),
            .I(N__54727));
    ClkMux I__13606 (
            .O(N__55214),
            .I(N__54727));
    ClkMux I__13605 (
            .O(N__55213),
            .I(N__54727));
    ClkMux I__13604 (
            .O(N__55212),
            .I(N__54727));
    ClkMux I__13603 (
            .O(N__55211),
            .I(N__54727));
    ClkMux I__13602 (
            .O(N__55210),
            .I(N__54727));
    ClkMux I__13601 (
            .O(N__55209),
            .I(N__54727));
    ClkMux I__13600 (
            .O(N__55208),
            .I(N__54727));
    ClkMux I__13599 (
            .O(N__55207),
            .I(N__54727));
    ClkMux I__13598 (
            .O(N__55206),
            .I(N__54727));
    ClkMux I__13597 (
            .O(N__55205),
            .I(N__54727));
    ClkMux I__13596 (
            .O(N__55204),
            .I(N__54727));
    ClkMux I__13595 (
            .O(N__55203),
            .I(N__54727));
    ClkMux I__13594 (
            .O(N__55202),
            .I(N__54727));
    ClkMux I__13593 (
            .O(N__55201),
            .I(N__54727));
    ClkMux I__13592 (
            .O(N__55200),
            .I(N__54727));
    ClkMux I__13591 (
            .O(N__55199),
            .I(N__54727));
    ClkMux I__13590 (
            .O(N__55198),
            .I(N__54727));
    ClkMux I__13589 (
            .O(N__55197),
            .I(N__54727));
    ClkMux I__13588 (
            .O(N__55196),
            .I(N__54727));
    ClkMux I__13587 (
            .O(N__55195),
            .I(N__54727));
    ClkMux I__13586 (
            .O(N__55194),
            .I(N__54727));
    ClkMux I__13585 (
            .O(N__55193),
            .I(N__54727));
    ClkMux I__13584 (
            .O(N__55192),
            .I(N__54727));
    ClkMux I__13583 (
            .O(N__55191),
            .I(N__54727));
    ClkMux I__13582 (
            .O(N__55190),
            .I(N__54727));
    ClkMux I__13581 (
            .O(N__55189),
            .I(N__54727));
    ClkMux I__13580 (
            .O(N__55188),
            .I(N__54727));
    ClkMux I__13579 (
            .O(N__55187),
            .I(N__54727));
    ClkMux I__13578 (
            .O(N__55186),
            .I(N__54727));
    ClkMux I__13577 (
            .O(N__55185),
            .I(N__54727));
    ClkMux I__13576 (
            .O(N__55184),
            .I(N__54727));
    ClkMux I__13575 (
            .O(N__55183),
            .I(N__54727));
    ClkMux I__13574 (
            .O(N__55182),
            .I(N__54727));
    ClkMux I__13573 (
            .O(N__55181),
            .I(N__54727));
    ClkMux I__13572 (
            .O(N__55180),
            .I(N__54727));
    ClkMux I__13571 (
            .O(N__55179),
            .I(N__54727));
    ClkMux I__13570 (
            .O(N__55178),
            .I(N__54727));
    ClkMux I__13569 (
            .O(N__55177),
            .I(N__54727));
    ClkMux I__13568 (
            .O(N__55176),
            .I(N__54727));
    ClkMux I__13567 (
            .O(N__55175),
            .I(N__54727));
    ClkMux I__13566 (
            .O(N__55174),
            .I(N__54727));
    ClkMux I__13565 (
            .O(N__55173),
            .I(N__54727));
    ClkMux I__13564 (
            .O(N__55172),
            .I(N__54727));
    ClkMux I__13563 (
            .O(N__55171),
            .I(N__54727));
    ClkMux I__13562 (
            .O(N__55170),
            .I(N__54727));
    ClkMux I__13561 (
            .O(N__55169),
            .I(N__54727));
    ClkMux I__13560 (
            .O(N__55168),
            .I(N__54727));
    ClkMux I__13559 (
            .O(N__55167),
            .I(N__54727));
    ClkMux I__13558 (
            .O(N__55166),
            .I(N__54727));
    ClkMux I__13557 (
            .O(N__55165),
            .I(N__54727));
    ClkMux I__13556 (
            .O(N__55164),
            .I(N__54727));
    ClkMux I__13555 (
            .O(N__55163),
            .I(N__54727));
    ClkMux I__13554 (
            .O(N__55162),
            .I(N__54727));
    ClkMux I__13553 (
            .O(N__55161),
            .I(N__54727));
    ClkMux I__13552 (
            .O(N__55160),
            .I(N__54727));
    ClkMux I__13551 (
            .O(N__55159),
            .I(N__54727));
    ClkMux I__13550 (
            .O(N__55158),
            .I(N__54727));
    ClkMux I__13549 (
            .O(N__55157),
            .I(N__54727));
    ClkMux I__13548 (
            .O(N__55156),
            .I(N__54727));
    ClkMux I__13547 (
            .O(N__55155),
            .I(N__54727));
    ClkMux I__13546 (
            .O(N__55154),
            .I(N__54727));
    ClkMux I__13545 (
            .O(N__55153),
            .I(N__54727));
    ClkMux I__13544 (
            .O(N__55152),
            .I(N__54727));
    ClkMux I__13543 (
            .O(N__55151),
            .I(N__54727));
    ClkMux I__13542 (
            .O(N__55150),
            .I(N__54727));
    ClkMux I__13541 (
            .O(N__55149),
            .I(N__54727));
    ClkMux I__13540 (
            .O(N__55148),
            .I(N__54727));
    ClkMux I__13539 (
            .O(N__55147),
            .I(N__54727));
    ClkMux I__13538 (
            .O(N__55146),
            .I(N__54727));
    ClkMux I__13537 (
            .O(N__55145),
            .I(N__54727));
    ClkMux I__13536 (
            .O(N__55144),
            .I(N__54727));
    ClkMux I__13535 (
            .O(N__55143),
            .I(N__54727));
    ClkMux I__13534 (
            .O(N__55142),
            .I(N__54727));
    ClkMux I__13533 (
            .O(N__55141),
            .I(N__54727));
    ClkMux I__13532 (
            .O(N__55140),
            .I(N__54727));
    ClkMux I__13531 (
            .O(N__55139),
            .I(N__54727));
    ClkMux I__13530 (
            .O(N__55138),
            .I(N__54727));
    ClkMux I__13529 (
            .O(N__55137),
            .I(N__54727));
    ClkMux I__13528 (
            .O(N__55136),
            .I(N__54727));
    ClkMux I__13527 (
            .O(N__55135),
            .I(N__54727));
    ClkMux I__13526 (
            .O(N__55134),
            .I(N__54727));
    ClkMux I__13525 (
            .O(N__55133),
            .I(N__54727));
    ClkMux I__13524 (
            .O(N__55132),
            .I(N__54727));
    ClkMux I__13523 (
            .O(N__55131),
            .I(N__54727));
    ClkMux I__13522 (
            .O(N__55130),
            .I(N__54727));
    ClkMux I__13521 (
            .O(N__55129),
            .I(N__54727));
    ClkMux I__13520 (
            .O(N__55128),
            .I(N__54727));
    ClkMux I__13519 (
            .O(N__55127),
            .I(N__54727));
    ClkMux I__13518 (
            .O(N__55126),
            .I(N__54727));
    ClkMux I__13517 (
            .O(N__55125),
            .I(N__54727));
    ClkMux I__13516 (
            .O(N__55124),
            .I(N__54727));
    ClkMux I__13515 (
            .O(N__55123),
            .I(N__54727));
    ClkMux I__13514 (
            .O(N__55122),
            .I(N__54727));
    ClkMux I__13513 (
            .O(N__55121),
            .I(N__54727));
    ClkMux I__13512 (
            .O(N__55120),
            .I(N__54727));
    ClkMux I__13511 (
            .O(N__55119),
            .I(N__54727));
    ClkMux I__13510 (
            .O(N__55118),
            .I(N__54727));
    ClkMux I__13509 (
            .O(N__55117),
            .I(N__54727));
    ClkMux I__13508 (
            .O(N__55116),
            .I(N__54727));
    ClkMux I__13507 (
            .O(N__55115),
            .I(N__54727));
    ClkMux I__13506 (
            .O(N__55114),
            .I(N__54727));
    ClkMux I__13505 (
            .O(N__55113),
            .I(N__54727));
    ClkMux I__13504 (
            .O(N__55112),
            .I(N__54727));
    ClkMux I__13503 (
            .O(N__55111),
            .I(N__54727));
    ClkMux I__13502 (
            .O(N__55110),
            .I(N__54727));
    ClkMux I__13501 (
            .O(N__55109),
            .I(N__54727));
    ClkMux I__13500 (
            .O(N__55108),
            .I(N__54727));
    ClkMux I__13499 (
            .O(N__55107),
            .I(N__54727));
    ClkMux I__13498 (
            .O(N__55106),
            .I(N__54727));
    ClkMux I__13497 (
            .O(N__55105),
            .I(N__54727));
    ClkMux I__13496 (
            .O(N__55104),
            .I(N__54727));
    ClkMux I__13495 (
            .O(N__55103),
            .I(N__54727));
    ClkMux I__13494 (
            .O(N__55102),
            .I(N__54727));
    ClkMux I__13493 (
            .O(N__55101),
            .I(N__54727));
    ClkMux I__13492 (
            .O(N__55100),
            .I(N__54727));
    ClkMux I__13491 (
            .O(N__55099),
            .I(N__54727));
    ClkMux I__13490 (
            .O(N__55098),
            .I(N__54727));
    ClkMux I__13489 (
            .O(N__55097),
            .I(N__54727));
    ClkMux I__13488 (
            .O(N__55096),
            .I(N__54727));
    ClkMux I__13487 (
            .O(N__55095),
            .I(N__54727));
    ClkMux I__13486 (
            .O(N__55094),
            .I(N__54727));
    ClkMux I__13485 (
            .O(N__55093),
            .I(N__54727));
    ClkMux I__13484 (
            .O(N__55092),
            .I(N__54727));
    ClkMux I__13483 (
            .O(N__55091),
            .I(N__54727));
    ClkMux I__13482 (
            .O(N__55090),
            .I(N__54727));
    ClkMux I__13481 (
            .O(N__55089),
            .I(N__54727));
    ClkMux I__13480 (
            .O(N__55088),
            .I(N__54727));
    ClkMux I__13479 (
            .O(N__55087),
            .I(N__54727));
    ClkMux I__13478 (
            .O(N__55086),
            .I(N__54727));
    ClkMux I__13477 (
            .O(N__55085),
            .I(N__54727));
    ClkMux I__13476 (
            .O(N__55084),
            .I(N__54727));
    ClkMux I__13475 (
            .O(N__55083),
            .I(N__54727));
    ClkMux I__13474 (
            .O(N__55082),
            .I(N__54727));
    ClkMux I__13473 (
            .O(N__55081),
            .I(N__54727));
    ClkMux I__13472 (
            .O(N__55080),
            .I(N__54727));
    ClkMux I__13471 (
            .O(N__55079),
            .I(N__54727));
    ClkMux I__13470 (
            .O(N__55078),
            .I(N__54727));
    ClkMux I__13469 (
            .O(N__55077),
            .I(N__54727));
    ClkMux I__13468 (
            .O(N__55076),
            .I(N__54727));
    ClkMux I__13467 (
            .O(N__55075),
            .I(N__54727));
    ClkMux I__13466 (
            .O(N__55074),
            .I(N__54727));
    GlobalMux I__13465 (
            .O(N__54727),
            .I(clk_32MHz));
    InMux I__13464 (
            .O(N__54724),
            .I(N__54706));
    InMux I__13463 (
            .O(N__54723),
            .I(N__54696));
    InMux I__13462 (
            .O(N__54722),
            .I(N__54690));
    InMux I__13461 (
            .O(N__54721),
            .I(N__54687));
    InMux I__13460 (
            .O(N__54720),
            .I(N__54684));
    InMux I__13459 (
            .O(N__54719),
            .I(N__54681));
    InMux I__13458 (
            .O(N__54718),
            .I(N__54676));
    InMux I__13457 (
            .O(N__54717),
            .I(N__54676));
    CascadeMux I__13456 (
            .O(N__54716),
            .I(N__54653));
    CascadeMux I__13455 (
            .O(N__54715),
            .I(N__54650));
    CascadeMux I__13454 (
            .O(N__54714),
            .I(N__54646));
    CascadeMux I__13453 (
            .O(N__54713),
            .I(N__54642));
    CascadeMux I__13452 (
            .O(N__54712),
            .I(N__54639));
    CascadeMux I__13451 (
            .O(N__54711),
            .I(N__54636));
    InMux I__13450 (
            .O(N__54710),
            .I(N__54632));
    InMux I__13449 (
            .O(N__54709),
            .I(N__54629));
    LocalMux I__13448 (
            .O(N__54706),
            .I(N__54626));
    InMux I__13447 (
            .O(N__54705),
            .I(N__54620));
    InMux I__13446 (
            .O(N__54704),
            .I(N__54617));
    InMux I__13445 (
            .O(N__54703),
            .I(N__54612));
    InMux I__13444 (
            .O(N__54702),
            .I(N__54612));
    InMux I__13443 (
            .O(N__54701),
            .I(N__54604));
    InMux I__13442 (
            .O(N__54700),
            .I(N__54604));
    InMux I__13441 (
            .O(N__54699),
            .I(N__54601));
    LocalMux I__13440 (
            .O(N__54696),
            .I(N__54593));
    CascadeMux I__13439 (
            .O(N__54695),
            .I(N__54585));
    CascadeMux I__13438 (
            .O(N__54694),
            .I(N__54581));
    CascadeMux I__13437 (
            .O(N__54693),
            .I(N__54577));
    LocalMux I__13436 (
            .O(N__54690),
            .I(N__54571));
    LocalMux I__13435 (
            .O(N__54687),
            .I(N__54571));
    LocalMux I__13434 (
            .O(N__54684),
            .I(N__54564));
    LocalMux I__13433 (
            .O(N__54681),
            .I(N__54564));
    LocalMux I__13432 (
            .O(N__54676),
            .I(N__54564));
    InMux I__13431 (
            .O(N__54675),
            .I(N__54558));
    InMux I__13430 (
            .O(N__54674),
            .I(N__54555));
    InMux I__13429 (
            .O(N__54673),
            .I(N__54550));
    InMux I__13428 (
            .O(N__54672),
            .I(N__54550));
    InMux I__13427 (
            .O(N__54671),
            .I(N__54545));
    InMux I__13426 (
            .O(N__54670),
            .I(N__54545));
    CascadeMux I__13425 (
            .O(N__54669),
            .I(N__54541));
    InMux I__13424 (
            .O(N__54668),
            .I(N__54538));
    InMux I__13423 (
            .O(N__54667),
            .I(N__54522));
    InMux I__13422 (
            .O(N__54666),
            .I(N__54522));
    InMux I__13421 (
            .O(N__54665),
            .I(N__54522));
    InMux I__13420 (
            .O(N__54664),
            .I(N__54522));
    InMux I__13419 (
            .O(N__54663),
            .I(N__54522));
    InMux I__13418 (
            .O(N__54662),
            .I(N__54522));
    InMux I__13417 (
            .O(N__54661),
            .I(N__54511));
    InMux I__13416 (
            .O(N__54660),
            .I(N__54511));
    InMux I__13415 (
            .O(N__54659),
            .I(N__54511));
    InMux I__13414 (
            .O(N__54658),
            .I(N__54511));
    InMux I__13413 (
            .O(N__54657),
            .I(N__54511));
    InMux I__13412 (
            .O(N__54656),
            .I(N__54508));
    InMux I__13411 (
            .O(N__54653),
            .I(N__54495));
    InMux I__13410 (
            .O(N__54650),
            .I(N__54495));
    InMux I__13409 (
            .O(N__54649),
            .I(N__54495));
    InMux I__13408 (
            .O(N__54646),
            .I(N__54495));
    InMux I__13407 (
            .O(N__54645),
            .I(N__54495));
    InMux I__13406 (
            .O(N__54642),
            .I(N__54495));
    InMux I__13405 (
            .O(N__54639),
            .I(N__54490));
    InMux I__13404 (
            .O(N__54636),
            .I(N__54490));
    InMux I__13403 (
            .O(N__54635),
            .I(N__54482));
    LocalMux I__13402 (
            .O(N__54632),
            .I(N__54475));
    LocalMux I__13401 (
            .O(N__54629),
            .I(N__54475));
    Span4Mux_h I__13400 (
            .O(N__54626),
            .I(N__54475));
    InMux I__13399 (
            .O(N__54625),
            .I(N__54472));
    InMux I__13398 (
            .O(N__54624),
            .I(N__54467));
    InMux I__13397 (
            .O(N__54623),
            .I(N__54467));
    LocalMux I__13396 (
            .O(N__54620),
            .I(N__54460));
    LocalMux I__13395 (
            .O(N__54617),
            .I(N__54460));
    LocalMux I__13394 (
            .O(N__54612),
            .I(N__54460));
    InMux I__13393 (
            .O(N__54611),
            .I(N__54455));
    InMux I__13392 (
            .O(N__54610),
            .I(N__54455));
    SRMux I__13391 (
            .O(N__54609),
            .I(N__54452));
    LocalMux I__13390 (
            .O(N__54604),
            .I(N__54448));
    LocalMux I__13389 (
            .O(N__54601),
            .I(N__54445));
    InMux I__13388 (
            .O(N__54600),
            .I(N__54442));
    CascadeMux I__13387 (
            .O(N__54599),
            .I(N__54437));
    CascadeMux I__13386 (
            .O(N__54598),
            .I(N__54434));
    InMux I__13385 (
            .O(N__54597),
            .I(N__54430));
    InMux I__13384 (
            .O(N__54596),
            .I(N__54427));
    Span4Mux_h I__13383 (
            .O(N__54593),
            .I(N__54424));
    InMux I__13382 (
            .O(N__54592),
            .I(N__54421));
    InMux I__13381 (
            .O(N__54591),
            .I(N__54416));
    InMux I__13380 (
            .O(N__54590),
            .I(N__54416));
    InMux I__13379 (
            .O(N__54589),
            .I(N__54399));
    InMux I__13378 (
            .O(N__54588),
            .I(N__54399));
    InMux I__13377 (
            .O(N__54585),
            .I(N__54399));
    InMux I__13376 (
            .O(N__54584),
            .I(N__54399));
    InMux I__13375 (
            .O(N__54581),
            .I(N__54399));
    InMux I__13374 (
            .O(N__54580),
            .I(N__54399));
    InMux I__13373 (
            .O(N__54577),
            .I(N__54399));
    InMux I__13372 (
            .O(N__54576),
            .I(N__54399));
    Span4Mux_v I__13371 (
            .O(N__54571),
            .I(N__54394));
    Span4Mux_v I__13370 (
            .O(N__54564),
            .I(N__54394));
    InMux I__13369 (
            .O(N__54563),
            .I(N__54389));
    InMux I__13368 (
            .O(N__54562),
            .I(N__54389));
    InMux I__13367 (
            .O(N__54561),
            .I(N__54384));
    LocalMux I__13366 (
            .O(N__54558),
            .I(N__54381));
    LocalMux I__13365 (
            .O(N__54555),
            .I(N__54376));
    LocalMux I__13364 (
            .O(N__54550),
            .I(N__54376));
    LocalMux I__13363 (
            .O(N__54545),
            .I(N__54373));
    InMux I__13362 (
            .O(N__54544),
            .I(N__54369));
    InMux I__13361 (
            .O(N__54541),
            .I(N__54364));
    LocalMux I__13360 (
            .O(N__54538),
            .I(N__54361));
    InMux I__13359 (
            .O(N__54537),
            .I(N__54358));
    InMux I__13358 (
            .O(N__54536),
            .I(N__54355));
    InMux I__13357 (
            .O(N__54535),
            .I(N__54352));
    LocalMux I__13356 (
            .O(N__54522),
            .I(N__54341));
    LocalMux I__13355 (
            .O(N__54511),
            .I(N__54341));
    LocalMux I__13354 (
            .O(N__54508),
            .I(N__54341));
    LocalMux I__13353 (
            .O(N__54495),
            .I(N__54341));
    LocalMux I__13352 (
            .O(N__54490),
            .I(N__54341));
    InMux I__13351 (
            .O(N__54489),
            .I(N__54336));
    InMux I__13350 (
            .O(N__54488),
            .I(N__54336));
    InMux I__13349 (
            .O(N__54487),
            .I(N__54329));
    InMux I__13348 (
            .O(N__54486),
            .I(N__54329));
    InMux I__13347 (
            .O(N__54485),
            .I(N__54329));
    LocalMux I__13346 (
            .O(N__54482),
            .I(N__54318));
    Span4Mux_h I__13345 (
            .O(N__54475),
            .I(N__54318));
    LocalMux I__13344 (
            .O(N__54472),
            .I(N__54318));
    LocalMux I__13343 (
            .O(N__54467),
            .I(N__54318));
    Span4Mux_v I__13342 (
            .O(N__54460),
            .I(N__54318));
    LocalMux I__13341 (
            .O(N__54455),
            .I(N__54315));
    LocalMux I__13340 (
            .O(N__54452),
            .I(N__54312));
    InMux I__13339 (
            .O(N__54451),
            .I(N__54309));
    Span4Mux_h I__13338 (
            .O(N__54448),
            .I(N__54306));
    Span4Mux_h I__13337 (
            .O(N__54445),
            .I(N__54301));
    LocalMux I__13336 (
            .O(N__54442),
            .I(N__54301));
    InMux I__13335 (
            .O(N__54441),
            .I(N__54298));
    InMux I__13334 (
            .O(N__54440),
            .I(N__54295));
    InMux I__13333 (
            .O(N__54437),
            .I(N__54288));
    InMux I__13332 (
            .O(N__54434),
            .I(N__54288));
    InMux I__13331 (
            .O(N__54433),
            .I(N__54288));
    LocalMux I__13330 (
            .O(N__54430),
            .I(N__54285));
    LocalMux I__13329 (
            .O(N__54427),
            .I(N__54280));
    Span4Mux_h I__13328 (
            .O(N__54424),
            .I(N__54280));
    LocalMux I__13327 (
            .O(N__54421),
            .I(N__54275));
    LocalMux I__13326 (
            .O(N__54416),
            .I(N__54275));
    LocalMux I__13325 (
            .O(N__54399),
            .I(N__54268));
    Span4Mux_h I__13324 (
            .O(N__54394),
            .I(N__54268));
    LocalMux I__13323 (
            .O(N__54389),
            .I(N__54268));
    InMux I__13322 (
            .O(N__54388),
            .I(N__54263));
    InMux I__13321 (
            .O(N__54387),
            .I(N__54263));
    LocalMux I__13320 (
            .O(N__54384),
            .I(N__54260));
    Span4Mux_v I__13319 (
            .O(N__54381),
            .I(N__54253));
    Span4Mux_h I__13318 (
            .O(N__54376),
            .I(N__54253));
    Span4Mux_v I__13317 (
            .O(N__54373),
            .I(N__54253));
    InMux I__13316 (
            .O(N__54372),
            .I(N__54250));
    LocalMux I__13315 (
            .O(N__54369),
            .I(N__54246));
    CascadeMux I__13314 (
            .O(N__54368),
            .I(N__54241));
    InMux I__13313 (
            .O(N__54367),
            .I(N__54235));
    LocalMux I__13312 (
            .O(N__54364),
            .I(N__54228));
    Span4Mux_v I__13311 (
            .O(N__54361),
            .I(N__54228));
    LocalMux I__13310 (
            .O(N__54358),
            .I(N__54228));
    LocalMux I__13309 (
            .O(N__54355),
            .I(N__54223));
    LocalMux I__13308 (
            .O(N__54352),
            .I(N__54223));
    Span4Mux_v I__13307 (
            .O(N__54341),
            .I(N__54220));
    LocalMux I__13306 (
            .O(N__54336),
            .I(N__54211));
    LocalMux I__13305 (
            .O(N__54329),
            .I(N__54211));
    Span4Mux_v I__13304 (
            .O(N__54318),
            .I(N__54211));
    Span4Mux_v I__13303 (
            .O(N__54315),
            .I(N__54211));
    Span4Mux_v I__13302 (
            .O(N__54312),
            .I(N__54200));
    LocalMux I__13301 (
            .O(N__54309),
            .I(N__54200));
    Span4Mux_h I__13300 (
            .O(N__54306),
            .I(N__54200));
    Span4Mux_h I__13299 (
            .O(N__54301),
            .I(N__54200));
    LocalMux I__13298 (
            .O(N__54298),
            .I(N__54200));
    LocalMux I__13297 (
            .O(N__54295),
            .I(N__54193));
    LocalMux I__13296 (
            .O(N__54288),
            .I(N__54193));
    Span4Mux_h I__13295 (
            .O(N__54285),
            .I(N__54193));
    Sp12to4 I__13294 (
            .O(N__54280),
            .I(N__54184));
    Sp12to4 I__13293 (
            .O(N__54275),
            .I(N__54184));
    Sp12to4 I__13292 (
            .O(N__54268),
            .I(N__54184));
    LocalMux I__13291 (
            .O(N__54263),
            .I(N__54184));
    Span4Mux_h I__13290 (
            .O(N__54260),
            .I(N__54177));
    Span4Mux_v I__13289 (
            .O(N__54253),
            .I(N__54177));
    LocalMux I__13288 (
            .O(N__54250),
            .I(N__54177));
    InMux I__13287 (
            .O(N__54249),
            .I(N__54172));
    Span4Mux_h I__13286 (
            .O(N__54246),
            .I(N__54169));
    InMux I__13285 (
            .O(N__54245),
            .I(N__54166));
    InMux I__13284 (
            .O(N__54244),
            .I(N__54157));
    InMux I__13283 (
            .O(N__54241),
            .I(N__54157));
    InMux I__13282 (
            .O(N__54240),
            .I(N__54157));
    InMux I__13281 (
            .O(N__54239),
            .I(N__54157));
    InMux I__13280 (
            .O(N__54238),
            .I(N__54154));
    LocalMux I__13279 (
            .O(N__54235),
            .I(N__54143));
    Span4Mux_v I__13278 (
            .O(N__54228),
            .I(N__54143));
    Span4Mux_v I__13277 (
            .O(N__54223),
            .I(N__54143));
    Span4Mux_h I__13276 (
            .O(N__54220),
            .I(N__54143));
    Span4Mux_v I__13275 (
            .O(N__54211),
            .I(N__54143));
    Sp12to4 I__13274 (
            .O(N__54200),
            .I(N__54138));
    Sp12to4 I__13273 (
            .O(N__54193),
            .I(N__54138));
    Span12Mux_v I__13272 (
            .O(N__54184),
            .I(N__54135));
    Span4Mux_h I__13271 (
            .O(N__54177),
            .I(N__54132));
    InMux I__13270 (
            .O(N__54176),
            .I(N__54127));
    InMux I__13269 (
            .O(N__54175),
            .I(N__54127));
    LocalMux I__13268 (
            .O(N__54172),
            .I(comm_state_3));
    Odrv4 I__13267 (
            .O(N__54169),
            .I(comm_state_3));
    LocalMux I__13266 (
            .O(N__54166),
            .I(comm_state_3));
    LocalMux I__13265 (
            .O(N__54157),
            .I(comm_state_3));
    LocalMux I__13264 (
            .O(N__54154),
            .I(comm_state_3));
    Odrv4 I__13263 (
            .O(N__54143),
            .I(comm_state_3));
    Odrv12 I__13262 (
            .O(N__54138),
            .I(comm_state_3));
    Odrv12 I__13261 (
            .O(N__54135),
            .I(comm_state_3));
    Odrv4 I__13260 (
            .O(N__54132),
            .I(comm_state_3));
    LocalMux I__13259 (
            .O(N__54127),
            .I(comm_state_3));
    InMux I__13258 (
            .O(N__54106),
            .I(N__54076));
    InMux I__13257 (
            .O(N__54105),
            .I(N__54067));
    InMux I__13256 (
            .O(N__54104),
            .I(N__54067));
    InMux I__13255 (
            .O(N__54103),
            .I(N__54067));
    InMux I__13254 (
            .O(N__54102),
            .I(N__54067));
    InMux I__13253 (
            .O(N__54101),
            .I(N__54064));
    InMux I__13252 (
            .O(N__54100),
            .I(N__54061));
    InMux I__13251 (
            .O(N__54099),
            .I(N__54052));
    InMux I__13250 (
            .O(N__54098),
            .I(N__54052));
    InMux I__13249 (
            .O(N__54097),
            .I(N__54052));
    InMux I__13248 (
            .O(N__54096),
            .I(N__54052));
    InMux I__13247 (
            .O(N__54095),
            .I(N__54048));
    InMux I__13246 (
            .O(N__54094),
            .I(N__54045));
    InMux I__13245 (
            .O(N__54093),
            .I(N__54042));
    InMux I__13244 (
            .O(N__54092),
            .I(N__54039));
    InMux I__13243 (
            .O(N__54091),
            .I(N__54036));
    InMux I__13242 (
            .O(N__54090),
            .I(N__54028));
    InMux I__13241 (
            .O(N__54089),
            .I(N__54010));
    InMux I__13240 (
            .O(N__54088),
            .I(N__54010));
    InMux I__13239 (
            .O(N__54087),
            .I(N__54010));
    InMux I__13238 (
            .O(N__54086),
            .I(N__54010));
    InMux I__13237 (
            .O(N__54085),
            .I(N__54010));
    InMux I__13236 (
            .O(N__54084),
            .I(N__54010));
    InMux I__13235 (
            .O(N__54083),
            .I(N__54010));
    InMux I__13234 (
            .O(N__54082),
            .I(N__54010));
    InMux I__13233 (
            .O(N__54081),
            .I(N__54005));
    InMux I__13232 (
            .O(N__54080),
            .I(N__54005));
    InMux I__13231 (
            .O(N__54079),
            .I(N__54002));
    LocalMux I__13230 (
            .O(N__54076),
            .I(N__53997));
    LocalMux I__13229 (
            .O(N__54067),
            .I(N__53988));
    LocalMux I__13228 (
            .O(N__54064),
            .I(N__53988));
    LocalMux I__13227 (
            .O(N__54061),
            .I(N__53988));
    LocalMux I__13226 (
            .O(N__54052),
            .I(N__53988));
    InMux I__13225 (
            .O(N__54051),
            .I(N__53972));
    LocalMux I__13224 (
            .O(N__54048),
            .I(N__53967));
    LocalMux I__13223 (
            .O(N__54045),
            .I(N__53967));
    LocalMux I__13222 (
            .O(N__54042),
            .I(N__53964));
    LocalMux I__13221 (
            .O(N__54039),
            .I(N__53961));
    LocalMux I__13220 (
            .O(N__54036),
            .I(N__53958));
    InMux I__13219 (
            .O(N__54035),
            .I(N__53953));
    InMux I__13218 (
            .O(N__54034),
            .I(N__53950));
    InMux I__13217 (
            .O(N__54033),
            .I(N__53932));
    InMux I__13216 (
            .O(N__54032),
            .I(N__53929));
    InMux I__13215 (
            .O(N__54031),
            .I(N__53926));
    LocalMux I__13214 (
            .O(N__54028),
            .I(N__53923));
    InMux I__13213 (
            .O(N__54027),
            .I(N__53920));
    LocalMux I__13212 (
            .O(N__54010),
            .I(N__53913));
    LocalMux I__13211 (
            .O(N__54005),
            .I(N__53913));
    LocalMux I__13210 (
            .O(N__54002),
            .I(N__53913));
    CascadeMux I__13209 (
            .O(N__54001),
            .I(N__53910));
    InMux I__13208 (
            .O(N__54000),
            .I(N__53905));
    Span4Mux_v I__13207 (
            .O(N__53997),
            .I(N__53895));
    Span4Mux_v I__13206 (
            .O(N__53988),
            .I(N__53895));
    InMux I__13205 (
            .O(N__53987),
            .I(N__53892));
    InMux I__13204 (
            .O(N__53986),
            .I(N__53889));
    InMux I__13203 (
            .O(N__53985),
            .I(N__53886));
    InMux I__13202 (
            .O(N__53984),
            .I(N__53878));
    InMux I__13201 (
            .O(N__53983),
            .I(N__53875));
    InMux I__13200 (
            .O(N__53982),
            .I(N__53854));
    InMux I__13199 (
            .O(N__53981),
            .I(N__53854));
    InMux I__13198 (
            .O(N__53980),
            .I(N__53854));
    InMux I__13197 (
            .O(N__53979),
            .I(N__53854));
    InMux I__13196 (
            .O(N__53978),
            .I(N__53854));
    InMux I__13195 (
            .O(N__53977),
            .I(N__53854));
    InMux I__13194 (
            .O(N__53976),
            .I(N__53854));
    InMux I__13193 (
            .O(N__53975),
            .I(N__53854));
    LocalMux I__13192 (
            .O(N__53972),
            .I(N__53851));
    Span4Mux_v I__13191 (
            .O(N__53967),
            .I(N__53848));
    Span4Mux_v I__13190 (
            .O(N__53964),
            .I(N__53843));
    Span4Mux_v I__13189 (
            .O(N__53961),
            .I(N__53843));
    Span4Mux_v I__13188 (
            .O(N__53958),
            .I(N__53840));
    InMux I__13187 (
            .O(N__53957),
            .I(N__53834));
    InMux I__13186 (
            .O(N__53956),
            .I(N__53831));
    LocalMux I__13185 (
            .O(N__53953),
            .I(N__53823));
    LocalMux I__13184 (
            .O(N__53950),
            .I(N__53823));
    InMux I__13183 (
            .O(N__53949),
            .I(N__53806));
    InMux I__13182 (
            .O(N__53948),
            .I(N__53806));
    InMux I__13181 (
            .O(N__53947),
            .I(N__53806));
    InMux I__13180 (
            .O(N__53946),
            .I(N__53806));
    InMux I__13179 (
            .O(N__53945),
            .I(N__53806));
    InMux I__13178 (
            .O(N__53944),
            .I(N__53806));
    InMux I__13177 (
            .O(N__53943),
            .I(N__53806));
    InMux I__13176 (
            .O(N__53942),
            .I(N__53806));
    InMux I__13175 (
            .O(N__53941),
            .I(N__53791));
    InMux I__13174 (
            .O(N__53940),
            .I(N__53791));
    InMux I__13173 (
            .O(N__53939),
            .I(N__53791));
    InMux I__13172 (
            .O(N__53938),
            .I(N__53791));
    InMux I__13171 (
            .O(N__53937),
            .I(N__53791));
    InMux I__13170 (
            .O(N__53936),
            .I(N__53791));
    InMux I__13169 (
            .O(N__53935),
            .I(N__53791));
    LocalMux I__13168 (
            .O(N__53932),
            .I(N__53780));
    LocalMux I__13167 (
            .O(N__53929),
            .I(N__53780));
    LocalMux I__13166 (
            .O(N__53926),
            .I(N__53780));
    Span4Mux_v I__13165 (
            .O(N__53923),
            .I(N__53780));
    LocalMux I__13164 (
            .O(N__53920),
            .I(N__53780));
    Span4Mux_v I__13163 (
            .O(N__53913),
            .I(N__53777));
    InMux I__13162 (
            .O(N__53910),
            .I(N__53774));
    InMux I__13161 (
            .O(N__53909),
            .I(N__53771));
    InMux I__13160 (
            .O(N__53908),
            .I(N__53768));
    LocalMux I__13159 (
            .O(N__53905),
            .I(N__53765));
    InMux I__13158 (
            .O(N__53904),
            .I(N__53756));
    InMux I__13157 (
            .O(N__53903),
            .I(N__53756));
    InMux I__13156 (
            .O(N__53902),
            .I(N__53756));
    InMux I__13155 (
            .O(N__53901),
            .I(N__53756));
    InMux I__13154 (
            .O(N__53900),
            .I(N__53753));
    Span4Mux_h I__13153 (
            .O(N__53895),
            .I(N__53750));
    LocalMux I__13152 (
            .O(N__53892),
            .I(N__53743));
    LocalMux I__13151 (
            .O(N__53889),
            .I(N__53743));
    LocalMux I__13150 (
            .O(N__53886),
            .I(N__53743));
    InMux I__13149 (
            .O(N__53885),
            .I(N__53733));
    InMux I__13148 (
            .O(N__53884),
            .I(N__53733));
    InMux I__13147 (
            .O(N__53883),
            .I(N__53733));
    InMux I__13146 (
            .O(N__53882),
            .I(N__53728));
    InMux I__13145 (
            .O(N__53881),
            .I(N__53728));
    LocalMux I__13144 (
            .O(N__53878),
            .I(N__53723));
    LocalMux I__13143 (
            .O(N__53875),
            .I(N__53723));
    InMux I__13142 (
            .O(N__53874),
            .I(N__53720));
    InMux I__13141 (
            .O(N__53873),
            .I(N__53713));
    InMux I__13140 (
            .O(N__53872),
            .I(N__53713));
    InMux I__13139 (
            .O(N__53871),
            .I(N__53713));
    LocalMux I__13138 (
            .O(N__53854),
            .I(N__53704));
    Span4Mux_v I__13137 (
            .O(N__53851),
            .I(N__53704));
    Span4Mux_h I__13136 (
            .O(N__53848),
            .I(N__53704));
    Span4Mux_h I__13135 (
            .O(N__53843),
            .I(N__53704));
    Span4Mux_h I__13134 (
            .O(N__53840),
            .I(N__53701));
    InMux I__13133 (
            .O(N__53839),
            .I(N__53696));
    InMux I__13132 (
            .O(N__53838),
            .I(N__53696));
    InMux I__13131 (
            .O(N__53837),
            .I(N__53693));
    LocalMux I__13130 (
            .O(N__53834),
            .I(N__53688));
    LocalMux I__13129 (
            .O(N__53831),
            .I(N__53688));
    CascadeMux I__13128 (
            .O(N__53830),
            .I(N__53682));
    InMux I__13127 (
            .O(N__53829),
            .I(N__53676));
    InMux I__13126 (
            .O(N__53828),
            .I(N__53673));
    Span4Mux_v I__13125 (
            .O(N__53823),
            .I(N__53670));
    LocalMux I__13124 (
            .O(N__53806),
            .I(N__53659));
    LocalMux I__13123 (
            .O(N__53791),
            .I(N__53659));
    Span4Mux_v I__13122 (
            .O(N__53780),
            .I(N__53659));
    Span4Mux_h I__13121 (
            .O(N__53777),
            .I(N__53659));
    LocalMux I__13120 (
            .O(N__53774),
            .I(N__53659));
    LocalMux I__13119 (
            .O(N__53771),
            .I(N__53645));
    LocalMux I__13118 (
            .O(N__53768),
            .I(N__53645));
    Sp12to4 I__13117 (
            .O(N__53765),
            .I(N__53645));
    LocalMux I__13116 (
            .O(N__53756),
            .I(N__53645));
    LocalMux I__13115 (
            .O(N__53753),
            .I(N__53638));
    Span4Mux_h I__13114 (
            .O(N__53750),
            .I(N__53638));
    Span4Mux_v I__13113 (
            .O(N__53743),
            .I(N__53638));
    InMux I__13112 (
            .O(N__53742),
            .I(N__53630));
    InMux I__13111 (
            .O(N__53741),
            .I(N__53630));
    InMux I__13110 (
            .O(N__53740),
            .I(N__53630));
    LocalMux I__13109 (
            .O(N__53733),
            .I(N__53623));
    LocalMux I__13108 (
            .O(N__53728),
            .I(N__53623));
    Span4Mux_v I__13107 (
            .O(N__53723),
            .I(N__53623));
    LocalMux I__13106 (
            .O(N__53720),
            .I(N__53608));
    LocalMux I__13105 (
            .O(N__53713),
            .I(N__53608));
    Span4Mux_h I__13104 (
            .O(N__53704),
            .I(N__53608));
    Span4Mux_h I__13103 (
            .O(N__53701),
            .I(N__53608));
    LocalMux I__13102 (
            .O(N__53696),
            .I(N__53608));
    LocalMux I__13101 (
            .O(N__53693),
            .I(N__53608));
    Span4Mux_v I__13100 (
            .O(N__53688),
            .I(N__53608));
    InMux I__13099 (
            .O(N__53687),
            .I(N__53601));
    InMux I__13098 (
            .O(N__53686),
            .I(N__53601));
    InMux I__13097 (
            .O(N__53685),
            .I(N__53601));
    InMux I__13096 (
            .O(N__53682),
            .I(N__53592));
    InMux I__13095 (
            .O(N__53681),
            .I(N__53592));
    InMux I__13094 (
            .O(N__53680),
            .I(N__53592));
    InMux I__13093 (
            .O(N__53679),
            .I(N__53592));
    LocalMux I__13092 (
            .O(N__53676),
            .I(N__53587));
    LocalMux I__13091 (
            .O(N__53673),
            .I(N__53587));
    Span4Mux_h I__13090 (
            .O(N__53670),
            .I(N__53582));
    Span4Mux_v I__13089 (
            .O(N__53659),
            .I(N__53582));
    InMux I__13088 (
            .O(N__53658),
            .I(N__53571));
    InMux I__13087 (
            .O(N__53657),
            .I(N__53571));
    InMux I__13086 (
            .O(N__53656),
            .I(N__53571));
    InMux I__13085 (
            .O(N__53655),
            .I(N__53571));
    InMux I__13084 (
            .O(N__53654),
            .I(N__53571));
    Span12Mux_v I__13083 (
            .O(N__53645),
            .I(N__53568));
    Span4Mux_v I__13082 (
            .O(N__53638),
            .I(N__53565));
    InMux I__13081 (
            .O(N__53637),
            .I(N__53562));
    LocalMux I__13080 (
            .O(N__53630),
            .I(N__53555));
    Span4Mux_v I__13079 (
            .O(N__53623),
            .I(N__53555));
    Span4Mux_v I__13078 (
            .O(N__53608),
            .I(N__53555));
    LocalMux I__13077 (
            .O(N__53601),
            .I(comm_state_1));
    LocalMux I__13076 (
            .O(N__53592),
            .I(comm_state_1));
    Odrv12 I__13075 (
            .O(N__53587),
            .I(comm_state_1));
    Odrv4 I__13074 (
            .O(N__53582),
            .I(comm_state_1));
    LocalMux I__13073 (
            .O(N__53571),
            .I(comm_state_1));
    Odrv12 I__13072 (
            .O(N__53568),
            .I(comm_state_1));
    Odrv4 I__13071 (
            .O(N__53565),
            .I(comm_state_1));
    LocalMux I__13070 (
            .O(N__53562),
            .I(comm_state_1));
    Odrv4 I__13069 (
            .O(N__53555),
            .I(comm_state_1));
    InMux I__13068 (
            .O(N__53536),
            .I(N__53533));
    LocalMux I__13067 (
            .O(N__53533),
            .I(N__53526));
    CascadeMux I__13066 (
            .O(N__53532),
            .I(N__53523));
    CascadeMux I__13065 (
            .O(N__53531),
            .I(N__53518));
    InMux I__13064 (
            .O(N__53530),
            .I(N__53513));
    InMux I__13063 (
            .O(N__53529),
            .I(N__53513));
    Span4Mux_h I__13062 (
            .O(N__53526),
            .I(N__53506));
    InMux I__13061 (
            .O(N__53523),
            .I(N__53503));
    InMux I__13060 (
            .O(N__53522),
            .I(N__53500));
    CascadeMux I__13059 (
            .O(N__53521),
            .I(N__53482));
    InMux I__13058 (
            .O(N__53518),
            .I(N__53479));
    LocalMux I__13057 (
            .O(N__53513),
            .I(N__53476));
    InMux I__13056 (
            .O(N__53512),
            .I(N__53467));
    InMux I__13055 (
            .O(N__53511),
            .I(N__53467));
    InMux I__13054 (
            .O(N__53510),
            .I(N__53467));
    InMux I__13053 (
            .O(N__53509),
            .I(N__53463));
    Span4Mux_h I__13052 (
            .O(N__53506),
            .I(N__53454));
    LocalMux I__13051 (
            .O(N__53503),
            .I(N__53454));
    LocalMux I__13050 (
            .O(N__53500),
            .I(N__53454));
    InMux I__13049 (
            .O(N__53499),
            .I(N__53451));
    InMux I__13048 (
            .O(N__53498),
            .I(N__53439));
    InMux I__13047 (
            .O(N__53497),
            .I(N__53439));
    InMux I__13046 (
            .O(N__53496),
            .I(N__53439));
    InMux I__13045 (
            .O(N__53495),
            .I(N__53439));
    InMux I__13044 (
            .O(N__53494),
            .I(N__53432));
    InMux I__13043 (
            .O(N__53493),
            .I(N__53432));
    InMux I__13042 (
            .O(N__53492),
            .I(N__53421));
    InMux I__13041 (
            .O(N__53491),
            .I(N__53421));
    InMux I__13040 (
            .O(N__53490),
            .I(N__53421));
    InMux I__13039 (
            .O(N__53489),
            .I(N__53421));
    InMux I__13038 (
            .O(N__53488),
            .I(N__53421));
    InMux I__13037 (
            .O(N__53487),
            .I(N__53418));
    InMux I__13036 (
            .O(N__53486),
            .I(N__53414));
    InMux I__13035 (
            .O(N__53485),
            .I(N__53411));
    InMux I__13034 (
            .O(N__53482),
            .I(N__53408));
    LocalMux I__13033 (
            .O(N__53479),
            .I(N__53403));
    Span4Mux_v I__13032 (
            .O(N__53476),
            .I(N__53403));
    InMux I__13031 (
            .O(N__53475),
            .I(N__53398));
    InMux I__13030 (
            .O(N__53474),
            .I(N__53398));
    LocalMux I__13029 (
            .O(N__53467),
            .I(N__53395));
    InMux I__13028 (
            .O(N__53466),
            .I(N__53392));
    LocalMux I__13027 (
            .O(N__53463),
            .I(N__53389));
    InMux I__13026 (
            .O(N__53462),
            .I(N__53384));
    InMux I__13025 (
            .O(N__53461),
            .I(N__53384));
    Span4Mux_v I__13024 (
            .O(N__53454),
            .I(N__53379));
    LocalMux I__13023 (
            .O(N__53451),
            .I(N__53379));
    InMux I__13022 (
            .O(N__53450),
            .I(N__53372));
    InMux I__13021 (
            .O(N__53449),
            .I(N__53372));
    InMux I__13020 (
            .O(N__53448),
            .I(N__53372));
    LocalMux I__13019 (
            .O(N__53439),
            .I(N__53368));
    InMux I__13018 (
            .O(N__53438),
            .I(N__53365));
    InMux I__13017 (
            .O(N__53437),
            .I(N__53362));
    LocalMux I__13016 (
            .O(N__53432),
            .I(N__53358));
    LocalMux I__13015 (
            .O(N__53421),
            .I(N__53353));
    LocalMux I__13014 (
            .O(N__53418),
            .I(N__53353));
    InMux I__13013 (
            .O(N__53417),
            .I(N__53350));
    LocalMux I__13012 (
            .O(N__53414),
            .I(N__53345));
    LocalMux I__13011 (
            .O(N__53411),
            .I(N__53345));
    LocalMux I__13010 (
            .O(N__53408),
            .I(N__53340));
    Span4Mux_h I__13009 (
            .O(N__53403),
            .I(N__53340));
    LocalMux I__13008 (
            .O(N__53398),
            .I(N__53337));
    Span4Mux_v I__13007 (
            .O(N__53395),
            .I(N__53332));
    LocalMux I__13006 (
            .O(N__53392),
            .I(N__53332));
    Sp12to4 I__13005 (
            .O(N__53389),
            .I(N__53327));
    LocalMux I__13004 (
            .O(N__53384),
            .I(N__53327));
    Span4Mux_h I__13003 (
            .O(N__53379),
            .I(N__53324));
    LocalMux I__13002 (
            .O(N__53372),
            .I(N__53321));
    InMux I__13001 (
            .O(N__53371),
            .I(N__53318));
    Span4Mux_h I__13000 (
            .O(N__53368),
            .I(N__53311));
    LocalMux I__12999 (
            .O(N__53365),
            .I(N__53311));
    LocalMux I__12998 (
            .O(N__53362),
            .I(N__53311));
    InMux I__12997 (
            .O(N__53361),
            .I(N__53308));
    Span4Mux_v I__12996 (
            .O(N__53358),
            .I(N__53303));
    Span4Mux_v I__12995 (
            .O(N__53353),
            .I(N__53303));
    LocalMux I__12994 (
            .O(N__53350),
            .I(N__53300));
    Span4Mux_v I__12993 (
            .O(N__53345),
            .I(N__53291));
    Span4Mux_h I__12992 (
            .O(N__53340),
            .I(N__53291));
    Span4Mux_v I__12991 (
            .O(N__53337),
            .I(N__53291));
    Span4Mux_v I__12990 (
            .O(N__53332),
            .I(N__53291));
    Span12Mux_v I__12989 (
            .O(N__53327),
            .I(N__53288));
    Span4Mux_h I__12988 (
            .O(N__53324),
            .I(N__53285));
    Odrv12 I__12987 (
            .O(N__53321),
            .I(comm_state_0));
    LocalMux I__12986 (
            .O(N__53318),
            .I(comm_state_0));
    Odrv4 I__12985 (
            .O(N__53311),
            .I(comm_state_0));
    LocalMux I__12984 (
            .O(N__53308),
            .I(comm_state_0));
    Odrv4 I__12983 (
            .O(N__53303),
            .I(comm_state_0));
    Odrv4 I__12982 (
            .O(N__53300),
            .I(comm_state_0));
    Odrv4 I__12981 (
            .O(N__53291),
            .I(comm_state_0));
    Odrv12 I__12980 (
            .O(N__53288),
            .I(comm_state_0));
    Odrv4 I__12979 (
            .O(N__53285),
            .I(comm_state_0));
    CEMux I__12978 (
            .O(N__53266),
            .I(N__53263));
    LocalMux I__12977 (
            .O(N__53263),
            .I(n11347));
    InMux I__12976 (
            .O(N__53260),
            .I(N__53255));
    InMux I__12975 (
            .O(N__53259),
            .I(N__53250));
    InMux I__12974 (
            .O(N__53258),
            .I(N__53250));
    LocalMux I__12973 (
            .O(N__53255),
            .I(N__53247));
    LocalMux I__12972 (
            .O(N__53250),
            .I(N__53244));
    Span4Mux_v I__12971 (
            .O(N__53247),
            .I(N__53239));
    Span4Mux_v I__12970 (
            .O(N__53244),
            .I(N__53239));
    Span4Mux_h I__12969 (
            .O(N__53239),
            .I(N__53236));
    Odrv4 I__12968 (
            .O(N__53236),
            .I(comm_tx_buf_0));
    InMux I__12967 (
            .O(N__53233),
            .I(N__53230));
    LocalMux I__12966 (
            .O(N__53230),
            .I(N__53225));
    InMux I__12965 (
            .O(N__53229),
            .I(N__53222));
    InMux I__12964 (
            .O(N__53228),
            .I(N__53219));
    Odrv4 I__12963 (
            .O(N__53225),
            .I(\comm_spi.n22650 ));
    LocalMux I__12962 (
            .O(N__53222),
            .I(\comm_spi.n22650 ));
    LocalMux I__12961 (
            .O(N__53219),
            .I(\comm_spi.n22650 ));
    SRMux I__12960 (
            .O(N__53212),
            .I(N__53209));
    LocalMux I__12959 (
            .O(N__53209),
            .I(N__53206));
    Span4Mux_v I__12958 (
            .O(N__53206),
            .I(N__53203));
    Odrv4 I__12957 (
            .O(N__53203),
            .I(\comm_spi.data_tx_7__N_764 ));
    InMux I__12956 (
            .O(N__53200),
            .I(N__53194));
    InMux I__12955 (
            .O(N__53199),
            .I(N__53194));
    LocalMux I__12954 (
            .O(N__53194),
            .I(N__53190));
    InMux I__12953 (
            .O(N__53193),
            .I(N__53187));
    Span4Mux_v I__12952 (
            .O(N__53190),
            .I(N__53184));
    LocalMux I__12951 (
            .O(N__53187),
            .I(N__53181));
    Odrv4 I__12950 (
            .O(N__53184),
            .I(comm_tx_buf_1));
    Odrv4 I__12949 (
            .O(N__53181),
            .I(comm_tx_buf_1));
    SRMux I__12948 (
            .O(N__53176),
            .I(N__53173));
    LocalMux I__12947 (
            .O(N__53173),
            .I(N__53170));
    Sp12to4 I__12946 (
            .O(N__53170),
            .I(N__53167));
    Odrv12 I__12945 (
            .O(N__53167),
            .I(\comm_spi.data_tx_7__N_784 ));
    InMux I__12944 (
            .O(N__53164),
            .I(N__53161));
    LocalMux I__12943 (
            .O(N__53161),
            .I(N__53157));
    InMux I__12942 (
            .O(N__53160),
            .I(N__53154));
    Span4Mux_h I__12941 (
            .O(N__53157),
            .I(N__53149));
    LocalMux I__12940 (
            .O(N__53154),
            .I(N__53149));
    Span4Mux_v I__12939 (
            .O(N__53149),
            .I(N__53145));
    InMux I__12938 (
            .O(N__53148),
            .I(N__53142));
    Span4Mux_h I__12937 (
            .O(N__53145),
            .I(N__53139));
    LocalMux I__12936 (
            .O(N__53142),
            .I(N__53136));
    Odrv4 I__12935 (
            .O(N__53139),
            .I(comm_tx_buf_4));
    Odrv4 I__12934 (
            .O(N__53136),
            .I(comm_tx_buf_4));
    SRMux I__12933 (
            .O(N__53131),
            .I(N__53128));
    LocalMux I__12932 (
            .O(N__53128),
            .I(N__53125));
    Span4Mux_v I__12931 (
            .O(N__53125),
            .I(N__53122));
    Odrv4 I__12930 (
            .O(N__53122),
            .I(\comm_spi.data_tx_7__N_775 ));
    CascadeMux I__12929 (
            .O(N__53119),
            .I(n20502_cascade_));
    InMux I__12928 (
            .O(N__53116),
            .I(N__53113));
    LocalMux I__12927 (
            .O(N__53113),
            .I(n12_adj_1583));
    InMux I__12926 (
            .O(N__53110),
            .I(N__53107));
    LocalMux I__12925 (
            .O(N__53107),
            .I(n20502));
    InMux I__12924 (
            .O(N__53104),
            .I(N__53100));
    InMux I__12923 (
            .O(N__53103),
            .I(N__53097));
    LocalMux I__12922 (
            .O(N__53100),
            .I(N__53094));
    LocalMux I__12921 (
            .O(N__53097),
            .I(secclk_cnt_19));
    Odrv12 I__12920 (
            .O(N__53094),
            .I(secclk_cnt_19));
    InMux I__12919 (
            .O(N__53089),
            .I(N__53085));
    InMux I__12918 (
            .O(N__53088),
            .I(N__53082));
    LocalMux I__12917 (
            .O(N__53085),
            .I(N__53079));
    LocalMux I__12916 (
            .O(N__53082),
            .I(secclk_cnt_21));
    Odrv12 I__12915 (
            .O(N__53079),
            .I(secclk_cnt_21));
    CascadeMux I__12914 (
            .O(N__53074),
            .I(N__53071));
    InMux I__12913 (
            .O(N__53071),
            .I(N__53068));
    LocalMux I__12912 (
            .O(N__53068),
            .I(N__53064));
    InMux I__12911 (
            .O(N__53067),
            .I(N__53061));
    Span4Mux_v I__12910 (
            .O(N__53064),
            .I(N__53058));
    LocalMux I__12909 (
            .O(N__53061),
            .I(secclk_cnt_12));
    Odrv4 I__12908 (
            .O(N__53058),
            .I(secclk_cnt_12));
    InMux I__12907 (
            .O(N__53053),
            .I(N__53049));
    InMux I__12906 (
            .O(N__53052),
            .I(N__53046));
    LocalMux I__12905 (
            .O(N__53049),
            .I(N__53043));
    LocalMux I__12904 (
            .O(N__53046),
            .I(secclk_cnt_22));
    Odrv12 I__12903 (
            .O(N__53043),
            .I(secclk_cnt_22));
    InMux I__12902 (
            .O(N__53038),
            .I(N__53035));
    LocalMux I__12901 (
            .O(N__53035),
            .I(N__53032));
    Span4Mux_h I__12900 (
            .O(N__53032),
            .I(N__53029));
    Odrv4 I__12899 (
            .O(N__53029),
            .I(n14_adj_1578));
    CascadeMux I__12898 (
            .O(N__53026),
            .I(N__53022));
    CascadeMux I__12897 (
            .O(N__53025),
            .I(N__53019));
    InMux I__12896 (
            .O(N__53022),
            .I(N__53015));
    InMux I__12895 (
            .O(N__53019),
            .I(N__53012));
    CascadeMux I__12894 (
            .O(N__53018),
            .I(N__53009));
    LocalMux I__12893 (
            .O(N__53015),
            .I(N__53006));
    LocalMux I__12892 (
            .O(N__53012),
            .I(N__53002));
    InMux I__12891 (
            .O(N__53009),
            .I(N__52999));
    Span4Mux_h I__12890 (
            .O(N__53006),
            .I(N__52996));
    CascadeMux I__12889 (
            .O(N__53005),
            .I(N__52993));
    Span4Mux_h I__12888 (
            .O(N__53002),
            .I(N__52990));
    LocalMux I__12887 (
            .O(N__52999),
            .I(N__52985));
    Span4Mux_h I__12886 (
            .O(N__52996),
            .I(N__52985));
    InMux I__12885 (
            .O(N__52993),
            .I(N__52982));
    Span4Mux_h I__12884 (
            .O(N__52990),
            .I(N__52979));
    Span4Mux_h I__12883 (
            .O(N__52985),
            .I(N__52976));
    LocalMux I__12882 (
            .O(N__52982),
            .I(trig_dds0));
    Odrv4 I__12881 (
            .O(N__52979),
            .I(trig_dds0));
    Odrv4 I__12880 (
            .O(N__52976),
            .I(trig_dds0));
    InMux I__12879 (
            .O(N__52969),
            .I(N__52966));
    LocalMux I__12878 (
            .O(N__52966),
            .I(N__52963));
    Odrv12 I__12877 (
            .O(N__52963),
            .I(\comm_spi.n14582 ));
    InMux I__12876 (
            .O(N__52960),
            .I(N__52957));
    LocalMux I__12875 (
            .O(N__52957),
            .I(N__52954));
    Span4Mux_v I__12874 (
            .O(N__52954),
            .I(N__52949));
    InMux I__12873 (
            .O(N__52953),
            .I(N__52946));
    InMux I__12872 (
            .O(N__52952),
            .I(N__52943));
    Sp12to4 I__12871 (
            .O(N__52949),
            .I(N__52938));
    LocalMux I__12870 (
            .O(N__52946),
            .I(N__52933));
    LocalMux I__12869 (
            .O(N__52943),
            .I(N__52933));
    InMux I__12868 (
            .O(N__52942),
            .I(N__52930));
    InMux I__12867 (
            .O(N__52941),
            .I(N__52927));
    Span12Mux_h I__12866 (
            .O(N__52938),
            .I(N__52924));
    Sp12to4 I__12865 (
            .O(N__52933),
            .I(N__52917));
    LocalMux I__12864 (
            .O(N__52930),
            .I(N__52917));
    LocalMux I__12863 (
            .O(N__52927),
            .I(N__52917));
    Span12Mux_v I__12862 (
            .O(N__52924),
            .I(N__52914));
    Span12Mux_v I__12861 (
            .O(N__52917),
            .I(N__52911));
    Odrv12 I__12860 (
            .O(N__52914),
            .I(ICE_SPI_SCLK));
    Odrv12 I__12859 (
            .O(N__52911),
            .I(ICE_SPI_SCLK));
    SRMux I__12858 (
            .O(N__52906),
            .I(N__52903));
    LocalMux I__12857 (
            .O(N__52903),
            .I(N__52900));
    Odrv4 I__12856 (
            .O(N__52900),
            .I(\comm_spi.iclk_N_755 ));
    SRMux I__12855 (
            .O(N__52897),
            .I(N__52894));
    LocalMux I__12854 (
            .O(N__52894),
            .I(N__52891));
    Odrv4 I__12853 (
            .O(N__52891),
            .I(\comm_spi.data_tx_7__N_765 ));
    SRMux I__12852 (
            .O(N__52888),
            .I(N__52883));
    SRMux I__12851 (
            .O(N__52887),
            .I(N__52880));
    SRMux I__12850 (
            .O(N__52886),
            .I(N__52874));
    LocalMux I__12849 (
            .O(N__52883),
            .I(N__52868));
    LocalMux I__12848 (
            .O(N__52880),
            .I(N__52868));
    SRMux I__12847 (
            .O(N__52879),
            .I(N__52865));
    SRMux I__12846 (
            .O(N__52878),
            .I(N__52862));
    IoInMux I__12845 (
            .O(N__52877),
            .I(N__52857));
    LocalMux I__12844 (
            .O(N__52874),
            .I(N__52854));
    SRMux I__12843 (
            .O(N__52873),
            .I(N__52851));
    Span4Mux_v I__12842 (
            .O(N__52868),
            .I(N__52844));
    LocalMux I__12841 (
            .O(N__52865),
            .I(N__52844));
    LocalMux I__12840 (
            .O(N__52862),
            .I(N__52844));
    SRMux I__12839 (
            .O(N__52861),
            .I(N__52841));
    SRMux I__12838 (
            .O(N__52860),
            .I(N__52838));
    LocalMux I__12837 (
            .O(N__52857),
            .I(N__52832));
    Span4Mux_v I__12836 (
            .O(N__52854),
            .I(N__52823));
    LocalMux I__12835 (
            .O(N__52851),
            .I(N__52823));
    Span4Mux_v I__12834 (
            .O(N__52844),
            .I(N__52816));
    LocalMux I__12833 (
            .O(N__52841),
            .I(N__52816));
    LocalMux I__12832 (
            .O(N__52838),
            .I(N__52816));
    SRMux I__12831 (
            .O(N__52837),
            .I(N__52813));
    SRMux I__12830 (
            .O(N__52836),
            .I(N__52806));
    SRMux I__12829 (
            .O(N__52835),
            .I(N__52796));
    Span4Mux_s0_v I__12828 (
            .O(N__52832),
            .I(N__52788));
    CascadeMux I__12827 (
            .O(N__52831),
            .I(N__52785));
    CascadeMux I__12826 (
            .O(N__52830),
            .I(N__52781));
    CascadeMux I__12825 (
            .O(N__52829),
            .I(N__52777));
    CascadeMux I__12824 (
            .O(N__52828),
            .I(N__52773));
    Span4Mux_h I__12823 (
            .O(N__52823),
            .I(N__52766));
    Span4Mux_v I__12822 (
            .O(N__52816),
            .I(N__52766));
    LocalMux I__12821 (
            .O(N__52813),
            .I(N__52766));
    CascadeMux I__12820 (
            .O(N__52812),
            .I(N__52763));
    CascadeMux I__12819 (
            .O(N__52811),
            .I(N__52759));
    CascadeMux I__12818 (
            .O(N__52810),
            .I(N__52755));
    CascadeMux I__12817 (
            .O(N__52809),
            .I(N__52751));
    LocalMux I__12816 (
            .O(N__52806),
            .I(N__52744));
    InMux I__12815 (
            .O(N__52805),
            .I(N__52737));
    InMux I__12814 (
            .O(N__52804),
            .I(N__52737));
    InMux I__12813 (
            .O(N__52803),
            .I(N__52737));
    InMux I__12812 (
            .O(N__52802),
            .I(N__52728));
    InMux I__12811 (
            .O(N__52801),
            .I(N__52728));
    InMux I__12810 (
            .O(N__52800),
            .I(N__52728));
    InMux I__12809 (
            .O(N__52799),
            .I(N__52728));
    LocalMux I__12808 (
            .O(N__52796),
            .I(N__52725));
    InMux I__12807 (
            .O(N__52795),
            .I(N__52720));
    CascadeMux I__12806 (
            .O(N__52794),
            .I(N__52716));
    CascadeMux I__12805 (
            .O(N__52793),
            .I(N__52712));
    CascadeMux I__12804 (
            .O(N__52792),
            .I(N__52708));
    CascadeMux I__12803 (
            .O(N__52791),
            .I(N__52704));
    Span4Mux_v I__12802 (
            .O(N__52788),
            .I(N__52701));
    InMux I__12801 (
            .O(N__52785),
            .I(N__52686));
    InMux I__12800 (
            .O(N__52784),
            .I(N__52686));
    InMux I__12799 (
            .O(N__52781),
            .I(N__52686));
    InMux I__12798 (
            .O(N__52780),
            .I(N__52686));
    InMux I__12797 (
            .O(N__52777),
            .I(N__52686));
    InMux I__12796 (
            .O(N__52776),
            .I(N__52686));
    InMux I__12795 (
            .O(N__52773),
            .I(N__52686));
    Span4Mux_v I__12794 (
            .O(N__52766),
            .I(N__52683));
    InMux I__12793 (
            .O(N__52763),
            .I(N__52668));
    InMux I__12792 (
            .O(N__52762),
            .I(N__52668));
    InMux I__12791 (
            .O(N__52759),
            .I(N__52668));
    InMux I__12790 (
            .O(N__52758),
            .I(N__52668));
    InMux I__12789 (
            .O(N__52755),
            .I(N__52668));
    InMux I__12788 (
            .O(N__52754),
            .I(N__52668));
    InMux I__12787 (
            .O(N__52751),
            .I(N__52668));
    CascadeMux I__12786 (
            .O(N__52750),
            .I(N__52664));
    CascadeMux I__12785 (
            .O(N__52749),
            .I(N__52660));
    CascadeMux I__12784 (
            .O(N__52748),
            .I(N__52656));
    CascadeMux I__12783 (
            .O(N__52747),
            .I(N__52652));
    Span4Mux_v I__12782 (
            .O(N__52744),
            .I(N__52649));
    LocalMux I__12781 (
            .O(N__52737),
            .I(N__52644));
    LocalMux I__12780 (
            .O(N__52728),
            .I(N__52644));
    Span4Mux_v I__12779 (
            .O(N__52725),
            .I(N__52641));
    InMux I__12778 (
            .O(N__52724),
            .I(N__52638));
    SRMux I__12777 (
            .O(N__52723),
            .I(N__52635));
    LocalMux I__12776 (
            .O(N__52720),
            .I(N__52632));
    InMux I__12775 (
            .O(N__52719),
            .I(N__52615));
    InMux I__12774 (
            .O(N__52716),
            .I(N__52615));
    InMux I__12773 (
            .O(N__52715),
            .I(N__52615));
    InMux I__12772 (
            .O(N__52712),
            .I(N__52615));
    InMux I__12771 (
            .O(N__52711),
            .I(N__52615));
    InMux I__12770 (
            .O(N__52708),
            .I(N__52615));
    InMux I__12769 (
            .O(N__52707),
            .I(N__52615));
    InMux I__12768 (
            .O(N__52704),
            .I(N__52615));
    Span4Mux_v I__12767 (
            .O(N__52701),
            .I(N__52610));
    LocalMux I__12766 (
            .O(N__52686),
            .I(N__52610));
    Span4Mux_h I__12765 (
            .O(N__52683),
            .I(N__52605));
    LocalMux I__12764 (
            .O(N__52668),
            .I(N__52605));
    InMux I__12763 (
            .O(N__52667),
            .I(N__52588));
    InMux I__12762 (
            .O(N__52664),
            .I(N__52588));
    InMux I__12761 (
            .O(N__52663),
            .I(N__52588));
    InMux I__12760 (
            .O(N__52660),
            .I(N__52588));
    InMux I__12759 (
            .O(N__52659),
            .I(N__52588));
    InMux I__12758 (
            .O(N__52656),
            .I(N__52588));
    InMux I__12757 (
            .O(N__52655),
            .I(N__52588));
    InMux I__12756 (
            .O(N__52652),
            .I(N__52588));
    Span4Mux_h I__12755 (
            .O(N__52649),
            .I(N__52585));
    Span4Mux_v I__12754 (
            .O(N__52644),
            .I(N__52582));
    Sp12to4 I__12753 (
            .O(N__52641),
            .I(N__52577));
    LocalMux I__12752 (
            .O(N__52638),
            .I(N__52577));
    LocalMux I__12751 (
            .O(N__52635),
            .I(N__52574));
    Span4Mux_v I__12750 (
            .O(N__52632),
            .I(N__52571));
    LocalMux I__12749 (
            .O(N__52615),
            .I(N__52568));
    Span4Mux_h I__12748 (
            .O(N__52610),
            .I(N__52561));
    Span4Mux_h I__12747 (
            .O(N__52605),
            .I(N__52561));
    LocalMux I__12746 (
            .O(N__52588),
            .I(N__52561));
    Span4Mux_h I__12745 (
            .O(N__52585),
            .I(N__52556));
    Span4Mux_v I__12744 (
            .O(N__52582),
            .I(N__52556));
    Span12Mux_s10_h I__12743 (
            .O(N__52577),
            .I(N__52551));
    Span12Mux_s9_h I__12742 (
            .O(N__52574),
            .I(N__52551));
    Span4Mux_h I__12741 (
            .O(N__52571),
            .I(N__52546));
    Span4Mux_v I__12740 (
            .O(N__52568),
            .I(N__52546));
    Sp12to4 I__12739 (
            .O(N__52561),
            .I(N__52543));
    Odrv4 I__12738 (
            .O(N__52556),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__12737 (
            .O(N__52551),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__12736 (
            .O(N__52546),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__12735 (
            .O(N__52543),
            .I(CONSTANT_ONE_NET));
    SRMux I__12734 (
            .O(N__52534),
            .I(N__52531));
    LocalMux I__12733 (
            .O(N__52531),
            .I(N__52528));
    Sp12to4 I__12732 (
            .O(N__52528),
            .I(N__52525));
    Odrv12 I__12731 (
            .O(N__52525),
            .I(\comm_spi.data_tx_7__N_787 ));
    InMux I__12730 (
            .O(N__52522),
            .I(N__52519));
    LocalMux I__12729 (
            .O(N__52519),
            .I(N__52515));
    InMux I__12728 (
            .O(N__52518),
            .I(N__52512));
    Span4Mux_v I__12727 (
            .O(N__52515),
            .I(N__52507));
    LocalMux I__12726 (
            .O(N__52512),
            .I(N__52507));
    Span4Mux_h I__12725 (
            .O(N__52507),
            .I(N__52504));
    Odrv4 I__12724 (
            .O(N__52504),
            .I(\comm_spi.n14604 ));
    InMux I__12723 (
            .O(N__52501),
            .I(N__52498));
    LocalMux I__12722 (
            .O(N__52498),
            .I(N__52494));
    InMux I__12721 (
            .O(N__52497),
            .I(N__52491));
    Odrv4 I__12720 (
            .O(N__52494),
            .I(\comm_spi.n14578 ));
    LocalMux I__12719 (
            .O(N__52491),
            .I(\comm_spi.n14578 ));
    InMux I__12718 (
            .O(N__52486),
            .I(N__52483));
    LocalMux I__12717 (
            .O(N__52483),
            .I(N__52479));
    InMux I__12716 (
            .O(N__52482),
            .I(N__52476));
    Span4Mux_v I__12715 (
            .O(N__52479),
            .I(N__52471));
    LocalMux I__12714 (
            .O(N__52476),
            .I(N__52471));
    Odrv4 I__12713 (
            .O(N__52471),
            .I(\comm_spi.n14577 ));
    InMux I__12712 (
            .O(N__52468),
            .I(N__52465));
    LocalMux I__12711 (
            .O(N__52465),
            .I(N__52462));
    Span4Mux_h I__12710 (
            .O(N__52462),
            .I(N__52458));
    InMux I__12709 (
            .O(N__52461),
            .I(N__52455));
    Span4Mux_h I__12708 (
            .O(N__52458),
            .I(N__52452));
    LocalMux I__12707 (
            .O(N__52455),
            .I(N__52449));
    Odrv4 I__12706 (
            .O(N__52452),
            .I(\comm_spi.n14603 ));
    Odrv12 I__12705 (
            .O(N__52449),
            .I(\comm_spi.n14603 ));
    ClkMux I__12704 (
            .O(N__52444),
            .I(N__52438));
    ClkMux I__12703 (
            .O(N__52443),
            .I(N__52434));
    ClkMux I__12702 (
            .O(N__52442),
            .I(N__52431));
    ClkMux I__12701 (
            .O(N__52441),
            .I(N__52427));
    LocalMux I__12700 (
            .O(N__52438),
            .I(N__52421));
    ClkMux I__12699 (
            .O(N__52437),
            .I(N__52418));
    LocalMux I__12698 (
            .O(N__52434),
            .I(N__52408));
    LocalMux I__12697 (
            .O(N__52431),
            .I(N__52408));
    ClkMux I__12696 (
            .O(N__52430),
            .I(N__52404));
    LocalMux I__12695 (
            .O(N__52427),
            .I(N__52401));
    ClkMux I__12694 (
            .O(N__52426),
            .I(N__52398));
    ClkMux I__12693 (
            .O(N__52425),
            .I(N__52395));
    ClkMux I__12692 (
            .O(N__52424),
            .I(N__52392));
    Span4Mux_v I__12691 (
            .O(N__52421),
            .I(N__52386));
    LocalMux I__12690 (
            .O(N__52418),
            .I(N__52386));
    ClkMux I__12689 (
            .O(N__52417),
            .I(N__52383));
    ClkMux I__12688 (
            .O(N__52416),
            .I(N__52380));
    ClkMux I__12687 (
            .O(N__52415),
            .I(N__52376));
    ClkMux I__12686 (
            .O(N__52414),
            .I(N__52372));
    ClkMux I__12685 (
            .O(N__52413),
            .I(N__52369));
    Span4Mux_v I__12684 (
            .O(N__52408),
            .I(N__52365));
    ClkMux I__12683 (
            .O(N__52407),
            .I(N__52361));
    LocalMux I__12682 (
            .O(N__52404),
            .I(N__52353));
    Span4Mux_h I__12681 (
            .O(N__52401),
            .I(N__52353));
    LocalMux I__12680 (
            .O(N__52398),
            .I(N__52353));
    LocalMux I__12679 (
            .O(N__52395),
            .I(N__52348));
    LocalMux I__12678 (
            .O(N__52392),
            .I(N__52348));
    ClkMux I__12677 (
            .O(N__52391),
            .I(N__52345));
    Span4Mux_v I__12676 (
            .O(N__52386),
            .I(N__52340));
    LocalMux I__12675 (
            .O(N__52383),
            .I(N__52340));
    LocalMux I__12674 (
            .O(N__52380),
            .I(N__52337));
    ClkMux I__12673 (
            .O(N__52379),
            .I(N__52334));
    LocalMux I__12672 (
            .O(N__52376),
            .I(N__52331));
    ClkMux I__12671 (
            .O(N__52375),
            .I(N__52328));
    LocalMux I__12670 (
            .O(N__52372),
            .I(N__52323));
    LocalMux I__12669 (
            .O(N__52369),
            .I(N__52323));
    ClkMux I__12668 (
            .O(N__52368),
            .I(N__52320));
    Span4Mux_h I__12667 (
            .O(N__52365),
            .I(N__52316));
    ClkMux I__12666 (
            .O(N__52364),
            .I(N__52313));
    LocalMux I__12665 (
            .O(N__52361),
            .I(N__52310));
    ClkMux I__12664 (
            .O(N__52360),
            .I(N__52307));
    Span4Mux_v I__12663 (
            .O(N__52353),
            .I(N__52304));
    Span4Mux_h I__12662 (
            .O(N__52348),
            .I(N__52293));
    LocalMux I__12661 (
            .O(N__52345),
            .I(N__52293));
    Span4Mux_h I__12660 (
            .O(N__52340),
            .I(N__52293));
    Span4Mux_v I__12659 (
            .O(N__52337),
            .I(N__52293));
    LocalMux I__12658 (
            .O(N__52334),
            .I(N__52293));
    Span4Mux_v I__12657 (
            .O(N__52331),
            .I(N__52288));
    LocalMux I__12656 (
            .O(N__52328),
            .I(N__52288));
    Span4Mux_v I__12655 (
            .O(N__52323),
            .I(N__52283));
    LocalMux I__12654 (
            .O(N__52320),
            .I(N__52283));
    ClkMux I__12653 (
            .O(N__52319),
            .I(N__52280));
    Span4Mux_v I__12652 (
            .O(N__52316),
            .I(N__52277));
    LocalMux I__12651 (
            .O(N__52313),
            .I(N__52274));
    Span4Mux_h I__12650 (
            .O(N__52310),
            .I(N__52267));
    LocalMux I__12649 (
            .O(N__52307),
            .I(N__52267));
    Span4Mux_h I__12648 (
            .O(N__52304),
            .I(N__52267));
    Span4Mux_v I__12647 (
            .O(N__52293),
            .I(N__52264));
    Span4Mux_h I__12646 (
            .O(N__52288),
            .I(N__52257));
    Span4Mux_h I__12645 (
            .O(N__52283),
            .I(N__52257));
    LocalMux I__12644 (
            .O(N__52280),
            .I(N__52257));
    Odrv4 I__12643 (
            .O(N__52277),
            .I(\comm_spi.iclk ));
    Odrv12 I__12642 (
            .O(N__52274),
            .I(\comm_spi.iclk ));
    Odrv4 I__12641 (
            .O(N__52267),
            .I(\comm_spi.iclk ));
    Odrv4 I__12640 (
            .O(N__52264),
            .I(\comm_spi.iclk ));
    Odrv4 I__12639 (
            .O(N__52257),
            .I(\comm_spi.iclk ));
    InMux I__12638 (
            .O(N__52246),
            .I(N__52243));
    LocalMux I__12637 (
            .O(N__52243),
            .I(N__52240));
    Span4Mux_h I__12636 (
            .O(N__52240),
            .I(N__52237));
    Odrv4 I__12635 (
            .O(N__52237),
            .I(n20863));
    InMux I__12634 (
            .O(N__52234),
            .I(N__52229));
    InMux I__12633 (
            .O(N__52233),
            .I(N__52226));
    CascadeMux I__12632 (
            .O(N__52232),
            .I(N__52223));
    LocalMux I__12631 (
            .O(N__52229),
            .I(N__52220));
    LocalMux I__12630 (
            .O(N__52226),
            .I(N__52217));
    InMux I__12629 (
            .O(N__52223),
            .I(N__52214));
    Span4Mux_h I__12628 (
            .O(N__52220),
            .I(N__52211));
    Span4Mux_h I__12627 (
            .O(N__52217),
            .I(N__52208));
    LocalMux I__12626 (
            .O(N__52214),
            .I(N__52205));
    Odrv4 I__12625 (
            .O(N__52211),
            .I(n14514));
    Odrv4 I__12624 (
            .O(N__52208),
            .I(n14514));
    Odrv4 I__12623 (
            .O(N__52205),
            .I(n14514));
    CascadeMux I__12622 (
            .O(N__52198),
            .I(n21658_cascade_));
    InMux I__12621 (
            .O(N__52195),
            .I(N__52186));
    CascadeMux I__12620 (
            .O(N__52194),
            .I(N__52182));
    CascadeMux I__12619 (
            .O(N__52193),
            .I(N__52178));
    CascadeMux I__12618 (
            .O(N__52192),
            .I(N__52163));
    InMux I__12617 (
            .O(N__52191),
            .I(N__52151));
    InMux I__12616 (
            .O(N__52190),
            .I(N__52151));
    InMux I__12615 (
            .O(N__52189),
            .I(N__52151));
    LocalMux I__12614 (
            .O(N__52186),
            .I(N__52148));
    InMux I__12613 (
            .O(N__52185),
            .I(N__52140));
    InMux I__12612 (
            .O(N__52182),
            .I(N__52140));
    InMux I__12611 (
            .O(N__52181),
            .I(N__52140));
    InMux I__12610 (
            .O(N__52178),
            .I(N__52135));
    InMux I__12609 (
            .O(N__52177),
            .I(N__52135));
    InMux I__12608 (
            .O(N__52176),
            .I(N__52132));
    InMux I__12607 (
            .O(N__52175),
            .I(N__52125));
    InMux I__12606 (
            .O(N__52174),
            .I(N__52125));
    InMux I__12605 (
            .O(N__52173),
            .I(N__52125));
    CascadeMux I__12604 (
            .O(N__52172),
            .I(N__52120));
    CascadeMux I__12603 (
            .O(N__52171),
            .I(N__52117));
    CascadeMux I__12602 (
            .O(N__52170),
            .I(N__52114));
    InMux I__12601 (
            .O(N__52169),
            .I(N__52105));
    InMux I__12600 (
            .O(N__52168),
            .I(N__52102));
    CascadeMux I__12599 (
            .O(N__52167),
            .I(N__52099));
    CascadeMux I__12598 (
            .O(N__52166),
            .I(N__52096));
    InMux I__12597 (
            .O(N__52163),
            .I(N__52093));
    InMux I__12596 (
            .O(N__52162),
            .I(N__52088));
    CascadeMux I__12595 (
            .O(N__52161),
            .I(N__52084));
    CascadeMux I__12594 (
            .O(N__52160),
            .I(N__52081));
    CascadeMux I__12593 (
            .O(N__52159),
            .I(N__52078));
    CascadeMux I__12592 (
            .O(N__52158),
            .I(N__52074));
    LocalMux I__12591 (
            .O(N__52151),
            .I(N__52069));
    Span4Mux_v I__12590 (
            .O(N__52148),
            .I(N__52069));
    CascadeMux I__12589 (
            .O(N__52147),
            .I(N__52066));
    LocalMux I__12588 (
            .O(N__52140),
            .I(N__52050));
    LocalMux I__12587 (
            .O(N__52135),
            .I(N__52050));
    LocalMux I__12586 (
            .O(N__52132),
            .I(N__52050));
    LocalMux I__12585 (
            .O(N__52125),
            .I(N__52050));
    CascadeMux I__12584 (
            .O(N__52124),
            .I(N__52047));
    CascadeMux I__12583 (
            .O(N__52123),
            .I(N__52044));
    InMux I__12582 (
            .O(N__52120),
            .I(N__52037));
    InMux I__12581 (
            .O(N__52117),
            .I(N__52037));
    InMux I__12580 (
            .O(N__52114),
            .I(N__52034));
    CascadeMux I__12579 (
            .O(N__52113),
            .I(N__52030));
    InMux I__12578 (
            .O(N__52112),
            .I(N__52027));
    InMux I__12577 (
            .O(N__52111),
            .I(N__52024));
    InMux I__12576 (
            .O(N__52110),
            .I(N__52017));
    InMux I__12575 (
            .O(N__52109),
            .I(N__52017));
    InMux I__12574 (
            .O(N__52108),
            .I(N__52017));
    LocalMux I__12573 (
            .O(N__52105),
            .I(N__52012));
    LocalMux I__12572 (
            .O(N__52102),
            .I(N__52012));
    InMux I__12571 (
            .O(N__52099),
            .I(N__52007));
    InMux I__12570 (
            .O(N__52096),
            .I(N__52007));
    LocalMux I__12569 (
            .O(N__52093),
            .I(N__52004));
    CascadeMux I__12568 (
            .O(N__52092),
            .I(N__52001));
    CascadeMux I__12567 (
            .O(N__52091),
            .I(N__51998));
    LocalMux I__12566 (
            .O(N__52088),
            .I(N__51995));
    InMux I__12565 (
            .O(N__52087),
            .I(N__51986));
    InMux I__12564 (
            .O(N__52084),
            .I(N__51986));
    InMux I__12563 (
            .O(N__52081),
            .I(N__51986));
    InMux I__12562 (
            .O(N__52078),
            .I(N__51986));
    CascadeMux I__12561 (
            .O(N__52077),
            .I(N__51980));
    InMux I__12560 (
            .O(N__52074),
            .I(N__51971));
    Span4Mux_h I__12559 (
            .O(N__52069),
            .I(N__51968));
    InMux I__12558 (
            .O(N__52066),
            .I(N__51963));
    InMux I__12557 (
            .O(N__52065),
            .I(N__51963));
    InMux I__12556 (
            .O(N__52064),
            .I(N__51958));
    InMux I__12555 (
            .O(N__52063),
            .I(N__51958));
    CascadeMux I__12554 (
            .O(N__52062),
            .I(N__51955));
    CascadeMux I__12553 (
            .O(N__52061),
            .I(N__51952));
    InMux I__12552 (
            .O(N__52060),
            .I(N__51945));
    InMux I__12551 (
            .O(N__52059),
            .I(N__51945));
    Span4Mux_v I__12550 (
            .O(N__52050),
            .I(N__51942));
    InMux I__12549 (
            .O(N__52047),
            .I(N__51937));
    InMux I__12548 (
            .O(N__52044),
            .I(N__51937));
    CascadeMux I__12547 (
            .O(N__52043),
            .I(N__51934));
    CascadeMux I__12546 (
            .O(N__52042),
            .I(N__51931));
    LocalMux I__12545 (
            .O(N__52037),
            .I(N__51924));
    LocalMux I__12544 (
            .O(N__52034),
            .I(N__51924));
    CascadeMux I__12543 (
            .O(N__52033),
            .I(N__51921));
    InMux I__12542 (
            .O(N__52030),
            .I(N__51916));
    LocalMux I__12541 (
            .O(N__52027),
            .I(N__51907));
    LocalMux I__12540 (
            .O(N__52024),
            .I(N__51907));
    LocalMux I__12539 (
            .O(N__52017),
            .I(N__51907));
    Span4Mux_v I__12538 (
            .O(N__52012),
            .I(N__51900));
    LocalMux I__12537 (
            .O(N__52007),
            .I(N__51900));
    Span4Mux_v I__12536 (
            .O(N__52004),
            .I(N__51900));
    InMux I__12535 (
            .O(N__52001),
            .I(N__51895));
    InMux I__12534 (
            .O(N__51998),
            .I(N__51895));
    Span4Mux_h I__12533 (
            .O(N__51995),
            .I(N__51888));
    LocalMux I__12532 (
            .O(N__51986),
            .I(N__51888));
    CascadeMux I__12531 (
            .O(N__51985),
            .I(N__51885));
    CascadeMux I__12530 (
            .O(N__51984),
            .I(N__51882));
    InMux I__12529 (
            .O(N__51983),
            .I(N__51878));
    InMux I__12528 (
            .O(N__51980),
            .I(N__51873));
    InMux I__12527 (
            .O(N__51979),
            .I(N__51873));
    InMux I__12526 (
            .O(N__51978),
            .I(N__51870));
    InMux I__12525 (
            .O(N__51977),
            .I(N__51861));
    InMux I__12524 (
            .O(N__51976),
            .I(N__51861));
    InMux I__12523 (
            .O(N__51975),
            .I(N__51861));
    InMux I__12522 (
            .O(N__51974),
            .I(N__51861));
    LocalMux I__12521 (
            .O(N__51971),
            .I(N__51852));
    Span4Mux_h I__12520 (
            .O(N__51968),
            .I(N__51852));
    LocalMux I__12519 (
            .O(N__51963),
            .I(N__51852));
    LocalMux I__12518 (
            .O(N__51958),
            .I(N__51852));
    InMux I__12517 (
            .O(N__51955),
            .I(N__51849));
    InMux I__12516 (
            .O(N__51952),
            .I(N__51842));
    InMux I__12515 (
            .O(N__51951),
            .I(N__51842));
    InMux I__12514 (
            .O(N__51950),
            .I(N__51842));
    LocalMux I__12513 (
            .O(N__51945),
            .I(N__51835));
    Span4Mux_h I__12512 (
            .O(N__51942),
            .I(N__51835));
    LocalMux I__12511 (
            .O(N__51937),
            .I(N__51835));
    InMux I__12510 (
            .O(N__51934),
            .I(N__51826));
    InMux I__12509 (
            .O(N__51931),
            .I(N__51826));
    InMux I__12508 (
            .O(N__51930),
            .I(N__51826));
    InMux I__12507 (
            .O(N__51929),
            .I(N__51826));
    Span4Mux_h I__12506 (
            .O(N__51924),
            .I(N__51823));
    InMux I__12505 (
            .O(N__51921),
            .I(N__51818));
    InMux I__12504 (
            .O(N__51920),
            .I(N__51818));
    InMux I__12503 (
            .O(N__51919),
            .I(N__51815));
    LocalMux I__12502 (
            .O(N__51916),
            .I(N__51812));
    InMux I__12501 (
            .O(N__51915),
            .I(N__51807));
    InMux I__12500 (
            .O(N__51914),
            .I(N__51807));
    Span4Mux_v I__12499 (
            .O(N__51907),
            .I(N__51800));
    Span4Mux_h I__12498 (
            .O(N__51900),
            .I(N__51800));
    LocalMux I__12497 (
            .O(N__51895),
            .I(N__51800));
    InMux I__12496 (
            .O(N__51894),
            .I(N__51795));
    InMux I__12495 (
            .O(N__51893),
            .I(N__51795));
    Span4Mux_v I__12494 (
            .O(N__51888),
            .I(N__51792));
    InMux I__12493 (
            .O(N__51885),
            .I(N__51787));
    InMux I__12492 (
            .O(N__51882),
            .I(N__51787));
    InMux I__12491 (
            .O(N__51881),
            .I(N__51783));
    LocalMux I__12490 (
            .O(N__51878),
            .I(N__51763));
    LocalMux I__12489 (
            .O(N__51873),
            .I(N__51763));
    LocalMux I__12488 (
            .O(N__51870),
            .I(N__51763));
    LocalMux I__12487 (
            .O(N__51861),
            .I(N__51763));
    Span4Mux_v I__12486 (
            .O(N__51852),
            .I(N__51763));
    LocalMux I__12485 (
            .O(N__51849),
            .I(N__51763));
    LocalMux I__12484 (
            .O(N__51842),
            .I(N__51763));
    Span4Mux_v I__12483 (
            .O(N__51835),
            .I(N__51763));
    LocalMux I__12482 (
            .O(N__51826),
            .I(N__51763));
    Span4Mux_h I__12481 (
            .O(N__51823),
            .I(N__51758));
    LocalMux I__12480 (
            .O(N__51818),
            .I(N__51758));
    LocalMux I__12479 (
            .O(N__51815),
            .I(N__51755));
    Span4Mux_h I__12478 (
            .O(N__51812),
            .I(N__51752));
    LocalMux I__12477 (
            .O(N__51807),
            .I(N__51747));
    Span4Mux_h I__12476 (
            .O(N__51800),
            .I(N__51747));
    LocalMux I__12475 (
            .O(N__51795),
            .I(N__51740));
    Span4Mux_h I__12474 (
            .O(N__51792),
            .I(N__51740));
    LocalMux I__12473 (
            .O(N__51787),
            .I(N__51740));
    InMux I__12472 (
            .O(N__51786),
            .I(N__51737));
    LocalMux I__12471 (
            .O(N__51783),
            .I(N__51734));
    InMux I__12470 (
            .O(N__51782),
            .I(N__51731));
    Span4Mux_v I__12469 (
            .O(N__51763),
            .I(N__51728));
    Span4Mux_h I__12468 (
            .O(N__51758),
            .I(N__51725));
    Span4Mux_v I__12467 (
            .O(N__51755),
            .I(N__51716));
    Span4Mux_v I__12466 (
            .O(N__51752),
            .I(N__51716));
    Span4Mux_h I__12465 (
            .O(N__51747),
            .I(N__51716));
    Span4Mux_h I__12464 (
            .O(N__51740),
            .I(N__51716));
    LocalMux I__12463 (
            .O(N__51737),
            .I(n9273));
    Odrv4 I__12462 (
            .O(N__51734),
            .I(n9273));
    LocalMux I__12461 (
            .O(N__51731),
            .I(n9273));
    Odrv4 I__12460 (
            .O(N__51728),
            .I(n9273));
    Odrv4 I__12459 (
            .O(N__51725),
            .I(n9273));
    Odrv4 I__12458 (
            .O(N__51716),
            .I(n9273));
    CascadeMux I__12457 (
            .O(N__51703),
            .I(n20865_cascade_));
    CEMux I__12456 (
            .O(N__51700),
            .I(N__51697));
    LocalMux I__12455 (
            .O(N__51697),
            .I(N__51694));
    Span4Mux_v I__12454 (
            .O(N__51694),
            .I(N__51691));
    Span4Mux_h I__12453 (
            .O(N__51691),
            .I(N__51688));
    Odrv4 I__12452 (
            .O(N__51688),
            .I(n20536));
    InMux I__12451 (
            .O(N__51685),
            .I(N__51681));
    InMux I__12450 (
            .O(N__51684),
            .I(N__51678));
    LocalMux I__12449 (
            .O(N__51681),
            .I(N__51674));
    LocalMux I__12448 (
            .O(N__51678),
            .I(N__51671));
    InMux I__12447 (
            .O(N__51677),
            .I(N__51668));
    Span4Mux_v I__12446 (
            .O(N__51674),
            .I(N__51665));
    Span4Mux_v I__12445 (
            .O(N__51671),
            .I(N__51660));
    LocalMux I__12444 (
            .O(N__51668),
            .I(N__51660));
    Sp12to4 I__12443 (
            .O(N__51665),
            .I(N__51656));
    Span4Mux_h I__12442 (
            .O(N__51660),
            .I(N__51653));
    InMux I__12441 (
            .O(N__51659),
            .I(N__51650));
    Odrv12 I__12440 (
            .O(N__51656),
            .I(n10540));
    Odrv4 I__12439 (
            .O(N__51653),
            .I(n10540));
    LocalMux I__12438 (
            .O(N__51650),
            .I(n10540));
    InMux I__12437 (
            .O(N__51643),
            .I(N__51633));
    InMux I__12436 (
            .O(N__51642),
            .I(N__51633));
    InMux I__12435 (
            .O(N__51641),
            .I(N__51610));
    InMux I__12434 (
            .O(N__51640),
            .I(N__51610));
    InMux I__12433 (
            .O(N__51639),
            .I(N__51610));
    InMux I__12432 (
            .O(N__51638),
            .I(N__51610));
    LocalMux I__12431 (
            .O(N__51633),
            .I(N__51607));
    InMux I__12430 (
            .O(N__51632),
            .I(N__51601));
    InMux I__12429 (
            .O(N__51631),
            .I(N__51592));
    InMux I__12428 (
            .O(N__51630),
            .I(N__51592));
    InMux I__12427 (
            .O(N__51629),
            .I(N__51592));
    InMux I__12426 (
            .O(N__51628),
            .I(N__51592));
    InMux I__12425 (
            .O(N__51627),
            .I(N__51583));
    InMux I__12424 (
            .O(N__51626),
            .I(N__51583));
    InMux I__12423 (
            .O(N__51625),
            .I(N__51583));
    InMux I__12422 (
            .O(N__51624),
            .I(N__51583));
    InMux I__12421 (
            .O(N__51623),
            .I(N__51580));
    InMux I__12420 (
            .O(N__51622),
            .I(N__51570));
    InMux I__12419 (
            .O(N__51621),
            .I(N__51570));
    InMux I__12418 (
            .O(N__51620),
            .I(N__51570));
    CascadeMux I__12417 (
            .O(N__51619),
            .I(N__51567));
    LocalMux I__12416 (
            .O(N__51610),
            .I(N__51564));
    Span4Mux_v I__12415 (
            .O(N__51607),
            .I(N__51561));
    InMux I__12414 (
            .O(N__51606),
            .I(N__51554));
    InMux I__12413 (
            .O(N__51605),
            .I(N__51554));
    InMux I__12412 (
            .O(N__51604),
            .I(N__51554));
    LocalMux I__12411 (
            .O(N__51601),
            .I(N__51551));
    LocalMux I__12410 (
            .O(N__51592),
            .I(N__51544));
    LocalMux I__12409 (
            .O(N__51583),
            .I(N__51544));
    LocalMux I__12408 (
            .O(N__51580),
            .I(N__51544));
    InMux I__12407 (
            .O(N__51579),
            .I(N__51541));
    InMux I__12406 (
            .O(N__51578),
            .I(N__51538));
    CascadeMux I__12405 (
            .O(N__51577),
            .I(N__51534));
    LocalMux I__12404 (
            .O(N__51570),
            .I(N__51530));
    InMux I__12403 (
            .O(N__51567),
            .I(N__51526));
    Span4Mux_v I__12402 (
            .O(N__51564),
            .I(N__51519));
    Span4Mux_h I__12401 (
            .O(N__51561),
            .I(N__51519));
    LocalMux I__12400 (
            .O(N__51554),
            .I(N__51519));
    Span4Mux_v I__12399 (
            .O(N__51551),
            .I(N__51510));
    Span4Mux_v I__12398 (
            .O(N__51544),
            .I(N__51510));
    LocalMux I__12397 (
            .O(N__51541),
            .I(N__51505));
    LocalMux I__12396 (
            .O(N__51538),
            .I(N__51505));
    InMux I__12395 (
            .O(N__51537),
            .I(N__51498));
    InMux I__12394 (
            .O(N__51534),
            .I(N__51498));
    InMux I__12393 (
            .O(N__51533),
            .I(N__51498));
    Span12Mux_v I__12392 (
            .O(N__51530),
            .I(N__51495));
    InMux I__12391 (
            .O(N__51529),
            .I(N__51492));
    LocalMux I__12390 (
            .O(N__51526),
            .I(N__51487));
    Span4Mux_h I__12389 (
            .O(N__51519),
            .I(N__51487));
    InMux I__12388 (
            .O(N__51518),
            .I(N__51478));
    InMux I__12387 (
            .O(N__51517),
            .I(N__51478));
    InMux I__12386 (
            .O(N__51516),
            .I(N__51478));
    InMux I__12385 (
            .O(N__51515),
            .I(N__51478));
    Span4Mux_h I__12384 (
            .O(N__51510),
            .I(N__51473));
    Span4Mux_v I__12383 (
            .O(N__51505),
            .I(N__51473));
    LocalMux I__12382 (
            .O(N__51498),
            .I(comm_index_0));
    Odrv12 I__12381 (
            .O(N__51495),
            .I(comm_index_0));
    LocalMux I__12380 (
            .O(N__51492),
            .I(comm_index_0));
    Odrv4 I__12379 (
            .O(N__51487),
            .I(comm_index_0));
    LocalMux I__12378 (
            .O(N__51478),
            .I(comm_index_0));
    Odrv4 I__12377 (
            .O(N__51473),
            .I(comm_index_0));
    InMux I__12376 (
            .O(N__51460),
            .I(N__51457));
    LocalMux I__12375 (
            .O(N__51457),
            .I(n20563));
    InMux I__12374 (
            .O(N__51454),
            .I(N__51451));
    LocalMux I__12373 (
            .O(N__51451),
            .I(N__51448));
    Span4Mux_h I__12372 (
            .O(N__51448),
            .I(N__51445));
    Odrv4 I__12371 (
            .O(N__51445),
            .I(n12_adj_1585));
    InMux I__12370 (
            .O(N__51442),
            .I(N__51439));
    LocalMux I__12369 (
            .O(N__51439),
            .I(N__51435));
    CascadeMux I__12368 (
            .O(N__51438),
            .I(N__51432));
    Span4Mux_v I__12367 (
            .O(N__51435),
            .I(N__51425));
    InMux I__12366 (
            .O(N__51432),
            .I(N__51420));
    InMux I__12365 (
            .O(N__51431),
            .I(N__51420));
    CascadeMux I__12364 (
            .O(N__51430),
            .I(N__51417));
    CascadeMux I__12363 (
            .O(N__51429),
            .I(N__51414));
    InMux I__12362 (
            .O(N__51428),
            .I(N__51411));
    Span4Mux_v I__12361 (
            .O(N__51425),
            .I(N__51406));
    LocalMux I__12360 (
            .O(N__51420),
            .I(N__51406));
    InMux I__12359 (
            .O(N__51417),
            .I(N__51403));
    InMux I__12358 (
            .O(N__51414),
            .I(N__51400));
    LocalMux I__12357 (
            .O(N__51411),
            .I(N__51397));
    Span4Mux_h I__12356 (
            .O(N__51406),
            .I(N__51394));
    LocalMux I__12355 (
            .O(N__51403),
            .I(N__51391));
    LocalMux I__12354 (
            .O(N__51400),
            .I(N__51386));
    Span4Mux_h I__12353 (
            .O(N__51397),
            .I(N__51386));
    Span4Mux_h I__12352 (
            .O(N__51394),
            .I(N__51383));
    Odrv12 I__12351 (
            .O(N__51391),
            .I(comm_buf_1_6));
    Odrv4 I__12350 (
            .O(N__51386),
            .I(comm_buf_1_6));
    Odrv4 I__12349 (
            .O(N__51383),
            .I(comm_buf_1_6));
    InMux I__12348 (
            .O(N__51376),
            .I(N__51372));
    InMux I__12347 (
            .O(N__51375),
            .I(N__51369));
    LocalMux I__12346 (
            .O(N__51372),
            .I(N__51364));
    LocalMux I__12345 (
            .O(N__51369),
            .I(N__51364));
    Span12Mux_h I__12344 (
            .O(N__51364),
            .I(N__51361));
    Odrv12 I__12343 (
            .O(N__51361),
            .I(n14_adj_1526));
    InMux I__12342 (
            .O(N__51358),
            .I(N__51355));
    LocalMux I__12341 (
            .O(N__51355),
            .I(N__51352));
    Span4Mux_v I__12340 (
            .O(N__51352),
            .I(N__51349));
    Span4Mux_v I__12339 (
            .O(N__51349),
            .I(N__51346));
    Sp12to4 I__12338 (
            .O(N__51346),
            .I(N__51343));
    Span12Mux_h I__12337 (
            .O(N__51343),
            .I(N__51339));
    InMux I__12336 (
            .O(N__51342),
            .I(N__51336));
    Odrv12 I__12335 (
            .O(N__51339),
            .I(buf_adcdata_vdc_4));
    LocalMux I__12334 (
            .O(N__51336),
            .I(buf_adcdata_vdc_4));
    InMux I__12333 (
            .O(N__51331),
            .I(N__51327));
    InMux I__12332 (
            .O(N__51330),
            .I(N__51323));
    LocalMux I__12331 (
            .O(N__51327),
            .I(N__51320));
    InMux I__12330 (
            .O(N__51326),
            .I(N__51317));
    LocalMux I__12329 (
            .O(N__51323),
            .I(buf_adcdata_vac_4));
    Odrv4 I__12328 (
            .O(N__51320),
            .I(buf_adcdata_vac_4));
    LocalMux I__12327 (
            .O(N__51317),
            .I(buf_adcdata_vac_4));
    InMux I__12326 (
            .O(N__51310),
            .I(N__51307));
    LocalMux I__12325 (
            .O(N__51307),
            .I(N__51304));
    Span12Mux_h I__12324 (
            .O(N__51304),
            .I(N__51301));
    Odrv12 I__12323 (
            .O(N__51301),
            .I(n19_adj_1605));
    InMux I__12322 (
            .O(N__51298),
            .I(N__51294));
    CascadeMux I__12321 (
            .O(N__51297),
            .I(N__51290));
    LocalMux I__12320 (
            .O(N__51294),
            .I(N__51287));
    InMux I__12319 (
            .O(N__51293),
            .I(N__51279));
    InMux I__12318 (
            .O(N__51290),
            .I(N__51276));
    Span4Mux_v I__12317 (
            .O(N__51287),
            .I(N__51273));
    InMux I__12316 (
            .O(N__51286),
            .I(N__51268));
    InMux I__12315 (
            .O(N__51285),
            .I(N__51268));
    InMux I__12314 (
            .O(N__51284),
            .I(N__51265));
    InMux I__12313 (
            .O(N__51283),
            .I(N__51254));
    InMux I__12312 (
            .O(N__51282),
            .I(N__51254));
    LocalMux I__12311 (
            .O(N__51279),
            .I(N__51251));
    LocalMux I__12310 (
            .O(N__51276),
            .I(N__51244));
    Span4Mux_h I__12309 (
            .O(N__51273),
            .I(N__51244));
    LocalMux I__12308 (
            .O(N__51268),
            .I(N__51244));
    LocalMux I__12307 (
            .O(N__51265),
            .I(N__51241));
    CascadeMux I__12306 (
            .O(N__51264),
            .I(N__51235));
    CascadeMux I__12305 (
            .O(N__51263),
            .I(N__51231));
    InMux I__12304 (
            .O(N__51262),
            .I(N__51222));
    CascadeMux I__12303 (
            .O(N__51261),
            .I(N__51214));
    CascadeMux I__12302 (
            .O(N__51260),
            .I(N__51211));
    CascadeMux I__12301 (
            .O(N__51259),
            .I(N__51201));
    LocalMux I__12300 (
            .O(N__51254),
            .I(N__51193));
    Span4Mux_v I__12299 (
            .O(N__51251),
            .I(N__51186));
    Span4Mux_v I__12298 (
            .O(N__51244),
            .I(N__51186));
    Span4Mux_h I__12297 (
            .O(N__51241),
            .I(N__51186));
    InMux I__12296 (
            .O(N__51240),
            .I(N__51181));
    InMux I__12295 (
            .O(N__51239),
            .I(N__51181));
    InMux I__12294 (
            .O(N__51238),
            .I(N__51178));
    InMux I__12293 (
            .O(N__51235),
            .I(N__51169));
    InMux I__12292 (
            .O(N__51234),
            .I(N__51169));
    InMux I__12291 (
            .O(N__51231),
            .I(N__51169));
    InMux I__12290 (
            .O(N__51230),
            .I(N__51169));
    InMux I__12289 (
            .O(N__51229),
            .I(N__51166));
    InMux I__12288 (
            .O(N__51228),
            .I(N__51163));
    InMux I__12287 (
            .O(N__51227),
            .I(N__51156));
    InMux I__12286 (
            .O(N__51226),
            .I(N__51156));
    InMux I__12285 (
            .O(N__51225),
            .I(N__51156));
    LocalMux I__12284 (
            .O(N__51222),
            .I(N__51153));
    InMux I__12283 (
            .O(N__51221),
            .I(N__51150));
    InMux I__12282 (
            .O(N__51220),
            .I(N__51143));
    InMux I__12281 (
            .O(N__51219),
            .I(N__51143));
    InMux I__12280 (
            .O(N__51218),
            .I(N__51143));
    InMux I__12279 (
            .O(N__51217),
            .I(N__51134));
    InMux I__12278 (
            .O(N__51214),
            .I(N__51134));
    InMux I__12277 (
            .O(N__51211),
            .I(N__51134));
    InMux I__12276 (
            .O(N__51210),
            .I(N__51134));
    InMux I__12275 (
            .O(N__51209),
            .I(N__51129));
    InMux I__12274 (
            .O(N__51208),
            .I(N__51129));
    InMux I__12273 (
            .O(N__51207),
            .I(N__51126));
    InMux I__12272 (
            .O(N__51206),
            .I(N__51123));
    InMux I__12271 (
            .O(N__51205),
            .I(N__51118));
    InMux I__12270 (
            .O(N__51204),
            .I(N__51118));
    InMux I__12269 (
            .O(N__51201),
            .I(N__51115));
    InMux I__12268 (
            .O(N__51200),
            .I(N__51112));
    CascadeMux I__12267 (
            .O(N__51199),
            .I(N__51107));
    InMux I__12266 (
            .O(N__51198),
            .I(N__51101));
    InMux I__12265 (
            .O(N__51197),
            .I(N__51096));
    InMux I__12264 (
            .O(N__51196),
            .I(N__51096));
    Span4Mux_v I__12263 (
            .O(N__51193),
            .I(N__51087));
    Span4Mux_h I__12262 (
            .O(N__51186),
            .I(N__51087));
    LocalMux I__12261 (
            .O(N__51181),
            .I(N__51087));
    LocalMux I__12260 (
            .O(N__51178),
            .I(N__51087));
    LocalMux I__12259 (
            .O(N__51169),
            .I(N__51084));
    LocalMux I__12258 (
            .O(N__51166),
            .I(N__51075));
    LocalMux I__12257 (
            .O(N__51163),
            .I(N__51075));
    LocalMux I__12256 (
            .O(N__51156),
            .I(N__51075));
    Span4Mux_v I__12255 (
            .O(N__51153),
            .I(N__51075));
    LocalMux I__12254 (
            .O(N__51150),
            .I(N__51070));
    LocalMux I__12253 (
            .O(N__51143),
            .I(N__51063));
    LocalMux I__12252 (
            .O(N__51134),
            .I(N__51063));
    LocalMux I__12251 (
            .O(N__51129),
            .I(N__51063));
    LocalMux I__12250 (
            .O(N__51126),
            .I(N__51058));
    LocalMux I__12249 (
            .O(N__51123),
            .I(N__51049));
    LocalMux I__12248 (
            .O(N__51118),
            .I(N__51049));
    LocalMux I__12247 (
            .O(N__51115),
            .I(N__51049));
    LocalMux I__12246 (
            .O(N__51112),
            .I(N__51049));
    InMux I__12245 (
            .O(N__51111),
            .I(N__51044));
    InMux I__12244 (
            .O(N__51110),
            .I(N__51044));
    InMux I__12243 (
            .O(N__51107),
            .I(N__51041));
    InMux I__12242 (
            .O(N__51106),
            .I(N__51038));
    InMux I__12241 (
            .O(N__51105),
            .I(N__51033));
    InMux I__12240 (
            .O(N__51104),
            .I(N__51033));
    LocalMux I__12239 (
            .O(N__51101),
            .I(N__51022));
    LocalMux I__12238 (
            .O(N__51096),
            .I(N__51022));
    Span4Mux_v I__12237 (
            .O(N__51087),
            .I(N__51022));
    Span4Mux_v I__12236 (
            .O(N__51084),
            .I(N__51022));
    Span4Mux_v I__12235 (
            .O(N__51075),
            .I(N__51022));
    InMux I__12234 (
            .O(N__51074),
            .I(N__51017));
    InMux I__12233 (
            .O(N__51073),
            .I(N__51017));
    Span4Mux_v I__12232 (
            .O(N__51070),
            .I(N__51014));
    Span12Mux_h I__12231 (
            .O(N__51063),
            .I(N__51011));
    InMux I__12230 (
            .O(N__51062),
            .I(N__51006));
    InMux I__12229 (
            .O(N__51061),
            .I(N__51006));
    Span4Mux_h I__12228 (
            .O(N__51058),
            .I(N__51001));
    Span4Mux_v I__12227 (
            .O(N__51049),
            .I(N__51001));
    LocalMux I__12226 (
            .O(N__51044),
            .I(comm_state_2));
    LocalMux I__12225 (
            .O(N__51041),
            .I(comm_state_2));
    LocalMux I__12224 (
            .O(N__51038),
            .I(comm_state_2));
    LocalMux I__12223 (
            .O(N__51033),
            .I(comm_state_2));
    Odrv4 I__12222 (
            .O(N__51022),
            .I(comm_state_2));
    LocalMux I__12221 (
            .O(N__51017),
            .I(comm_state_2));
    Odrv4 I__12220 (
            .O(N__51014),
            .I(comm_state_2));
    Odrv12 I__12219 (
            .O(N__51011),
            .I(comm_state_2));
    LocalMux I__12218 (
            .O(N__51006),
            .I(comm_state_2));
    Odrv4 I__12217 (
            .O(N__51001),
            .I(comm_state_2));
    CascadeMux I__12216 (
            .O(N__50980),
            .I(N__50977));
    InMux I__12215 (
            .O(N__50977),
            .I(N__50974));
    LocalMux I__12214 (
            .O(N__50974),
            .I(N__50971));
    Span4Mux_h I__12213 (
            .O(N__50971),
            .I(N__50968));
    Odrv4 I__12212 (
            .O(N__50968),
            .I(n20734));
    CascadeMux I__12211 (
            .O(N__50965),
            .I(N__50957));
    InMux I__12210 (
            .O(N__50964),
            .I(N__50945));
    InMux I__12209 (
            .O(N__50963),
            .I(N__50938));
    InMux I__12208 (
            .O(N__50962),
            .I(N__50938));
    InMux I__12207 (
            .O(N__50961),
            .I(N__50938));
    InMux I__12206 (
            .O(N__50960),
            .I(N__50931));
    InMux I__12205 (
            .O(N__50957),
            .I(N__50922));
    InMux I__12204 (
            .O(N__50956),
            .I(N__50922));
    InMux I__12203 (
            .O(N__50955),
            .I(N__50922));
    InMux I__12202 (
            .O(N__50954),
            .I(N__50922));
    InMux I__12201 (
            .O(N__50953),
            .I(N__50916));
    CascadeMux I__12200 (
            .O(N__50952),
            .I(N__50903));
    InMux I__12199 (
            .O(N__50951),
            .I(N__50896));
    InMux I__12198 (
            .O(N__50950),
            .I(N__50896));
    InMux I__12197 (
            .O(N__50949),
            .I(N__50896));
    InMux I__12196 (
            .O(N__50948),
            .I(N__50893));
    LocalMux I__12195 (
            .O(N__50945),
            .I(N__50888));
    LocalMux I__12194 (
            .O(N__50938),
            .I(N__50888));
    CascadeMux I__12193 (
            .O(N__50937),
            .I(N__50885));
    InMux I__12192 (
            .O(N__50936),
            .I(N__50877));
    InMux I__12191 (
            .O(N__50935),
            .I(N__50872));
    InMux I__12190 (
            .O(N__50934),
            .I(N__50872));
    LocalMux I__12189 (
            .O(N__50931),
            .I(N__50867));
    LocalMux I__12188 (
            .O(N__50922),
            .I(N__50867));
    InMux I__12187 (
            .O(N__50921),
            .I(N__50860));
    InMux I__12186 (
            .O(N__50920),
            .I(N__50860));
    InMux I__12185 (
            .O(N__50919),
            .I(N__50860));
    LocalMux I__12184 (
            .O(N__50916),
            .I(N__50857));
    InMux I__12183 (
            .O(N__50915),
            .I(N__50852));
    InMux I__12182 (
            .O(N__50914),
            .I(N__50849));
    InMux I__12181 (
            .O(N__50913),
            .I(N__50844));
    InMux I__12180 (
            .O(N__50912),
            .I(N__50844));
    InMux I__12179 (
            .O(N__50911),
            .I(N__50841));
    CascadeMux I__12178 (
            .O(N__50910),
            .I(N__50838));
    CascadeMux I__12177 (
            .O(N__50909),
            .I(N__50831));
    InMux I__12176 (
            .O(N__50908),
            .I(N__50825));
    InMux I__12175 (
            .O(N__50907),
            .I(N__50825));
    InMux I__12174 (
            .O(N__50906),
            .I(N__50822));
    InMux I__12173 (
            .O(N__50903),
            .I(N__50818));
    LocalMux I__12172 (
            .O(N__50896),
            .I(N__50813));
    LocalMux I__12171 (
            .O(N__50893),
            .I(N__50813));
    Span4Mux_h I__12170 (
            .O(N__50888),
            .I(N__50810));
    InMux I__12169 (
            .O(N__50885),
            .I(N__50805));
    InMux I__12168 (
            .O(N__50884),
            .I(N__50805));
    InMux I__12167 (
            .O(N__50883),
            .I(N__50802));
    InMux I__12166 (
            .O(N__50882),
            .I(N__50798));
    InMux I__12165 (
            .O(N__50881),
            .I(N__50793));
    InMux I__12164 (
            .O(N__50880),
            .I(N__50793));
    LocalMux I__12163 (
            .O(N__50877),
            .I(N__50788));
    LocalMux I__12162 (
            .O(N__50872),
            .I(N__50788));
    Span4Mux_v I__12161 (
            .O(N__50867),
            .I(N__50781));
    LocalMux I__12160 (
            .O(N__50860),
            .I(N__50781));
    Span4Mux_v I__12159 (
            .O(N__50857),
            .I(N__50781));
    InMux I__12158 (
            .O(N__50856),
            .I(N__50776));
    InMux I__12157 (
            .O(N__50855),
            .I(N__50776));
    LocalMux I__12156 (
            .O(N__50852),
            .I(N__50771));
    LocalMux I__12155 (
            .O(N__50849),
            .I(N__50771));
    LocalMux I__12154 (
            .O(N__50844),
            .I(N__50766));
    LocalMux I__12153 (
            .O(N__50841),
            .I(N__50766));
    InMux I__12152 (
            .O(N__50838),
            .I(N__50763));
    CascadeMux I__12151 (
            .O(N__50837),
            .I(N__50760));
    CascadeMux I__12150 (
            .O(N__50836),
            .I(N__50756));
    CascadeMux I__12149 (
            .O(N__50835),
            .I(N__50753));
    CascadeMux I__12148 (
            .O(N__50834),
            .I(N__50750));
    InMux I__12147 (
            .O(N__50831),
            .I(N__50741));
    InMux I__12146 (
            .O(N__50830),
            .I(N__50741));
    LocalMux I__12145 (
            .O(N__50825),
            .I(N__50736));
    LocalMux I__12144 (
            .O(N__50822),
            .I(N__50736));
    InMux I__12143 (
            .O(N__50821),
            .I(N__50733));
    LocalMux I__12142 (
            .O(N__50818),
            .I(N__50730));
    Span4Mux_h I__12141 (
            .O(N__50813),
            .I(N__50725));
    Span4Mux_v I__12140 (
            .O(N__50810),
            .I(N__50725));
    LocalMux I__12139 (
            .O(N__50805),
            .I(N__50718));
    LocalMux I__12138 (
            .O(N__50802),
            .I(N__50718));
    InMux I__12137 (
            .O(N__50801),
            .I(N__50707));
    LocalMux I__12136 (
            .O(N__50798),
            .I(N__50704));
    LocalMux I__12135 (
            .O(N__50793),
            .I(N__50695));
    Span4Mux_v I__12134 (
            .O(N__50788),
            .I(N__50695));
    Span4Mux_h I__12133 (
            .O(N__50781),
            .I(N__50695));
    LocalMux I__12132 (
            .O(N__50776),
            .I(N__50695));
    Span4Mux_v I__12131 (
            .O(N__50771),
            .I(N__50692));
    Sp12to4 I__12130 (
            .O(N__50766),
            .I(N__50689));
    LocalMux I__12129 (
            .O(N__50763),
            .I(N__50686));
    InMux I__12128 (
            .O(N__50760),
            .I(N__50681));
    InMux I__12127 (
            .O(N__50759),
            .I(N__50681));
    InMux I__12126 (
            .O(N__50756),
            .I(N__50666));
    InMux I__12125 (
            .O(N__50753),
            .I(N__50666));
    InMux I__12124 (
            .O(N__50750),
            .I(N__50666));
    InMux I__12123 (
            .O(N__50749),
            .I(N__50666));
    InMux I__12122 (
            .O(N__50748),
            .I(N__50666));
    InMux I__12121 (
            .O(N__50747),
            .I(N__50666));
    InMux I__12120 (
            .O(N__50746),
            .I(N__50666));
    LocalMux I__12119 (
            .O(N__50741),
            .I(N__50663));
    Span4Mux_h I__12118 (
            .O(N__50736),
            .I(N__50660));
    LocalMux I__12117 (
            .O(N__50733),
            .I(N__50657));
    Span4Mux_v I__12116 (
            .O(N__50730),
            .I(N__50652));
    Span4Mux_h I__12115 (
            .O(N__50725),
            .I(N__50652));
    InMux I__12114 (
            .O(N__50724),
            .I(N__50642));
    InMux I__12113 (
            .O(N__50723),
            .I(N__50639));
    Span4Mux_h I__12112 (
            .O(N__50718),
            .I(N__50636));
    InMux I__12111 (
            .O(N__50717),
            .I(N__50619));
    InMux I__12110 (
            .O(N__50716),
            .I(N__50619));
    InMux I__12109 (
            .O(N__50715),
            .I(N__50619));
    InMux I__12108 (
            .O(N__50714),
            .I(N__50619));
    InMux I__12107 (
            .O(N__50713),
            .I(N__50619));
    InMux I__12106 (
            .O(N__50712),
            .I(N__50619));
    InMux I__12105 (
            .O(N__50711),
            .I(N__50619));
    InMux I__12104 (
            .O(N__50710),
            .I(N__50619));
    LocalMux I__12103 (
            .O(N__50707),
            .I(N__50614));
    Span4Mux_v I__12102 (
            .O(N__50704),
            .I(N__50614));
    Span4Mux_v I__12101 (
            .O(N__50695),
            .I(N__50611));
    Sp12to4 I__12100 (
            .O(N__50692),
            .I(N__50606));
    Span12Mux_v I__12099 (
            .O(N__50689),
            .I(N__50606));
    Span12Mux_s11_h I__12098 (
            .O(N__50686),
            .I(N__50603));
    LocalMux I__12097 (
            .O(N__50681),
            .I(N__50594));
    LocalMux I__12096 (
            .O(N__50666),
            .I(N__50594));
    Span4Mux_h I__12095 (
            .O(N__50663),
            .I(N__50594));
    Span4Mux_v I__12094 (
            .O(N__50660),
            .I(N__50594));
    Span4Mux_h I__12093 (
            .O(N__50657),
            .I(N__50589));
    Span4Mux_h I__12092 (
            .O(N__50652),
            .I(N__50589));
    InMux I__12091 (
            .O(N__50651),
            .I(N__50582));
    InMux I__12090 (
            .O(N__50650),
            .I(N__50582));
    InMux I__12089 (
            .O(N__50649),
            .I(N__50582));
    InMux I__12088 (
            .O(N__50648),
            .I(N__50573));
    InMux I__12087 (
            .O(N__50647),
            .I(N__50573));
    InMux I__12086 (
            .O(N__50646),
            .I(N__50573));
    InMux I__12085 (
            .O(N__50645),
            .I(N__50573));
    LocalMux I__12084 (
            .O(N__50642),
            .I(adc_state_0));
    LocalMux I__12083 (
            .O(N__50639),
            .I(adc_state_0));
    Odrv4 I__12082 (
            .O(N__50636),
            .I(adc_state_0));
    LocalMux I__12081 (
            .O(N__50619),
            .I(adc_state_0));
    Odrv4 I__12080 (
            .O(N__50614),
            .I(adc_state_0));
    Odrv4 I__12079 (
            .O(N__50611),
            .I(adc_state_0));
    Odrv12 I__12078 (
            .O(N__50606),
            .I(adc_state_0));
    Odrv12 I__12077 (
            .O(N__50603),
            .I(adc_state_0));
    Odrv4 I__12076 (
            .O(N__50594),
            .I(adc_state_0));
    Odrv4 I__12075 (
            .O(N__50589),
            .I(adc_state_0));
    LocalMux I__12074 (
            .O(N__50582),
            .I(adc_state_0));
    LocalMux I__12073 (
            .O(N__50573),
            .I(adc_state_0));
    CascadeMux I__12072 (
            .O(N__50548),
            .I(N__50544));
    CascadeMux I__12071 (
            .O(N__50547),
            .I(N__50541));
    InMux I__12070 (
            .O(N__50544),
            .I(N__50537));
    InMux I__12069 (
            .O(N__50541),
            .I(N__50532));
    InMux I__12068 (
            .O(N__50540),
            .I(N__50532));
    LocalMux I__12067 (
            .O(N__50537),
            .I(cmd_rdadctmp_12));
    LocalMux I__12066 (
            .O(N__50532),
            .I(cmd_rdadctmp_12));
    InMux I__12065 (
            .O(N__50527),
            .I(N__50523));
    InMux I__12064 (
            .O(N__50526),
            .I(N__50520));
    LocalMux I__12063 (
            .O(N__50523),
            .I(N__50507));
    LocalMux I__12062 (
            .O(N__50520),
            .I(N__50507));
    InMux I__12061 (
            .O(N__50519),
            .I(N__50502));
    InMux I__12060 (
            .O(N__50518),
            .I(N__50502));
    InMux I__12059 (
            .O(N__50517),
            .I(N__50497));
    InMux I__12058 (
            .O(N__50516),
            .I(N__50486));
    InMux I__12057 (
            .O(N__50515),
            .I(N__50486));
    InMux I__12056 (
            .O(N__50514),
            .I(N__50483));
    InMux I__12055 (
            .O(N__50513),
            .I(N__50480));
    InMux I__12054 (
            .O(N__50512),
            .I(N__50476));
    Span4Mux_v I__12053 (
            .O(N__50507),
            .I(N__50471));
    LocalMux I__12052 (
            .O(N__50502),
            .I(N__50471));
    InMux I__12051 (
            .O(N__50501),
            .I(N__50466));
    InMux I__12050 (
            .O(N__50500),
            .I(N__50463));
    LocalMux I__12049 (
            .O(N__50497),
            .I(N__50460));
    InMux I__12048 (
            .O(N__50496),
            .I(N__50448));
    InMux I__12047 (
            .O(N__50495),
            .I(N__50448));
    InMux I__12046 (
            .O(N__50494),
            .I(N__50443));
    InMux I__12045 (
            .O(N__50493),
            .I(N__50443));
    InMux I__12044 (
            .O(N__50492),
            .I(N__50438));
    InMux I__12043 (
            .O(N__50491),
            .I(N__50438));
    LocalMux I__12042 (
            .O(N__50486),
            .I(N__50431));
    LocalMux I__12041 (
            .O(N__50483),
            .I(N__50431));
    LocalMux I__12040 (
            .O(N__50480),
            .I(N__50431));
    InMux I__12039 (
            .O(N__50479),
            .I(N__50428));
    LocalMux I__12038 (
            .O(N__50476),
            .I(N__50425));
    Span4Mux_h I__12037 (
            .O(N__50471),
            .I(N__50422));
    CascadeMux I__12036 (
            .O(N__50470),
            .I(N__50419));
    InMux I__12035 (
            .O(N__50469),
            .I(N__50412));
    LocalMux I__12034 (
            .O(N__50466),
            .I(N__50409));
    LocalMux I__12033 (
            .O(N__50463),
            .I(N__50406));
    Span12Mux_v I__12032 (
            .O(N__50460),
            .I(N__50403));
    InMux I__12031 (
            .O(N__50459),
            .I(N__50390));
    InMux I__12030 (
            .O(N__50458),
            .I(N__50390));
    InMux I__12029 (
            .O(N__50457),
            .I(N__50390));
    InMux I__12028 (
            .O(N__50456),
            .I(N__50390));
    InMux I__12027 (
            .O(N__50455),
            .I(N__50390));
    InMux I__12026 (
            .O(N__50454),
            .I(N__50390));
    InMux I__12025 (
            .O(N__50453),
            .I(N__50387));
    LocalMux I__12024 (
            .O(N__50448),
            .I(N__50378));
    LocalMux I__12023 (
            .O(N__50443),
            .I(N__50378));
    LocalMux I__12022 (
            .O(N__50438),
            .I(N__50378));
    Span4Mux_v I__12021 (
            .O(N__50431),
            .I(N__50378));
    LocalMux I__12020 (
            .O(N__50428),
            .I(N__50373));
    Span4Mux_v I__12019 (
            .O(N__50425),
            .I(N__50373));
    Span4Mux_h I__12018 (
            .O(N__50422),
            .I(N__50370));
    InMux I__12017 (
            .O(N__50419),
            .I(N__50367));
    InMux I__12016 (
            .O(N__50418),
            .I(N__50358));
    InMux I__12015 (
            .O(N__50417),
            .I(N__50358));
    InMux I__12014 (
            .O(N__50416),
            .I(N__50358));
    InMux I__12013 (
            .O(N__50415),
            .I(N__50358));
    LocalMux I__12012 (
            .O(N__50412),
            .I(N__50353));
    Span4Mux_v I__12011 (
            .O(N__50409),
            .I(N__50353));
    Span4Mux_h I__12010 (
            .O(N__50406),
            .I(N__50350));
    Span12Mux_h I__12009 (
            .O(N__50403),
            .I(N__50347));
    LocalMux I__12008 (
            .O(N__50390),
            .I(N__50336));
    LocalMux I__12007 (
            .O(N__50387),
            .I(N__50336));
    Span4Mux_v I__12006 (
            .O(N__50378),
            .I(N__50336));
    Span4Mux_v I__12005 (
            .O(N__50373),
            .I(N__50336));
    Span4Mux_v I__12004 (
            .O(N__50370),
            .I(N__50336));
    LocalMux I__12003 (
            .O(N__50367),
            .I(n12542));
    LocalMux I__12002 (
            .O(N__50358),
            .I(n12542));
    Odrv4 I__12001 (
            .O(N__50353),
            .I(n12542));
    Odrv4 I__12000 (
            .O(N__50350),
            .I(n12542));
    Odrv12 I__11999 (
            .O(N__50347),
            .I(n12542));
    Odrv4 I__11998 (
            .O(N__50336),
            .I(n12542));
    CascadeMux I__11997 (
            .O(N__50323),
            .I(N__50319));
    CascadeMux I__11996 (
            .O(N__50322),
            .I(N__50316));
    InMux I__11995 (
            .O(N__50319),
            .I(N__50312));
    InMux I__11994 (
            .O(N__50316),
            .I(N__50309));
    InMux I__11993 (
            .O(N__50315),
            .I(N__50306));
    LocalMux I__11992 (
            .O(N__50312),
            .I(cmd_rdadctmp_13));
    LocalMux I__11991 (
            .O(N__50309),
            .I(cmd_rdadctmp_13));
    LocalMux I__11990 (
            .O(N__50306),
            .I(cmd_rdadctmp_13));
    InMux I__11989 (
            .O(N__50299),
            .I(N__50296));
    LocalMux I__11988 (
            .O(N__50296),
            .I(N__50293));
    Span4Mux_h I__11987 (
            .O(N__50293),
            .I(N__50289));
    InMux I__11986 (
            .O(N__50292),
            .I(N__50286));
    Span4Mux_h I__11985 (
            .O(N__50289),
            .I(N__50282));
    LocalMux I__11984 (
            .O(N__50286),
            .I(N__50279));
    InMux I__11983 (
            .O(N__50285),
            .I(N__50276));
    Span4Mux_v I__11982 (
            .O(N__50282),
            .I(N__50273));
    Odrv12 I__11981 (
            .O(N__50279),
            .I(buf_control_0));
    LocalMux I__11980 (
            .O(N__50276),
            .I(buf_control_0));
    Odrv4 I__11979 (
            .O(N__50273),
            .I(buf_control_0));
    InMux I__11978 (
            .O(N__50266),
            .I(N__50263));
    LocalMux I__11977 (
            .O(N__50263),
            .I(N__50260));
    Sp12to4 I__11976 (
            .O(N__50260),
            .I(N__50257));
    Span12Mux_v I__11975 (
            .O(N__50257),
            .I(N__50252));
    InMux I__11974 (
            .O(N__50256),
            .I(N__50249));
    InMux I__11973 (
            .O(N__50255),
            .I(N__50246));
    Odrv12 I__11972 (
            .O(N__50252),
            .I(wdtick_flag));
    LocalMux I__11971 (
            .O(N__50249),
            .I(wdtick_flag));
    LocalMux I__11970 (
            .O(N__50246),
            .I(wdtick_flag));
    IoInMux I__11969 (
            .O(N__50239),
            .I(N__50236));
    LocalMux I__11968 (
            .O(N__50236),
            .I(N__50233));
    Span4Mux_s1_v I__11967 (
            .O(N__50233),
            .I(N__50230));
    Span4Mux_v I__11966 (
            .O(N__50230),
            .I(N__50227));
    Span4Mux_v I__11965 (
            .O(N__50227),
            .I(N__50224));
    Odrv4 I__11964 (
            .O(N__50224),
            .I(CONT_SD));
    InMux I__11963 (
            .O(N__50221),
            .I(N__50217));
    InMux I__11962 (
            .O(N__50220),
            .I(N__50214));
    LocalMux I__11961 (
            .O(N__50217),
            .I(N__50211));
    LocalMux I__11960 (
            .O(N__50214),
            .I(N__50206));
    Span4Mux_v I__11959 (
            .O(N__50211),
            .I(N__50206));
    Span4Mux_h I__11958 (
            .O(N__50206),
            .I(N__50202));
    InMux I__11957 (
            .O(N__50205),
            .I(N__50199));
    Odrv4 I__11956 (
            .O(N__50202),
            .I(\comm_spi.n22647 ));
    LocalMux I__11955 (
            .O(N__50199),
            .I(\comm_spi.n22647 ));
    InMux I__11954 (
            .O(N__50194),
            .I(N__50191));
    LocalMux I__11953 (
            .O(N__50191),
            .I(N__50187));
    CascadeMux I__11952 (
            .O(N__50190),
            .I(N__50184));
    Span4Mux_v I__11951 (
            .O(N__50187),
            .I(N__50178));
    InMux I__11950 (
            .O(N__50184),
            .I(N__50175));
    InMux I__11949 (
            .O(N__50183),
            .I(N__50172));
    InMux I__11948 (
            .O(N__50182),
            .I(N__50169));
    InMux I__11947 (
            .O(N__50181),
            .I(N__50166));
    Span4Mux_v I__11946 (
            .O(N__50178),
            .I(N__50163));
    LocalMux I__11945 (
            .O(N__50175),
            .I(N__50158));
    LocalMux I__11944 (
            .O(N__50172),
            .I(N__50158));
    LocalMux I__11943 (
            .O(N__50169),
            .I(N__50155));
    LocalMux I__11942 (
            .O(N__50166),
            .I(N__50148));
    Span4Mux_h I__11941 (
            .O(N__50163),
            .I(N__50148));
    Span4Mux_v I__11940 (
            .O(N__50158),
            .I(N__50148));
    Span4Mux_h I__11939 (
            .O(N__50155),
            .I(N__50145));
    Span4Mux_h I__11938 (
            .O(N__50148),
            .I(N__50142));
    Odrv4 I__11937 (
            .O(N__50145),
            .I(comm_buf_1_5));
    Odrv4 I__11936 (
            .O(N__50142),
            .I(comm_buf_1_5));
    CascadeMux I__11935 (
            .O(N__50137),
            .I(N__50133));
    InMux I__11934 (
            .O(N__50136),
            .I(N__50129));
    InMux I__11933 (
            .O(N__50133),
            .I(N__50126));
    InMux I__11932 (
            .O(N__50132),
            .I(N__50123));
    LocalMux I__11931 (
            .O(N__50129),
            .I(N__50120));
    LocalMux I__11930 (
            .O(N__50126),
            .I(N__50115));
    LocalMux I__11929 (
            .O(N__50123),
            .I(N__50115));
    Span4Mux_v I__11928 (
            .O(N__50120),
            .I(N__50110));
    Span4Mux_h I__11927 (
            .O(N__50115),
            .I(N__50110));
    Span4Mux_h I__11926 (
            .O(N__50110),
            .I(N__50107));
    Span4Mux_h I__11925 (
            .O(N__50107),
            .I(N__50104));
    Odrv4 I__11924 (
            .O(N__50104),
            .I(n14_adj_1557));
    InMux I__11923 (
            .O(N__50101),
            .I(N__50089));
    InMux I__11922 (
            .O(N__50100),
            .I(N__50089));
    InMux I__11921 (
            .O(N__50099),
            .I(N__50082));
    InMux I__11920 (
            .O(N__50098),
            .I(N__50082));
    InMux I__11919 (
            .O(N__50097),
            .I(N__50079));
    InMux I__11918 (
            .O(N__50096),
            .I(N__50070));
    InMux I__11917 (
            .O(N__50095),
            .I(N__50070));
    CascadeMux I__11916 (
            .O(N__50094),
            .I(N__50064));
    LocalMux I__11915 (
            .O(N__50089),
            .I(N__50061));
    InMux I__11914 (
            .O(N__50088),
            .I(N__50058));
    InMux I__11913 (
            .O(N__50087),
            .I(N__50055));
    LocalMux I__11912 (
            .O(N__50082),
            .I(N__50050));
    LocalMux I__11911 (
            .O(N__50079),
            .I(N__50050));
    InMux I__11910 (
            .O(N__50078),
            .I(N__50047));
    InMux I__11909 (
            .O(N__50077),
            .I(N__50040));
    InMux I__11908 (
            .O(N__50076),
            .I(N__50040));
    InMux I__11907 (
            .O(N__50075),
            .I(N__50040));
    LocalMux I__11906 (
            .O(N__50070),
            .I(N__50037));
    InMux I__11905 (
            .O(N__50069),
            .I(N__50030));
    InMux I__11904 (
            .O(N__50068),
            .I(N__50030));
    InMux I__11903 (
            .O(N__50067),
            .I(N__50030));
    InMux I__11902 (
            .O(N__50064),
            .I(N__50027));
    Span4Mux_v I__11901 (
            .O(N__50061),
            .I(N__50016));
    LocalMux I__11900 (
            .O(N__50058),
            .I(N__50016));
    LocalMux I__11899 (
            .O(N__50055),
            .I(N__50016));
    Span4Mux_h I__11898 (
            .O(N__50050),
            .I(N__50016));
    LocalMux I__11897 (
            .O(N__50047),
            .I(N__50016));
    LocalMux I__11896 (
            .O(N__50040),
            .I(N__50011));
    Span4Mux_v I__11895 (
            .O(N__50037),
            .I(N__50011));
    LocalMux I__11894 (
            .O(N__50030),
            .I(N__50003));
    LocalMux I__11893 (
            .O(N__50027),
            .I(N__49999));
    Span4Mux_v I__11892 (
            .O(N__50016),
            .I(N__49994));
    Span4Mux_h I__11891 (
            .O(N__50011),
            .I(N__49994));
    InMux I__11890 (
            .O(N__50010),
            .I(N__49989));
    InMux I__11889 (
            .O(N__50009),
            .I(N__49989));
    InMux I__11888 (
            .O(N__50008),
            .I(N__49986));
    InMux I__11887 (
            .O(N__50007),
            .I(N__49981));
    InMux I__11886 (
            .O(N__50006),
            .I(N__49981));
    Span12Mux_v I__11885 (
            .O(N__50003),
            .I(N__49978));
    InMux I__11884 (
            .O(N__50002),
            .I(N__49975));
    Span4Mux_h I__11883 (
            .O(N__49999),
            .I(N__49968));
    Span4Mux_h I__11882 (
            .O(N__49994),
            .I(N__49968));
    LocalMux I__11881 (
            .O(N__49989),
            .I(N__49968));
    LocalMux I__11880 (
            .O(N__49986),
            .I(comm_index_2));
    LocalMux I__11879 (
            .O(N__49981),
            .I(comm_index_2));
    Odrv12 I__11878 (
            .O(N__49978),
            .I(comm_index_2));
    LocalMux I__11877 (
            .O(N__49975),
            .I(comm_index_2));
    Odrv4 I__11876 (
            .O(N__49968),
            .I(comm_index_2));
    CascadeMux I__11875 (
            .O(N__49957),
            .I(N__49954));
    InMux I__11874 (
            .O(N__49954),
            .I(N__49951));
    LocalMux I__11873 (
            .O(N__49951),
            .I(N__49948));
    Span4Mux_h I__11872 (
            .O(N__49948),
            .I(N__49944));
    InMux I__11871 (
            .O(N__49947),
            .I(N__49941));
    Span4Mux_h I__11870 (
            .O(N__49944),
            .I(N__49936));
    LocalMux I__11869 (
            .O(N__49941),
            .I(N__49933));
    InMux I__11868 (
            .O(N__49940),
            .I(N__49930));
    InMux I__11867 (
            .O(N__49939),
            .I(N__49927));
    Odrv4 I__11866 (
            .O(N__49936),
            .I(n18824));
    Odrv12 I__11865 (
            .O(N__49933),
            .I(n18824));
    LocalMux I__11864 (
            .O(N__49930),
            .I(n18824));
    LocalMux I__11863 (
            .O(N__49927),
            .I(n18824));
    CascadeMux I__11862 (
            .O(N__49918),
            .I(n20563_cascade_));
    InMux I__11861 (
            .O(N__49915),
            .I(N__49911));
    InMux I__11860 (
            .O(N__49914),
            .I(N__49905));
    LocalMux I__11859 (
            .O(N__49911),
            .I(N__49902));
    InMux I__11858 (
            .O(N__49910),
            .I(N__49897));
    InMux I__11857 (
            .O(N__49909),
            .I(N__49897));
    InMux I__11856 (
            .O(N__49908),
            .I(N__49894));
    LocalMux I__11855 (
            .O(N__49905),
            .I(N__49891));
    Span4Mux_h I__11854 (
            .O(N__49902),
            .I(N__49888));
    LocalMux I__11853 (
            .O(N__49897),
            .I(N__49883));
    LocalMux I__11852 (
            .O(N__49894),
            .I(N__49883));
    Span4Mux_h I__11851 (
            .O(N__49891),
            .I(N__49876));
    Span4Mux_h I__11850 (
            .O(N__49888),
            .I(N__49876));
    Span4Mux_v I__11849 (
            .O(N__49883),
            .I(N__49876));
    Odrv4 I__11848 (
            .O(N__49876),
            .I(n20627));
    CascadeMux I__11847 (
            .O(N__49873),
            .I(n12_adj_1539_cascade_));
    InMux I__11846 (
            .O(N__49870),
            .I(N__49864));
    InMux I__11845 (
            .O(N__49869),
            .I(N__49864));
    LocalMux I__11844 (
            .O(N__49864),
            .I(N__49861));
    Span4Mux_h I__11843 (
            .O(N__49861),
            .I(N__49855));
    InMux I__11842 (
            .O(N__49860),
            .I(N__49850));
    InMux I__11841 (
            .O(N__49859),
            .I(N__49850));
    InMux I__11840 (
            .O(N__49858),
            .I(N__49847));
    Span4Mux_h I__11839 (
            .O(N__49855),
            .I(N__49839));
    LocalMux I__11838 (
            .O(N__49850),
            .I(N__49839));
    LocalMux I__11837 (
            .O(N__49847),
            .I(N__49839));
    InMux I__11836 (
            .O(N__49846),
            .I(N__49836));
    Span4Mux_v I__11835 (
            .O(N__49839),
            .I(N__49831));
    LocalMux I__11834 (
            .O(N__49836),
            .I(N__49831));
    Span4Mux_h I__11833 (
            .O(N__49831),
            .I(N__49828));
    Odrv4 I__11832 (
            .O(N__49828),
            .I(n20556));
    CEMux I__11831 (
            .O(N__49825),
            .I(N__49822));
    LocalMux I__11830 (
            .O(N__49822),
            .I(N__49818));
    InMux I__11829 (
            .O(N__49821),
            .I(N__49815));
    Span4Mux_v I__11828 (
            .O(N__49818),
            .I(N__49812));
    LocalMux I__11827 (
            .O(N__49815),
            .I(N__49809));
    Span4Mux_h I__11826 (
            .O(N__49812),
            .I(N__49804));
    Span4Mux_h I__11825 (
            .O(N__49809),
            .I(N__49804));
    Odrv4 I__11824 (
            .O(N__49804),
            .I(n12164));
    InMux I__11823 (
            .O(N__49801),
            .I(N__49792));
    InMux I__11822 (
            .O(N__49800),
            .I(N__49783));
    InMux I__11821 (
            .O(N__49799),
            .I(N__49783));
    InMux I__11820 (
            .O(N__49798),
            .I(N__49783));
    CascadeMux I__11819 (
            .O(N__49797),
            .I(N__49778));
    CascadeMux I__11818 (
            .O(N__49796),
            .I(N__49775));
    CascadeMux I__11817 (
            .O(N__49795),
            .I(N__49771));
    LocalMux I__11816 (
            .O(N__49792),
            .I(N__49764));
    InMux I__11815 (
            .O(N__49791),
            .I(N__49759));
    InMux I__11814 (
            .O(N__49790),
            .I(N__49759));
    LocalMux I__11813 (
            .O(N__49783),
            .I(N__49756));
    CascadeMux I__11812 (
            .O(N__49782),
            .I(N__49752));
    InMux I__11811 (
            .O(N__49781),
            .I(N__49747));
    InMux I__11810 (
            .O(N__49778),
            .I(N__49744));
    InMux I__11809 (
            .O(N__49775),
            .I(N__49735));
    InMux I__11808 (
            .O(N__49774),
            .I(N__49735));
    InMux I__11807 (
            .O(N__49771),
            .I(N__49735));
    InMux I__11806 (
            .O(N__49770),
            .I(N__49735));
    InMux I__11805 (
            .O(N__49769),
            .I(N__49730));
    InMux I__11804 (
            .O(N__49768),
            .I(N__49730));
    InMux I__11803 (
            .O(N__49767),
            .I(N__49727));
    Span4Mux_v I__11802 (
            .O(N__49764),
            .I(N__49722));
    LocalMux I__11801 (
            .O(N__49759),
            .I(N__49722));
    Span4Mux_v I__11800 (
            .O(N__49756),
            .I(N__49719));
    InMux I__11799 (
            .O(N__49755),
            .I(N__49712));
    InMux I__11798 (
            .O(N__49752),
            .I(N__49712));
    InMux I__11797 (
            .O(N__49751),
            .I(N__49712));
    InMux I__11796 (
            .O(N__49750),
            .I(N__49709));
    LocalMux I__11795 (
            .O(N__49747),
            .I(N__49700));
    LocalMux I__11794 (
            .O(N__49744),
            .I(N__49700));
    LocalMux I__11793 (
            .O(N__49735),
            .I(N__49700));
    LocalMux I__11792 (
            .O(N__49730),
            .I(N__49700));
    LocalMux I__11791 (
            .O(N__49727),
            .I(N__49696));
    Span4Mux_v I__11790 (
            .O(N__49722),
            .I(N__49693));
    Span4Mux_h I__11789 (
            .O(N__49719),
            .I(N__49690));
    LocalMux I__11788 (
            .O(N__49712),
            .I(N__49683));
    LocalMux I__11787 (
            .O(N__49709),
            .I(N__49683));
    Span4Mux_v I__11786 (
            .O(N__49700),
            .I(N__49683));
    InMux I__11785 (
            .O(N__49699),
            .I(N__49680));
    Sp12to4 I__11784 (
            .O(N__49696),
            .I(N__49677));
    Sp12to4 I__11783 (
            .O(N__49693),
            .I(N__49674));
    Span4Mux_h I__11782 (
            .O(N__49690),
            .I(N__49671));
    Sp12to4 I__11781 (
            .O(N__49683),
            .I(N__49666));
    LocalMux I__11780 (
            .O(N__49680),
            .I(N__49666));
    Span12Mux_v I__11779 (
            .O(N__49677),
            .I(N__49661));
    Span12Mux_s10_h I__11778 (
            .O(N__49674),
            .I(N__49661));
    Sp12to4 I__11777 (
            .O(N__49671),
            .I(N__49656));
    Span12Mux_h I__11776 (
            .O(N__49666),
            .I(N__49656));
    Span12Mux_v I__11775 (
            .O(N__49661),
            .I(N__49653));
    Span12Mux_v I__11774 (
            .O(N__49656),
            .I(N__49650));
    Odrv12 I__11773 (
            .O(N__49653),
            .I(ICE_SPI_CE0));
    Odrv12 I__11772 (
            .O(N__49650),
            .I(ICE_SPI_CE0));
    InMux I__11771 (
            .O(N__49645),
            .I(N__49642));
    LocalMux I__11770 (
            .O(N__49642),
            .I(N__49636));
    InMux I__11769 (
            .O(N__49641),
            .I(N__49629));
    InMux I__11768 (
            .O(N__49640),
            .I(N__49619));
    InMux I__11767 (
            .O(N__49639),
            .I(N__49619));
    Span4Mux_v I__11766 (
            .O(N__49636),
            .I(N__49616));
    InMux I__11765 (
            .O(N__49635),
            .I(N__49613));
    InMux I__11764 (
            .O(N__49634),
            .I(N__49610));
    InMux I__11763 (
            .O(N__49633),
            .I(N__49605));
    InMux I__11762 (
            .O(N__49632),
            .I(N__49605));
    LocalMux I__11761 (
            .O(N__49629),
            .I(N__49602));
    InMux I__11760 (
            .O(N__49628),
            .I(N__49593));
    InMux I__11759 (
            .O(N__49627),
            .I(N__49593));
    InMux I__11758 (
            .O(N__49626),
            .I(N__49593));
    InMux I__11757 (
            .O(N__49625),
            .I(N__49593));
    InMux I__11756 (
            .O(N__49624),
            .I(N__49590));
    LocalMux I__11755 (
            .O(N__49619),
            .I(comm_data_vld));
    Odrv4 I__11754 (
            .O(N__49616),
            .I(comm_data_vld));
    LocalMux I__11753 (
            .O(N__49613),
            .I(comm_data_vld));
    LocalMux I__11752 (
            .O(N__49610),
            .I(comm_data_vld));
    LocalMux I__11751 (
            .O(N__49605),
            .I(comm_data_vld));
    Odrv4 I__11750 (
            .O(N__49602),
            .I(comm_data_vld));
    LocalMux I__11749 (
            .O(N__49593),
            .I(comm_data_vld));
    LocalMux I__11748 (
            .O(N__49590),
            .I(comm_data_vld));
    InMux I__11747 (
            .O(N__49573),
            .I(N__49570));
    LocalMux I__11746 (
            .O(N__49570),
            .I(N__49567));
    Span4Mux_h I__11745 (
            .O(N__49567),
            .I(N__49564));
    Span4Mux_v I__11744 (
            .O(N__49564),
            .I(N__49561));
    Odrv4 I__11743 (
            .O(N__49561),
            .I(n23_adj_1574));
    CascadeMux I__11742 (
            .O(N__49558),
            .I(n21_adj_1573_cascade_));
    CEMux I__11741 (
            .O(N__49555),
            .I(N__49552));
    LocalMux I__11740 (
            .O(N__49552),
            .I(N__49549));
    Span4Mux_h I__11739 (
            .O(N__49549),
            .I(N__49546));
    Odrv4 I__11738 (
            .O(N__49546),
            .I(n18));
    CascadeMux I__11737 (
            .O(N__49543),
            .I(N__49540));
    InMux I__11736 (
            .O(N__49540),
            .I(N__49526));
    InMux I__11735 (
            .O(N__49539),
            .I(N__49515));
    InMux I__11734 (
            .O(N__49538),
            .I(N__49515));
    InMux I__11733 (
            .O(N__49537),
            .I(N__49506));
    InMux I__11732 (
            .O(N__49536),
            .I(N__49506));
    InMux I__11731 (
            .O(N__49535),
            .I(N__49506));
    InMux I__11730 (
            .O(N__49534),
            .I(N__49503));
    InMux I__11729 (
            .O(N__49533),
            .I(N__49500));
    InMux I__11728 (
            .O(N__49532),
            .I(N__49493));
    InMux I__11727 (
            .O(N__49531),
            .I(N__49493));
    InMux I__11726 (
            .O(N__49530),
            .I(N__49493));
    InMux I__11725 (
            .O(N__49529),
            .I(N__49489));
    LocalMux I__11724 (
            .O(N__49526),
            .I(N__49486));
    InMux I__11723 (
            .O(N__49525),
            .I(N__49481));
    InMux I__11722 (
            .O(N__49524),
            .I(N__49481));
    InMux I__11721 (
            .O(N__49523),
            .I(N__49476));
    InMux I__11720 (
            .O(N__49522),
            .I(N__49476));
    InMux I__11719 (
            .O(N__49521),
            .I(N__49471));
    InMux I__11718 (
            .O(N__49520),
            .I(N__49471));
    LocalMux I__11717 (
            .O(N__49515),
            .I(N__49468));
    CascadeMux I__11716 (
            .O(N__49514),
            .I(N__49464));
    CascadeMux I__11715 (
            .O(N__49513),
            .I(N__49459));
    LocalMux I__11714 (
            .O(N__49506),
            .I(N__49456));
    LocalMux I__11713 (
            .O(N__49503),
            .I(N__49451));
    LocalMux I__11712 (
            .O(N__49500),
            .I(N__49451));
    LocalMux I__11711 (
            .O(N__49493),
            .I(N__49448));
    InMux I__11710 (
            .O(N__49492),
            .I(N__49445));
    LocalMux I__11709 (
            .O(N__49489),
            .I(N__49442));
    Span4Mux_v I__11708 (
            .O(N__49486),
            .I(N__49435));
    LocalMux I__11707 (
            .O(N__49481),
            .I(N__49435));
    LocalMux I__11706 (
            .O(N__49476),
            .I(N__49435));
    LocalMux I__11705 (
            .O(N__49471),
            .I(N__49430));
    Span4Mux_h I__11704 (
            .O(N__49468),
            .I(N__49430));
    InMux I__11703 (
            .O(N__49467),
            .I(N__49426));
    InMux I__11702 (
            .O(N__49464),
            .I(N__49423));
    InMux I__11701 (
            .O(N__49463),
            .I(N__49420));
    InMux I__11700 (
            .O(N__49462),
            .I(N__49417));
    InMux I__11699 (
            .O(N__49459),
            .I(N__49414));
    Span4Mux_v I__11698 (
            .O(N__49456),
            .I(N__49407));
    Span4Mux_v I__11697 (
            .O(N__49451),
            .I(N__49407));
    Span4Mux_v I__11696 (
            .O(N__49448),
            .I(N__49407));
    LocalMux I__11695 (
            .O(N__49445),
            .I(N__49404));
    Span4Mux_v I__11694 (
            .O(N__49442),
            .I(N__49397));
    Span4Mux_v I__11693 (
            .O(N__49435),
            .I(N__49397));
    Span4Mux_h I__11692 (
            .O(N__49430),
            .I(N__49397));
    CascadeMux I__11691 (
            .O(N__49429),
            .I(N__49392));
    LocalMux I__11690 (
            .O(N__49426),
            .I(N__49387));
    LocalMux I__11689 (
            .O(N__49423),
            .I(N__49387));
    LocalMux I__11688 (
            .O(N__49420),
            .I(N__49384));
    LocalMux I__11687 (
            .O(N__49417),
            .I(N__49375));
    LocalMux I__11686 (
            .O(N__49414),
            .I(N__49375));
    Span4Mux_h I__11685 (
            .O(N__49407),
            .I(N__49375));
    Span4Mux_v I__11684 (
            .O(N__49404),
            .I(N__49375));
    Span4Mux_h I__11683 (
            .O(N__49397),
            .I(N__49372));
    InMux I__11682 (
            .O(N__49396),
            .I(N__49367));
    InMux I__11681 (
            .O(N__49395),
            .I(N__49367));
    InMux I__11680 (
            .O(N__49392),
            .I(N__49364));
    Span4Mux_h I__11679 (
            .O(N__49387),
            .I(N__49361));
    Odrv4 I__11678 (
            .O(N__49384),
            .I(comm_index_1));
    Odrv4 I__11677 (
            .O(N__49375),
            .I(comm_index_1));
    Odrv4 I__11676 (
            .O(N__49372),
            .I(comm_index_1));
    LocalMux I__11675 (
            .O(N__49367),
            .I(comm_index_1));
    LocalMux I__11674 (
            .O(N__49364),
            .I(comm_index_1));
    Odrv4 I__11673 (
            .O(N__49361),
            .I(comm_index_1));
    CascadeMux I__11672 (
            .O(N__49348),
            .I(N__49345));
    InMux I__11671 (
            .O(N__49345),
            .I(N__49341));
    InMux I__11670 (
            .O(N__49344),
            .I(N__49338));
    LocalMux I__11669 (
            .O(N__49341),
            .I(N__49335));
    LocalMux I__11668 (
            .O(N__49338),
            .I(N__49332));
    Span4Mux_v I__11667 (
            .O(N__49335),
            .I(N__49327));
    Span4Mux_h I__11666 (
            .O(N__49332),
            .I(N__49327));
    Odrv4 I__11665 (
            .O(N__49327),
            .I(comm_length_1));
    InMux I__11664 (
            .O(N__49324),
            .I(N__49320));
    InMux I__11663 (
            .O(N__49323),
            .I(N__49317));
    LocalMux I__11662 (
            .O(N__49320),
            .I(N__49314));
    LocalMux I__11661 (
            .O(N__49317),
            .I(N__49311));
    Span4Mux_v I__11660 (
            .O(N__49314),
            .I(N__49306));
    Span4Mux_h I__11659 (
            .O(N__49311),
            .I(N__49306));
    Odrv4 I__11658 (
            .O(N__49306),
            .I(n4_adj_1576));
    InMux I__11657 (
            .O(N__49303),
            .I(N__49299));
    InMux I__11656 (
            .O(N__49302),
            .I(N__49295));
    LocalMux I__11655 (
            .O(N__49299),
            .I(N__49292));
    InMux I__11654 (
            .O(N__49298),
            .I(N__49289));
    LocalMux I__11653 (
            .O(N__49295),
            .I(N__49281));
    Span4Mux_v I__11652 (
            .O(N__49292),
            .I(N__49281));
    LocalMux I__11651 (
            .O(N__49289),
            .I(N__49281));
    InMux I__11650 (
            .O(N__49288),
            .I(N__49278));
    Span4Mux_h I__11649 (
            .O(N__49281),
            .I(N__49275));
    LocalMux I__11648 (
            .O(N__49278),
            .I(comm_cmd_7));
    Odrv4 I__11647 (
            .O(N__49275),
            .I(comm_cmd_7));
    CascadeMux I__11646 (
            .O(N__49270),
            .I(n5_cascade_));
    IoInMux I__11645 (
            .O(N__49267),
            .I(N__49264));
    LocalMux I__11644 (
            .O(N__49264),
            .I(N__49261));
    Span4Mux_s1_h I__11643 (
            .O(N__49261),
            .I(N__49258));
    Sp12to4 I__11642 (
            .O(N__49258),
            .I(N__49255));
    Span12Mux_v I__11641 (
            .O(N__49255),
            .I(N__49252));
    Odrv12 I__11640 (
            .O(N__49252),
            .I(ICE_GPMI_0));
    CEMux I__11639 (
            .O(N__49249),
            .I(N__49246));
    LocalMux I__11638 (
            .O(N__49246),
            .I(N__49243));
    Odrv4 I__11637 (
            .O(N__49243),
            .I(n11406));
    InMux I__11636 (
            .O(N__49240),
            .I(N__49232));
    InMux I__11635 (
            .O(N__49239),
            .I(N__49229));
    InMux I__11634 (
            .O(N__49238),
            .I(N__49226));
    InMux I__11633 (
            .O(N__49237),
            .I(N__49223));
    InMux I__11632 (
            .O(N__49236),
            .I(N__49220));
    CascadeMux I__11631 (
            .O(N__49235),
            .I(N__49217));
    LocalMux I__11630 (
            .O(N__49232),
            .I(N__49212));
    LocalMux I__11629 (
            .O(N__49229),
            .I(N__49207));
    LocalMux I__11628 (
            .O(N__49226),
            .I(N__49200));
    LocalMux I__11627 (
            .O(N__49223),
            .I(N__49200));
    LocalMux I__11626 (
            .O(N__49220),
            .I(N__49200));
    InMux I__11625 (
            .O(N__49217),
            .I(N__49193));
    InMux I__11624 (
            .O(N__49216),
            .I(N__49193));
    InMux I__11623 (
            .O(N__49215),
            .I(N__49193));
    Span4Mux_h I__11622 (
            .O(N__49212),
            .I(N__49190));
    InMux I__11621 (
            .O(N__49211),
            .I(N__49187));
    InMux I__11620 (
            .O(N__49210),
            .I(N__49182));
    Sp12to4 I__11619 (
            .O(N__49207),
            .I(N__49179));
    Span4Mux_v I__11618 (
            .O(N__49200),
            .I(N__49176));
    LocalMux I__11617 (
            .O(N__49193),
            .I(N__49169));
    Span4Mux_v I__11616 (
            .O(N__49190),
            .I(N__49169));
    LocalMux I__11615 (
            .O(N__49187),
            .I(N__49169));
    InMux I__11614 (
            .O(N__49186),
            .I(N__49164));
    InMux I__11613 (
            .O(N__49185),
            .I(N__49164));
    LocalMux I__11612 (
            .O(N__49182),
            .I(N__49159));
    Span12Mux_v I__11611 (
            .O(N__49179),
            .I(N__49159));
    Span4Mux_h I__11610 (
            .O(N__49176),
            .I(N__49154));
    Span4Mux_v I__11609 (
            .O(N__49169),
            .I(N__49154));
    LocalMux I__11608 (
            .O(N__49164),
            .I(n12220));
    Odrv12 I__11607 (
            .O(N__49159),
            .I(n12220));
    Odrv4 I__11606 (
            .O(N__49154),
            .I(n12220));
    CascadeMux I__11605 (
            .O(N__49147),
            .I(n10_adj_1572_cascade_));
    CascadeMux I__11604 (
            .O(N__49144),
            .I(N__49141));
    InMux I__11603 (
            .O(N__49141),
            .I(N__49135));
    InMux I__11602 (
            .O(N__49140),
            .I(N__49135));
    LocalMux I__11601 (
            .O(N__49135),
            .I(N__49132));
    Span4Mux_h I__11600 (
            .O(N__49132),
            .I(N__49129));
    Odrv4 I__11599 (
            .O(N__49129),
            .I(n20643));
    InMux I__11598 (
            .O(N__49126),
            .I(N__49123));
    LocalMux I__11597 (
            .O(N__49123),
            .I(n4_adj_1596));
    InMux I__11596 (
            .O(N__49120),
            .I(N__49117));
    LocalMux I__11595 (
            .O(N__49117),
            .I(N__49114));
    Span4Mux_h I__11594 (
            .O(N__49114),
            .I(N__49110));
    InMux I__11593 (
            .O(N__49113),
            .I(N__49107));
    Odrv4 I__11592 (
            .O(N__49110),
            .I(n2342));
    LocalMux I__11591 (
            .O(N__49107),
            .I(n2342));
    CEMux I__11590 (
            .O(N__49102),
            .I(N__49099));
    LocalMux I__11589 (
            .O(N__49099),
            .I(N__49096));
    Odrv12 I__11588 (
            .O(N__49096),
            .I(n11836));
    SRMux I__11587 (
            .O(N__49093),
            .I(N__49090));
    LocalMux I__11586 (
            .O(N__49090),
            .I(N__49087));
    Span4Mux_h I__11585 (
            .O(N__49087),
            .I(N__49084));
    Span4Mux_h I__11584 (
            .O(N__49084),
            .I(N__49081));
    Odrv4 I__11583 (
            .O(N__49081),
            .I(n14722));
    InMux I__11582 (
            .O(N__49078),
            .I(N__49074));
    InMux I__11581 (
            .O(N__49077),
            .I(N__49071));
    LocalMux I__11580 (
            .O(N__49074),
            .I(N__49067));
    LocalMux I__11579 (
            .O(N__49071),
            .I(N__49064));
    InMux I__11578 (
            .O(N__49070),
            .I(N__49061));
    Span4Mux_h I__11577 (
            .O(N__49067),
            .I(N__49058));
    Span4Mux_h I__11576 (
            .O(N__49064),
            .I(N__49055));
    LocalMux I__11575 (
            .O(N__49061),
            .I(buf_adcdata_iac_5));
    Odrv4 I__11574 (
            .O(N__49058),
            .I(buf_adcdata_iac_5));
    Odrv4 I__11573 (
            .O(N__49055),
            .I(buf_adcdata_iac_5));
    CascadeMux I__11572 (
            .O(N__49048),
            .I(N__49045));
    InMux I__11571 (
            .O(N__49045),
            .I(N__49042));
    LocalMux I__11570 (
            .O(N__49042),
            .I(N__49038));
    CascadeMux I__11569 (
            .O(N__49041),
            .I(N__49035));
    Span4Mux_v I__11568 (
            .O(N__49038),
            .I(N__49032));
    InMux I__11567 (
            .O(N__49035),
            .I(N__49029));
    Sp12to4 I__11566 (
            .O(N__49032),
            .I(N__49026));
    LocalMux I__11565 (
            .O(N__49029),
            .I(N__49022));
    Span12Mux_h I__11564 (
            .O(N__49026),
            .I(N__49019));
    InMux I__11563 (
            .O(N__49025),
            .I(N__49016));
    Odrv4 I__11562 (
            .O(N__49022),
            .I(cmd_rdadctmp_11));
    Odrv12 I__11561 (
            .O(N__49019),
            .I(cmd_rdadctmp_11));
    LocalMux I__11560 (
            .O(N__49016),
            .I(cmd_rdadctmp_11));
    InMux I__11559 (
            .O(N__49009),
            .I(N__49005));
    InMux I__11558 (
            .O(N__49008),
            .I(N__49001));
    LocalMux I__11557 (
            .O(N__49005),
            .I(N__48994));
    InMux I__11556 (
            .O(N__49004),
            .I(N__48991));
    LocalMux I__11555 (
            .O(N__49001),
            .I(N__48987));
    InMux I__11554 (
            .O(N__49000),
            .I(N__48984));
    InMux I__11553 (
            .O(N__48999),
            .I(N__48979));
    InMux I__11552 (
            .O(N__48998),
            .I(N__48979));
    InMux I__11551 (
            .O(N__48997),
            .I(N__48976));
    Span4Mux_v I__11550 (
            .O(N__48994),
            .I(N__48970));
    LocalMux I__11549 (
            .O(N__48991),
            .I(N__48970));
    InMux I__11548 (
            .O(N__48990),
            .I(N__48963));
    Span4Mux_h I__11547 (
            .O(N__48987),
            .I(N__48954));
    LocalMux I__11546 (
            .O(N__48984),
            .I(N__48954));
    LocalMux I__11545 (
            .O(N__48979),
            .I(N__48948));
    LocalMux I__11544 (
            .O(N__48976),
            .I(N__48948));
    InMux I__11543 (
            .O(N__48975),
            .I(N__48945));
    Span4Mux_h I__11542 (
            .O(N__48970),
            .I(N__48942));
    InMux I__11541 (
            .O(N__48969),
            .I(N__48939));
    InMux I__11540 (
            .O(N__48968),
            .I(N__48936));
    InMux I__11539 (
            .O(N__48967),
            .I(N__48931));
    InMux I__11538 (
            .O(N__48966),
            .I(N__48931));
    LocalMux I__11537 (
            .O(N__48963),
            .I(N__48928));
    InMux I__11536 (
            .O(N__48962),
            .I(N__48923));
    InMux I__11535 (
            .O(N__48961),
            .I(N__48923));
    InMux I__11534 (
            .O(N__48960),
            .I(N__48918));
    InMux I__11533 (
            .O(N__48959),
            .I(N__48918));
    Span4Mux_v I__11532 (
            .O(N__48954),
            .I(N__48915));
    InMux I__11531 (
            .O(N__48953),
            .I(N__48912));
    Span4Mux_h I__11530 (
            .O(N__48948),
            .I(N__48905));
    LocalMux I__11529 (
            .O(N__48945),
            .I(N__48905));
    Span4Mux_h I__11528 (
            .O(N__48942),
            .I(N__48898));
    LocalMux I__11527 (
            .O(N__48939),
            .I(N__48898));
    LocalMux I__11526 (
            .O(N__48936),
            .I(N__48898));
    LocalMux I__11525 (
            .O(N__48931),
            .I(N__48895));
    Span4Mux_v I__11524 (
            .O(N__48928),
            .I(N__48887));
    LocalMux I__11523 (
            .O(N__48923),
            .I(N__48887));
    LocalMux I__11522 (
            .O(N__48918),
            .I(N__48884));
    Span4Mux_h I__11521 (
            .O(N__48915),
            .I(N__48879));
    LocalMux I__11520 (
            .O(N__48912),
            .I(N__48879));
    InMux I__11519 (
            .O(N__48911),
            .I(N__48874));
    InMux I__11518 (
            .O(N__48910),
            .I(N__48874));
    Span4Mux_v I__11517 (
            .O(N__48905),
            .I(N__48870));
    Span4Mux_h I__11516 (
            .O(N__48898),
            .I(N__48867));
    Span4Mux_h I__11515 (
            .O(N__48895),
            .I(N__48864));
    InMux I__11514 (
            .O(N__48894),
            .I(N__48859));
    InMux I__11513 (
            .O(N__48893),
            .I(N__48859));
    InMux I__11512 (
            .O(N__48892),
            .I(N__48856));
    Span4Mux_v I__11511 (
            .O(N__48887),
            .I(N__48847));
    Span4Mux_v I__11510 (
            .O(N__48884),
            .I(N__48847));
    Span4Mux_h I__11509 (
            .O(N__48879),
            .I(N__48847));
    LocalMux I__11508 (
            .O(N__48874),
            .I(N__48847));
    InMux I__11507 (
            .O(N__48873),
            .I(N__48844));
    Odrv4 I__11506 (
            .O(N__48870),
            .I(n20543));
    Odrv4 I__11505 (
            .O(N__48867),
            .I(n20543));
    Odrv4 I__11504 (
            .O(N__48864),
            .I(n20543));
    LocalMux I__11503 (
            .O(N__48859),
            .I(n20543));
    LocalMux I__11502 (
            .O(N__48856),
            .I(n20543));
    Odrv4 I__11501 (
            .O(N__48847),
            .I(n20543));
    LocalMux I__11500 (
            .O(N__48844),
            .I(n20543));
    InMux I__11499 (
            .O(N__48829),
            .I(N__48825));
    InMux I__11498 (
            .O(N__48828),
            .I(N__48822));
    LocalMux I__11497 (
            .O(N__48825),
            .I(N__48818));
    LocalMux I__11496 (
            .O(N__48822),
            .I(N__48815));
    InMux I__11495 (
            .O(N__48821),
            .I(N__48812));
    Span4Mux_h I__11494 (
            .O(N__48818),
            .I(N__48809));
    Span4Mux_h I__11493 (
            .O(N__48815),
            .I(N__48806));
    LocalMux I__11492 (
            .O(N__48812),
            .I(buf_adcdata_iac_4));
    Odrv4 I__11491 (
            .O(N__48809),
            .I(buf_adcdata_iac_4));
    Odrv4 I__11490 (
            .O(N__48806),
            .I(buf_adcdata_iac_4));
    CascadeMux I__11489 (
            .O(N__48799),
            .I(N__48795));
    InMux I__11488 (
            .O(N__48798),
            .I(N__48792));
    InMux I__11487 (
            .O(N__48795),
            .I(N__48789));
    LocalMux I__11486 (
            .O(N__48792),
            .I(N__48786));
    LocalMux I__11485 (
            .O(N__48789),
            .I(N__48782));
    Span4Mux_v I__11484 (
            .O(N__48786),
            .I(N__48779));
    InMux I__11483 (
            .O(N__48785),
            .I(N__48776));
    Odrv12 I__11482 (
            .O(N__48782),
            .I(cmd_rdadctmp_14));
    Odrv4 I__11481 (
            .O(N__48779),
            .I(cmd_rdadctmp_14));
    LocalMux I__11480 (
            .O(N__48776),
            .I(cmd_rdadctmp_14));
    InMux I__11479 (
            .O(N__48769),
            .I(N__48766));
    LocalMux I__11478 (
            .O(N__48766),
            .I(N__48763));
    Odrv4 I__11477 (
            .O(N__48763),
            .I(\comm_spi.n14581 ));
    SRMux I__11476 (
            .O(N__48760),
            .I(N__48757));
    LocalMux I__11475 (
            .O(N__48757),
            .I(N__48754));
    Span4Mux_h I__11474 (
            .O(N__48754),
            .I(N__48751));
    Odrv4 I__11473 (
            .O(N__48751),
            .I(\comm_spi.iclk_N_754 ));
    InMux I__11472 (
            .O(N__48748),
            .I(N__48745));
    LocalMux I__11471 (
            .O(N__48745),
            .I(N__48741));
    InMux I__11470 (
            .O(N__48744),
            .I(N__48738));
    Span4Mux_v I__11469 (
            .O(N__48741),
            .I(N__48734));
    LocalMux I__11468 (
            .O(N__48738),
            .I(N__48731));
    InMux I__11467 (
            .O(N__48737),
            .I(N__48728));
    Sp12to4 I__11466 (
            .O(N__48734),
            .I(N__48725));
    Span4Mux_h I__11465 (
            .O(N__48731),
            .I(N__48720));
    LocalMux I__11464 (
            .O(N__48728),
            .I(N__48720));
    Span12Mux_h I__11463 (
            .O(N__48725),
            .I(N__48717));
    Span4Mux_v I__11462 (
            .O(N__48720),
            .I(N__48714));
    Odrv12 I__11461 (
            .O(N__48717),
            .I(comm_tx_buf_5));
    Odrv4 I__11460 (
            .O(N__48714),
            .I(comm_tx_buf_5));
    SRMux I__11459 (
            .O(N__48709),
            .I(N__48706));
    LocalMux I__11458 (
            .O(N__48706),
            .I(N__48703));
    Odrv12 I__11457 (
            .O(N__48703),
            .I(\comm_spi.data_tx_7__N_760 ));
    InMux I__11456 (
            .O(N__48700),
            .I(N__48696));
    InMux I__11455 (
            .O(N__48699),
            .I(N__48693));
    LocalMux I__11454 (
            .O(N__48696),
            .I(data_cntvec_14));
    LocalMux I__11453 (
            .O(N__48693),
            .I(data_cntvec_14));
    InMux I__11452 (
            .O(N__48688),
            .I(n19309));
    InMux I__11451 (
            .O(N__48685),
            .I(n19310));
    InMux I__11450 (
            .O(N__48682),
            .I(N__48678));
    InMux I__11449 (
            .O(N__48681),
            .I(N__48675));
    LocalMux I__11448 (
            .O(N__48678),
            .I(N__48672));
    LocalMux I__11447 (
            .O(N__48675),
            .I(data_cntvec_15));
    Odrv4 I__11446 (
            .O(N__48672),
            .I(data_cntvec_15));
    CEMux I__11445 (
            .O(N__48667),
            .I(N__48664));
    LocalMux I__11444 (
            .O(N__48664),
            .I(N__48659));
    CEMux I__11443 (
            .O(N__48663),
            .I(N__48656));
    CEMux I__11442 (
            .O(N__48662),
            .I(N__48652));
    Span4Mux_h I__11441 (
            .O(N__48659),
            .I(N__48649));
    LocalMux I__11440 (
            .O(N__48656),
            .I(N__48646));
    CEMux I__11439 (
            .O(N__48655),
            .I(N__48643));
    LocalMux I__11438 (
            .O(N__48652),
            .I(N__48640));
    Span4Mux_v I__11437 (
            .O(N__48649),
            .I(N__48635));
    Span4Mux_v I__11436 (
            .O(N__48646),
            .I(N__48635));
    LocalMux I__11435 (
            .O(N__48643),
            .I(N__48632));
    Span4Mux_h I__11434 (
            .O(N__48640),
            .I(N__48628));
    Span4Mux_h I__11433 (
            .O(N__48635),
            .I(N__48623));
    Span4Mux_h I__11432 (
            .O(N__48632),
            .I(N__48623));
    InMux I__11431 (
            .O(N__48631),
            .I(N__48620));
    Span4Mux_h I__11430 (
            .O(N__48628),
            .I(N__48617));
    Span4Mux_h I__11429 (
            .O(N__48623),
            .I(N__48614));
    LocalMux I__11428 (
            .O(N__48620),
            .I(N__48611));
    Odrv4 I__11427 (
            .O(N__48617),
            .I(n13443));
    Odrv4 I__11426 (
            .O(N__48614),
            .I(n13443));
    Odrv12 I__11425 (
            .O(N__48611),
            .I(n13443));
    SRMux I__11424 (
            .O(N__48604),
            .I(N__48600));
    SRMux I__11423 (
            .O(N__48603),
            .I(N__48597));
    LocalMux I__11422 (
            .O(N__48600),
            .I(N__48593));
    LocalMux I__11421 (
            .O(N__48597),
            .I(N__48590));
    SRMux I__11420 (
            .O(N__48596),
            .I(N__48587));
    Span4Mux_h I__11419 (
            .O(N__48593),
            .I(N__48583));
    Span4Mux_v I__11418 (
            .O(N__48590),
            .I(N__48580));
    LocalMux I__11417 (
            .O(N__48587),
            .I(N__48577));
    SRMux I__11416 (
            .O(N__48586),
            .I(N__48574));
    Odrv4 I__11415 (
            .O(N__48583),
            .I(n14632));
    Odrv4 I__11414 (
            .O(N__48580),
            .I(n14632));
    Odrv12 I__11413 (
            .O(N__48577),
            .I(n14632));
    LocalMux I__11412 (
            .O(N__48574),
            .I(n14632));
    InMux I__11411 (
            .O(N__48565),
            .I(N__48561));
    InMux I__11410 (
            .O(N__48564),
            .I(N__48558));
    LocalMux I__11409 (
            .O(N__48561),
            .I(N__48554));
    LocalMux I__11408 (
            .O(N__48558),
            .I(N__48551));
    InMux I__11407 (
            .O(N__48557),
            .I(N__48548));
    Span4Mux_v I__11406 (
            .O(N__48554),
            .I(N__48545));
    Span4Mux_h I__11405 (
            .O(N__48551),
            .I(N__48542));
    LocalMux I__11404 (
            .O(N__48548),
            .I(buf_adcdata_iac_6));
    Odrv4 I__11403 (
            .O(N__48545),
            .I(buf_adcdata_iac_6));
    Odrv4 I__11402 (
            .O(N__48542),
            .I(buf_adcdata_iac_6));
    InMux I__11401 (
            .O(N__48535),
            .I(N__48530));
    InMux I__11400 (
            .O(N__48534),
            .I(N__48527));
    CascadeMux I__11399 (
            .O(N__48533),
            .I(N__48521));
    LocalMux I__11398 (
            .O(N__48530),
            .I(N__48518));
    LocalMux I__11397 (
            .O(N__48527),
            .I(N__48515));
    InMux I__11396 (
            .O(N__48526),
            .I(N__48512));
    InMux I__11395 (
            .O(N__48525),
            .I(N__48499));
    InMux I__11394 (
            .O(N__48524),
            .I(N__48499));
    InMux I__11393 (
            .O(N__48521),
            .I(N__48496));
    Span4Mux_h I__11392 (
            .O(N__48518),
            .I(N__48489));
    Span4Mux_h I__11391 (
            .O(N__48515),
            .I(N__48484));
    LocalMux I__11390 (
            .O(N__48512),
            .I(N__48484));
    CascadeMux I__11389 (
            .O(N__48511),
            .I(N__48481));
    InMux I__11388 (
            .O(N__48510),
            .I(N__48469));
    InMux I__11387 (
            .O(N__48509),
            .I(N__48469));
    InMux I__11386 (
            .O(N__48508),
            .I(N__48469));
    InMux I__11385 (
            .O(N__48507),
            .I(N__48469));
    InMux I__11384 (
            .O(N__48506),
            .I(N__48464));
    InMux I__11383 (
            .O(N__48505),
            .I(N__48464));
    InMux I__11382 (
            .O(N__48504),
            .I(N__48461));
    LocalMux I__11381 (
            .O(N__48499),
            .I(N__48456));
    LocalMux I__11380 (
            .O(N__48496),
            .I(N__48456));
    InMux I__11379 (
            .O(N__48495),
            .I(N__48453));
    InMux I__11378 (
            .O(N__48494),
            .I(N__48448));
    InMux I__11377 (
            .O(N__48493),
            .I(N__48448));
    InMux I__11376 (
            .O(N__48492),
            .I(N__48445));
    Span4Mux_h I__11375 (
            .O(N__48489),
            .I(N__48440));
    Span4Mux_h I__11374 (
            .O(N__48484),
            .I(N__48440));
    InMux I__11373 (
            .O(N__48481),
            .I(N__48432));
    InMux I__11372 (
            .O(N__48480),
            .I(N__48432));
    InMux I__11371 (
            .O(N__48479),
            .I(N__48427));
    InMux I__11370 (
            .O(N__48478),
            .I(N__48427));
    LocalMux I__11369 (
            .O(N__48469),
            .I(N__48422));
    LocalMux I__11368 (
            .O(N__48464),
            .I(N__48422));
    LocalMux I__11367 (
            .O(N__48461),
            .I(N__48419));
    Span4Mux_h I__11366 (
            .O(N__48456),
            .I(N__48416));
    LocalMux I__11365 (
            .O(N__48453),
            .I(N__48413));
    LocalMux I__11364 (
            .O(N__48448),
            .I(N__48408));
    LocalMux I__11363 (
            .O(N__48445),
            .I(N__48408));
    Span4Mux_h I__11362 (
            .O(N__48440),
            .I(N__48405));
    InMux I__11361 (
            .O(N__48439),
            .I(N__48402));
    InMux I__11360 (
            .O(N__48438),
            .I(N__48399));
    InMux I__11359 (
            .O(N__48437),
            .I(N__48396));
    LocalMux I__11358 (
            .O(N__48432),
            .I(N__48389));
    LocalMux I__11357 (
            .O(N__48427),
            .I(N__48389));
    Span4Mux_h I__11356 (
            .O(N__48422),
            .I(N__48389));
    Span12Mux_h I__11355 (
            .O(N__48419),
            .I(N__48386));
    Span4Mux_v I__11354 (
            .O(N__48416),
            .I(N__48383));
    Span4Mux_v I__11353 (
            .O(N__48413),
            .I(N__48378));
    Span4Mux_h I__11352 (
            .O(N__48408),
            .I(N__48378));
    Span4Mux_h I__11351 (
            .O(N__48405),
            .I(N__48375));
    LocalMux I__11350 (
            .O(N__48402),
            .I(n20540));
    LocalMux I__11349 (
            .O(N__48399),
            .I(n20540));
    LocalMux I__11348 (
            .O(N__48396),
            .I(n20540));
    Odrv4 I__11347 (
            .O(N__48389),
            .I(n20540));
    Odrv12 I__11346 (
            .O(N__48386),
            .I(n20540));
    Odrv4 I__11345 (
            .O(N__48383),
            .I(n20540));
    Odrv4 I__11344 (
            .O(N__48378),
            .I(n20540));
    Odrv4 I__11343 (
            .O(N__48375),
            .I(n20540));
    CascadeMux I__11342 (
            .O(N__48358),
            .I(N__48355));
    InMux I__11341 (
            .O(N__48355),
            .I(N__48352));
    LocalMux I__11340 (
            .O(N__48352),
            .I(N__48343));
    InMux I__11339 (
            .O(N__48351),
            .I(N__48336));
    InMux I__11338 (
            .O(N__48350),
            .I(N__48336));
    InMux I__11337 (
            .O(N__48349),
            .I(N__48336));
    InMux I__11336 (
            .O(N__48348),
            .I(N__48332));
    InMux I__11335 (
            .O(N__48347),
            .I(N__48329));
    CascadeMux I__11334 (
            .O(N__48346),
            .I(N__48326));
    Span4Mux_h I__11333 (
            .O(N__48343),
            .I(N__48316));
    LocalMux I__11332 (
            .O(N__48336),
            .I(N__48311));
    CascadeMux I__11331 (
            .O(N__48335),
            .I(N__48308));
    LocalMux I__11330 (
            .O(N__48332),
            .I(N__48305));
    LocalMux I__11329 (
            .O(N__48329),
            .I(N__48302));
    InMux I__11328 (
            .O(N__48326),
            .I(N__48293));
    InMux I__11327 (
            .O(N__48325),
            .I(N__48293));
    InMux I__11326 (
            .O(N__48324),
            .I(N__48293));
    InMux I__11325 (
            .O(N__48323),
            .I(N__48293));
    InMux I__11324 (
            .O(N__48322),
            .I(N__48288));
    InMux I__11323 (
            .O(N__48321),
            .I(N__48288));
    InMux I__11322 (
            .O(N__48320),
            .I(N__48275));
    InMux I__11321 (
            .O(N__48319),
            .I(N__48275));
    Span4Mux_h I__11320 (
            .O(N__48316),
            .I(N__48272));
    InMux I__11319 (
            .O(N__48315),
            .I(N__48269));
    InMux I__11318 (
            .O(N__48314),
            .I(N__48266));
    Span4Mux_v I__11317 (
            .O(N__48311),
            .I(N__48259));
    InMux I__11316 (
            .O(N__48308),
            .I(N__48256));
    Span4Mux_v I__11315 (
            .O(N__48305),
            .I(N__48251));
    Span4Mux_v I__11314 (
            .O(N__48302),
            .I(N__48251));
    LocalMux I__11313 (
            .O(N__48293),
            .I(N__48248));
    LocalMux I__11312 (
            .O(N__48288),
            .I(N__48245));
    InMux I__11311 (
            .O(N__48287),
            .I(N__48242));
    InMux I__11310 (
            .O(N__48286),
            .I(N__48235));
    InMux I__11309 (
            .O(N__48285),
            .I(N__48235));
    InMux I__11308 (
            .O(N__48284),
            .I(N__48235));
    CascadeMux I__11307 (
            .O(N__48283),
            .I(N__48232));
    CascadeMux I__11306 (
            .O(N__48282),
            .I(N__48229));
    CascadeMux I__11305 (
            .O(N__48281),
            .I(N__48226));
    CascadeMux I__11304 (
            .O(N__48280),
            .I(N__48220));
    LocalMux I__11303 (
            .O(N__48275),
            .I(N__48209));
    Span4Mux_v I__11302 (
            .O(N__48272),
            .I(N__48209));
    LocalMux I__11301 (
            .O(N__48269),
            .I(N__48209));
    LocalMux I__11300 (
            .O(N__48266),
            .I(N__48206));
    CascadeMux I__11299 (
            .O(N__48265),
            .I(N__48199));
    CascadeMux I__11298 (
            .O(N__48264),
            .I(N__48191));
    CascadeMux I__11297 (
            .O(N__48263),
            .I(N__48188));
    CascadeMux I__11296 (
            .O(N__48262),
            .I(N__48185));
    Span4Mux_h I__11295 (
            .O(N__48259),
            .I(N__48166));
    LocalMux I__11294 (
            .O(N__48256),
            .I(N__48166));
    Span4Mux_h I__11293 (
            .O(N__48251),
            .I(N__48166));
    Span4Mux_h I__11292 (
            .O(N__48248),
            .I(N__48157));
    Span4Mux_h I__11291 (
            .O(N__48245),
            .I(N__48157));
    LocalMux I__11290 (
            .O(N__48242),
            .I(N__48157));
    LocalMux I__11289 (
            .O(N__48235),
            .I(N__48157));
    InMux I__11288 (
            .O(N__48232),
            .I(N__48144));
    InMux I__11287 (
            .O(N__48229),
            .I(N__48144));
    InMux I__11286 (
            .O(N__48226),
            .I(N__48144));
    InMux I__11285 (
            .O(N__48225),
            .I(N__48144));
    InMux I__11284 (
            .O(N__48224),
            .I(N__48144));
    InMux I__11283 (
            .O(N__48223),
            .I(N__48144));
    InMux I__11282 (
            .O(N__48220),
            .I(N__48139));
    InMux I__11281 (
            .O(N__48219),
            .I(N__48139));
    InMux I__11280 (
            .O(N__48218),
            .I(N__48136));
    InMux I__11279 (
            .O(N__48217),
            .I(N__48131));
    InMux I__11278 (
            .O(N__48216),
            .I(N__48131));
    Span4Mux_h I__11277 (
            .O(N__48209),
            .I(N__48128));
    Span4Mux_h I__11276 (
            .O(N__48206),
            .I(N__48125));
    InMux I__11275 (
            .O(N__48205),
            .I(N__48118));
    InMux I__11274 (
            .O(N__48204),
            .I(N__48118));
    InMux I__11273 (
            .O(N__48203),
            .I(N__48118));
    CascadeMux I__11272 (
            .O(N__48202),
            .I(N__48114));
    InMux I__11271 (
            .O(N__48199),
            .I(N__48109));
    InMux I__11270 (
            .O(N__48198),
            .I(N__48098));
    InMux I__11269 (
            .O(N__48197),
            .I(N__48098));
    InMux I__11268 (
            .O(N__48196),
            .I(N__48098));
    InMux I__11267 (
            .O(N__48195),
            .I(N__48098));
    InMux I__11266 (
            .O(N__48194),
            .I(N__48098));
    InMux I__11265 (
            .O(N__48191),
            .I(N__48081));
    InMux I__11264 (
            .O(N__48188),
            .I(N__48081));
    InMux I__11263 (
            .O(N__48185),
            .I(N__48081));
    InMux I__11262 (
            .O(N__48184),
            .I(N__48081));
    InMux I__11261 (
            .O(N__48183),
            .I(N__48081));
    InMux I__11260 (
            .O(N__48182),
            .I(N__48081));
    InMux I__11259 (
            .O(N__48181),
            .I(N__48081));
    InMux I__11258 (
            .O(N__48180),
            .I(N__48081));
    InMux I__11257 (
            .O(N__48179),
            .I(N__48076));
    InMux I__11256 (
            .O(N__48178),
            .I(N__48076));
    InMux I__11255 (
            .O(N__48177),
            .I(N__48065));
    InMux I__11254 (
            .O(N__48176),
            .I(N__48065));
    InMux I__11253 (
            .O(N__48175),
            .I(N__48065));
    InMux I__11252 (
            .O(N__48174),
            .I(N__48065));
    InMux I__11251 (
            .O(N__48173),
            .I(N__48065));
    Span4Mux_h I__11250 (
            .O(N__48166),
            .I(N__48060));
    Span4Mux_v I__11249 (
            .O(N__48157),
            .I(N__48060));
    LocalMux I__11248 (
            .O(N__48144),
            .I(N__48051));
    LocalMux I__11247 (
            .O(N__48139),
            .I(N__48051));
    LocalMux I__11246 (
            .O(N__48136),
            .I(N__48051));
    LocalMux I__11245 (
            .O(N__48131),
            .I(N__48051));
    Span4Mux_v I__11244 (
            .O(N__48128),
            .I(N__48048));
    Span4Mux_h I__11243 (
            .O(N__48125),
            .I(N__48043));
    LocalMux I__11242 (
            .O(N__48118),
            .I(N__48043));
    InMux I__11241 (
            .O(N__48117),
            .I(N__48032));
    InMux I__11240 (
            .O(N__48114),
            .I(N__48025));
    InMux I__11239 (
            .O(N__48113),
            .I(N__48025));
    InMux I__11238 (
            .O(N__48112),
            .I(N__48025));
    LocalMux I__11237 (
            .O(N__48109),
            .I(N__48018));
    LocalMux I__11236 (
            .O(N__48098),
            .I(N__48018));
    LocalMux I__11235 (
            .O(N__48081),
            .I(N__48018));
    LocalMux I__11234 (
            .O(N__48076),
            .I(N__48013));
    LocalMux I__11233 (
            .O(N__48065),
            .I(N__48013));
    Sp12to4 I__11232 (
            .O(N__48060),
            .I(N__48010));
    Span4Mux_v I__11231 (
            .O(N__48051),
            .I(N__48003));
    Span4Mux_h I__11230 (
            .O(N__48048),
            .I(N__48003));
    Span4Mux_h I__11229 (
            .O(N__48043),
            .I(N__48003));
    InMux I__11228 (
            .O(N__48042),
            .I(N__47994));
    InMux I__11227 (
            .O(N__48041),
            .I(N__47994));
    InMux I__11226 (
            .O(N__48040),
            .I(N__47994));
    InMux I__11225 (
            .O(N__48039),
            .I(N__47994));
    InMux I__11224 (
            .O(N__48038),
            .I(N__47985));
    InMux I__11223 (
            .O(N__48037),
            .I(N__47985));
    InMux I__11222 (
            .O(N__48036),
            .I(N__47985));
    InMux I__11221 (
            .O(N__48035),
            .I(N__47985));
    LocalMux I__11220 (
            .O(N__48032),
            .I(adc_state_0_adj_1411));
    LocalMux I__11219 (
            .O(N__48025),
            .I(adc_state_0_adj_1411));
    Odrv4 I__11218 (
            .O(N__48018),
            .I(adc_state_0_adj_1411));
    Odrv12 I__11217 (
            .O(N__48013),
            .I(adc_state_0_adj_1411));
    Odrv12 I__11216 (
            .O(N__48010),
            .I(adc_state_0_adj_1411));
    Odrv4 I__11215 (
            .O(N__48003),
            .I(adc_state_0_adj_1411));
    LocalMux I__11214 (
            .O(N__47994),
            .I(adc_state_0_adj_1411));
    LocalMux I__11213 (
            .O(N__47985),
            .I(adc_state_0_adj_1411));
    CascadeMux I__11212 (
            .O(N__47968),
            .I(N__47964));
    InMux I__11211 (
            .O(N__47967),
            .I(N__47961));
    InMux I__11210 (
            .O(N__47964),
            .I(N__47958));
    LocalMux I__11209 (
            .O(N__47961),
            .I(N__47955));
    LocalMux I__11208 (
            .O(N__47958),
            .I(N__47952));
    Span4Mux_v I__11207 (
            .O(N__47955),
            .I(N__47949));
    Span12Mux_v I__11206 (
            .O(N__47952),
            .I(N__47945));
    Span4Mux_h I__11205 (
            .O(N__47949),
            .I(N__47942));
    InMux I__11204 (
            .O(N__47948),
            .I(N__47939));
    Odrv12 I__11203 (
            .O(N__47945),
            .I(cmd_rdadctmp_12_adj_1431));
    Odrv4 I__11202 (
            .O(N__47942),
            .I(cmd_rdadctmp_12_adj_1431));
    LocalMux I__11201 (
            .O(N__47939),
            .I(cmd_rdadctmp_12_adj_1431));
    InMux I__11200 (
            .O(N__47932),
            .I(N__47929));
    LocalMux I__11199 (
            .O(N__47929),
            .I(N__47925));
    InMux I__11198 (
            .O(N__47928),
            .I(N__47921));
    Span4Mux_v I__11197 (
            .O(N__47925),
            .I(N__47918));
    InMux I__11196 (
            .O(N__47924),
            .I(N__47915));
    LocalMux I__11195 (
            .O(N__47921),
            .I(buf_adcdata_vac_7));
    Odrv4 I__11194 (
            .O(N__47918),
            .I(buf_adcdata_vac_7));
    LocalMux I__11193 (
            .O(N__47915),
            .I(buf_adcdata_vac_7));
    InMux I__11192 (
            .O(N__47908),
            .I(N__47905));
    LocalMux I__11191 (
            .O(N__47905),
            .I(N__47902));
    Span4Mux_v I__11190 (
            .O(N__47902),
            .I(N__47899));
    Span4Mux_v I__11189 (
            .O(N__47899),
            .I(N__47895));
    CascadeMux I__11188 (
            .O(N__47898),
            .I(N__47892));
    Sp12to4 I__11187 (
            .O(N__47895),
            .I(N__47889));
    InMux I__11186 (
            .O(N__47892),
            .I(N__47886));
    Odrv12 I__11185 (
            .O(N__47889),
            .I(buf_adcdata_vdc_7));
    LocalMux I__11184 (
            .O(N__47886),
            .I(buf_adcdata_vdc_7));
    InMux I__11183 (
            .O(N__47881),
            .I(N__47877));
    CascadeMux I__11182 (
            .O(N__47880),
            .I(N__47874));
    LocalMux I__11181 (
            .O(N__47877),
            .I(N__47870));
    InMux I__11180 (
            .O(N__47874),
            .I(N__47867));
    InMux I__11179 (
            .O(N__47873),
            .I(N__47864));
    Span4Mux_h I__11178 (
            .O(N__47870),
            .I(N__47861));
    LocalMux I__11177 (
            .O(N__47867),
            .I(buf_adcdata_iac_7));
    LocalMux I__11176 (
            .O(N__47864),
            .I(buf_adcdata_iac_7));
    Odrv4 I__11175 (
            .O(N__47861),
            .I(buf_adcdata_iac_7));
    CascadeMux I__11174 (
            .O(N__47854),
            .I(n19_adj_1589_cascade_));
    InMux I__11173 (
            .O(N__47851),
            .I(N__47840));
    InMux I__11172 (
            .O(N__47850),
            .I(N__47837));
    CascadeMux I__11171 (
            .O(N__47849),
            .I(N__47826));
    InMux I__11170 (
            .O(N__47848),
            .I(N__47817));
    InMux I__11169 (
            .O(N__47847),
            .I(N__47814));
    InMux I__11168 (
            .O(N__47846),
            .I(N__47811));
    InMux I__11167 (
            .O(N__47845),
            .I(N__47806));
    InMux I__11166 (
            .O(N__47844),
            .I(N__47806));
    InMux I__11165 (
            .O(N__47843),
            .I(N__47803));
    LocalMux I__11164 (
            .O(N__47840),
            .I(N__47800));
    LocalMux I__11163 (
            .O(N__47837),
            .I(N__47797));
    InMux I__11162 (
            .O(N__47836),
            .I(N__47794));
    InMux I__11161 (
            .O(N__47835),
            .I(N__47791));
    InMux I__11160 (
            .O(N__47834),
            .I(N__47775));
    InMux I__11159 (
            .O(N__47833),
            .I(N__47771));
    InMux I__11158 (
            .O(N__47832),
            .I(N__47768));
    InMux I__11157 (
            .O(N__47831),
            .I(N__47763));
    InMux I__11156 (
            .O(N__47830),
            .I(N__47763));
    InMux I__11155 (
            .O(N__47829),
            .I(N__47758));
    InMux I__11154 (
            .O(N__47826),
            .I(N__47758));
    InMux I__11153 (
            .O(N__47825),
            .I(N__47755));
    InMux I__11152 (
            .O(N__47824),
            .I(N__47749));
    InMux I__11151 (
            .O(N__47823),
            .I(N__47738));
    InMux I__11150 (
            .O(N__47822),
            .I(N__47734));
    InMux I__11149 (
            .O(N__47821),
            .I(N__47731));
    InMux I__11148 (
            .O(N__47820),
            .I(N__47728));
    LocalMux I__11147 (
            .O(N__47817),
            .I(N__47721));
    LocalMux I__11146 (
            .O(N__47814),
            .I(N__47721));
    LocalMux I__11145 (
            .O(N__47811),
            .I(N__47718));
    LocalMux I__11144 (
            .O(N__47806),
            .I(N__47705));
    LocalMux I__11143 (
            .O(N__47803),
            .I(N__47705));
    Span4Mux_v I__11142 (
            .O(N__47800),
            .I(N__47705));
    Span4Mux_h I__11141 (
            .O(N__47797),
            .I(N__47705));
    LocalMux I__11140 (
            .O(N__47794),
            .I(N__47705));
    LocalMux I__11139 (
            .O(N__47791),
            .I(N__47705));
    InMux I__11138 (
            .O(N__47790),
            .I(N__47702));
    InMux I__11137 (
            .O(N__47789),
            .I(N__47691));
    InMux I__11136 (
            .O(N__47788),
            .I(N__47688));
    InMux I__11135 (
            .O(N__47787),
            .I(N__47683));
    InMux I__11134 (
            .O(N__47786),
            .I(N__47683));
    InMux I__11133 (
            .O(N__47785),
            .I(N__47674));
    InMux I__11132 (
            .O(N__47784),
            .I(N__47674));
    InMux I__11131 (
            .O(N__47783),
            .I(N__47674));
    InMux I__11130 (
            .O(N__47782),
            .I(N__47674));
    InMux I__11129 (
            .O(N__47781),
            .I(N__47665));
    InMux I__11128 (
            .O(N__47780),
            .I(N__47665));
    InMux I__11127 (
            .O(N__47779),
            .I(N__47665));
    InMux I__11126 (
            .O(N__47778),
            .I(N__47665));
    LocalMux I__11125 (
            .O(N__47775),
            .I(N__47662));
    InMux I__11124 (
            .O(N__47774),
            .I(N__47659));
    LocalMux I__11123 (
            .O(N__47771),
            .I(N__47654));
    LocalMux I__11122 (
            .O(N__47768),
            .I(N__47654));
    LocalMux I__11121 (
            .O(N__47763),
            .I(N__47649));
    LocalMux I__11120 (
            .O(N__47758),
            .I(N__47649));
    LocalMux I__11119 (
            .O(N__47755),
            .I(N__47646));
    InMux I__11118 (
            .O(N__47754),
            .I(N__47643));
    InMux I__11117 (
            .O(N__47753),
            .I(N__47640));
    InMux I__11116 (
            .O(N__47752),
            .I(N__47637));
    LocalMux I__11115 (
            .O(N__47749),
            .I(N__47634));
    InMux I__11114 (
            .O(N__47748),
            .I(N__47631));
    InMux I__11113 (
            .O(N__47747),
            .I(N__47628));
    InMux I__11112 (
            .O(N__47746),
            .I(N__47623));
    InMux I__11111 (
            .O(N__47745),
            .I(N__47623));
    InMux I__11110 (
            .O(N__47744),
            .I(N__47618));
    InMux I__11109 (
            .O(N__47743),
            .I(N__47618));
    InMux I__11108 (
            .O(N__47742),
            .I(N__47615));
    InMux I__11107 (
            .O(N__47741),
            .I(N__47612));
    LocalMux I__11106 (
            .O(N__47738),
            .I(N__47609));
    InMux I__11105 (
            .O(N__47737),
            .I(N__47606));
    LocalMux I__11104 (
            .O(N__47734),
            .I(N__47601));
    LocalMux I__11103 (
            .O(N__47731),
            .I(N__47601));
    LocalMux I__11102 (
            .O(N__47728),
            .I(N__47598));
    InMux I__11101 (
            .O(N__47727),
            .I(N__47593));
    InMux I__11100 (
            .O(N__47726),
            .I(N__47593));
    Span4Mux_v I__11099 (
            .O(N__47721),
            .I(N__47584));
    Span4Mux_v I__11098 (
            .O(N__47718),
            .I(N__47584));
    Span4Mux_v I__11097 (
            .O(N__47705),
            .I(N__47584));
    LocalMux I__11096 (
            .O(N__47702),
            .I(N__47584));
    CascadeMux I__11095 (
            .O(N__47701),
            .I(N__47581));
    InMux I__11094 (
            .O(N__47700),
            .I(N__47573));
    InMux I__11093 (
            .O(N__47699),
            .I(N__47573));
    InMux I__11092 (
            .O(N__47698),
            .I(N__47568));
    InMux I__11091 (
            .O(N__47697),
            .I(N__47568));
    InMux I__11090 (
            .O(N__47696),
            .I(N__47565));
    InMux I__11089 (
            .O(N__47695),
            .I(N__47562));
    InMux I__11088 (
            .O(N__47694),
            .I(N__47559));
    LocalMux I__11087 (
            .O(N__47691),
            .I(N__47556));
    LocalMux I__11086 (
            .O(N__47688),
            .I(N__47545));
    LocalMux I__11085 (
            .O(N__47683),
            .I(N__47545));
    LocalMux I__11084 (
            .O(N__47674),
            .I(N__47545));
    LocalMux I__11083 (
            .O(N__47665),
            .I(N__47545));
    Span4Mux_v I__11082 (
            .O(N__47662),
            .I(N__47545));
    LocalMux I__11081 (
            .O(N__47659),
            .I(N__47542));
    Span4Mux_v I__11080 (
            .O(N__47654),
            .I(N__47533));
    Span4Mux_v I__11079 (
            .O(N__47649),
            .I(N__47533));
    Span4Mux_v I__11078 (
            .O(N__47646),
            .I(N__47533));
    LocalMux I__11077 (
            .O(N__47643),
            .I(N__47533));
    LocalMux I__11076 (
            .O(N__47640),
            .I(N__47520));
    LocalMux I__11075 (
            .O(N__47637),
            .I(N__47520));
    Span4Mux_v I__11074 (
            .O(N__47634),
            .I(N__47520));
    LocalMux I__11073 (
            .O(N__47631),
            .I(N__47520));
    LocalMux I__11072 (
            .O(N__47628),
            .I(N__47520));
    LocalMux I__11071 (
            .O(N__47623),
            .I(N__47520));
    LocalMux I__11070 (
            .O(N__47618),
            .I(N__47509));
    LocalMux I__11069 (
            .O(N__47615),
            .I(N__47509));
    LocalMux I__11068 (
            .O(N__47612),
            .I(N__47509));
    Span4Mux_v I__11067 (
            .O(N__47609),
            .I(N__47509));
    LocalMux I__11066 (
            .O(N__47606),
            .I(N__47509));
    Span4Mux_v I__11065 (
            .O(N__47601),
            .I(N__47503));
    Span4Mux_v I__11064 (
            .O(N__47598),
            .I(N__47503));
    LocalMux I__11063 (
            .O(N__47593),
            .I(N__47498));
    Span4Mux_h I__11062 (
            .O(N__47584),
            .I(N__47498));
    InMux I__11061 (
            .O(N__47581),
            .I(N__47495));
    InMux I__11060 (
            .O(N__47580),
            .I(N__47488));
    InMux I__11059 (
            .O(N__47579),
            .I(N__47488));
    InMux I__11058 (
            .O(N__47578),
            .I(N__47488));
    LocalMux I__11057 (
            .O(N__47573),
            .I(N__47479));
    LocalMux I__11056 (
            .O(N__47568),
            .I(N__47479));
    LocalMux I__11055 (
            .O(N__47565),
            .I(N__47479));
    LocalMux I__11054 (
            .O(N__47562),
            .I(N__47479));
    LocalMux I__11053 (
            .O(N__47559),
            .I(N__47464));
    Span4Mux_v I__11052 (
            .O(N__47556),
            .I(N__47464));
    Span4Mux_v I__11051 (
            .O(N__47545),
            .I(N__47464));
    Span4Mux_v I__11050 (
            .O(N__47542),
            .I(N__47464));
    Span4Mux_h I__11049 (
            .O(N__47533),
            .I(N__47464));
    Span4Mux_v I__11048 (
            .O(N__47520),
            .I(N__47464));
    Span4Mux_h I__11047 (
            .O(N__47509),
            .I(N__47464));
    InMux I__11046 (
            .O(N__47508),
            .I(N__47461));
    Span4Mux_h I__11045 (
            .O(N__47503),
            .I(N__47456));
    Span4Mux_h I__11044 (
            .O(N__47498),
            .I(N__47456));
    LocalMux I__11043 (
            .O(N__47495),
            .I(comm_cmd_2));
    LocalMux I__11042 (
            .O(N__47488),
            .I(comm_cmd_2));
    Odrv12 I__11041 (
            .O(N__47479),
            .I(comm_cmd_2));
    Odrv4 I__11040 (
            .O(N__47464),
            .I(comm_cmd_2));
    LocalMux I__11039 (
            .O(N__47461),
            .I(comm_cmd_2));
    Odrv4 I__11038 (
            .O(N__47456),
            .I(comm_cmd_2));
    InMux I__11037 (
            .O(N__47443),
            .I(N__47440));
    LocalMux I__11036 (
            .O(N__47440),
            .I(N__47437));
    Span4Mux_h I__11035 (
            .O(N__47437),
            .I(N__47434));
    Odrv4 I__11034 (
            .O(N__47434),
            .I(buf_data_iac_7));
    CascadeMux I__11033 (
            .O(N__47431),
            .I(n22_adj_1590_cascade_));
    InMux I__11032 (
            .O(N__47428),
            .I(N__47425));
    LocalMux I__11031 (
            .O(N__47425),
            .I(N__47422));
    Span4Mux_v I__11030 (
            .O(N__47422),
            .I(N__47419));
    Span4Mux_h I__11029 (
            .O(N__47419),
            .I(N__47416));
    Odrv4 I__11028 (
            .O(N__47416),
            .I(n30_adj_1591));
    InMux I__11027 (
            .O(N__47413),
            .I(N__47409));
    InMux I__11026 (
            .O(N__47412),
            .I(N__47406));
    LocalMux I__11025 (
            .O(N__47409),
            .I(N__47403));
    LocalMux I__11024 (
            .O(N__47406),
            .I(N__47399));
    Span4Mux_h I__11023 (
            .O(N__47403),
            .I(N__47396));
    InMux I__11022 (
            .O(N__47402),
            .I(N__47393));
    Span4Mux_h I__11021 (
            .O(N__47399),
            .I(N__47390));
    Span4Mux_h I__11020 (
            .O(N__47396),
            .I(N__47387));
    LocalMux I__11019 (
            .O(N__47393),
            .I(data_cntvec_6));
    Odrv4 I__11018 (
            .O(N__47390),
            .I(data_cntvec_6));
    Odrv4 I__11017 (
            .O(N__47387),
            .I(data_cntvec_6));
    InMux I__11016 (
            .O(N__47380),
            .I(n19301));
    InMux I__11015 (
            .O(N__47377),
            .I(N__47373));
    InMux I__11014 (
            .O(N__47376),
            .I(N__47370));
    LocalMux I__11013 (
            .O(N__47373),
            .I(N__47366));
    LocalMux I__11012 (
            .O(N__47370),
            .I(N__47363));
    InMux I__11011 (
            .O(N__47369),
            .I(N__47360));
    Span4Mux_h I__11010 (
            .O(N__47366),
            .I(N__47357));
    Span4Mux_v I__11009 (
            .O(N__47363),
            .I(N__47354));
    LocalMux I__11008 (
            .O(N__47360),
            .I(data_cntvec_7));
    Odrv4 I__11007 (
            .O(N__47357),
            .I(data_cntvec_7));
    Odrv4 I__11006 (
            .O(N__47354),
            .I(data_cntvec_7));
    InMux I__11005 (
            .O(N__47347),
            .I(n19302));
    InMux I__11004 (
            .O(N__47344),
            .I(N__47340));
    InMux I__11003 (
            .O(N__47343),
            .I(N__47337));
    LocalMux I__11002 (
            .O(N__47340),
            .I(N__47333));
    LocalMux I__11001 (
            .O(N__47337),
            .I(N__47330));
    InMux I__11000 (
            .O(N__47336),
            .I(N__47327));
    Span4Mux_h I__10999 (
            .O(N__47333),
            .I(N__47324));
    Span4Mux_h I__10998 (
            .O(N__47330),
            .I(N__47321));
    LocalMux I__10997 (
            .O(N__47327),
            .I(data_cntvec_8));
    Odrv4 I__10996 (
            .O(N__47324),
            .I(data_cntvec_8));
    Odrv4 I__10995 (
            .O(N__47321),
            .I(data_cntvec_8));
    InMux I__10994 (
            .O(N__47314),
            .I(bfn_18_13_0_));
    InMux I__10993 (
            .O(N__47311),
            .I(N__47308));
    LocalMux I__10992 (
            .O(N__47308),
            .I(N__47304));
    InMux I__10991 (
            .O(N__47307),
            .I(N__47301));
    Span4Mux_v I__10990 (
            .O(N__47304),
            .I(N__47298));
    LocalMux I__10989 (
            .O(N__47301),
            .I(N__47292));
    Span4Mux_h I__10988 (
            .O(N__47298),
            .I(N__47292));
    InMux I__10987 (
            .O(N__47297),
            .I(N__47289));
    Span4Mux_h I__10986 (
            .O(N__47292),
            .I(N__47286));
    LocalMux I__10985 (
            .O(N__47289),
            .I(data_cntvec_9));
    Odrv4 I__10984 (
            .O(N__47286),
            .I(data_cntvec_9));
    InMux I__10983 (
            .O(N__47281),
            .I(n19304));
    CascadeMux I__10982 (
            .O(N__47278),
            .I(N__47275));
    InMux I__10981 (
            .O(N__47275),
            .I(N__47271));
    InMux I__10980 (
            .O(N__47274),
            .I(N__47268));
    LocalMux I__10979 (
            .O(N__47271),
            .I(N__47264));
    LocalMux I__10978 (
            .O(N__47268),
            .I(N__47261));
    InMux I__10977 (
            .O(N__47267),
            .I(N__47258));
    Span4Mux_v I__10976 (
            .O(N__47264),
            .I(N__47255));
    Span12Mux_h I__10975 (
            .O(N__47261),
            .I(N__47252));
    LocalMux I__10974 (
            .O(N__47258),
            .I(data_cntvec_10));
    Odrv4 I__10973 (
            .O(N__47255),
            .I(data_cntvec_10));
    Odrv12 I__10972 (
            .O(N__47252),
            .I(data_cntvec_10));
    InMux I__10971 (
            .O(N__47245),
            .I(n19305));
    InMux I__10970 (
            .O(N__47242),
            .I(N__47237));
    InMux I__10969 (
            .O(N__47241),
            .I(N__47234));
    InMux I__10968 (
            .O(N__47240),
            .I(N__47231));
    LocalMux I__10967 (
            .O(N__47237),
            .I(data_cntvec_11));
    LocalMux I__10966 (
            .O(N__47234),
            .I(data_cntvec_11));
    LocalMux I__10965 (
            .O(N__47231),
            .I(data_cntvec_11));
    InMux I__10964 (
            .O(N__47224),
            .I(n19306));
    InMux I__10963 (
            .O(N__47221),
            .I(N__47218));
    LocalMux I__10962 (
            .O(N__47218),
            .I(N__47214));
    InMux I__10961 (
            .O(N__47217),
            .I(N__47211));
    Span4Mux_v I__10960 (
            .O(N__47214),
            .I(N__47208));
    LocalMux I__10959 (
            .O(N__47211),
            .I(data_cntvec_12));
    Odrv4 I__10958 (
            .O(N__47208),
            .I(data_cntvec_12));
    InMux I__10957 (
            .O(N__47203),
            .I(n19307));
    InMux I__10956 (
            .O(N__47200),
            .I(N__47197));
    LocalMux I__10955 (
            .O(N__47197),
            .I(N__47193));
    InMux I__10954 (
            .O(N__47196),
            .I(N__47190));
    Span4Mux_v I__10953 (
            .O(N__47193),
            .I(N__47187));
    LocalMux I__10952 (
            .O(N__47190),
            .I(data_cntvec_13));
    Odrv4 I__10951 (
            .O(N__47187),
            .I(data_cntvec_13));
    InMux I__10950 (
            .O(N__47182),
            .I(n19308));
    CascadeMux I__10949 (
            .O(N__47179),
            .I(n4_adj_1569_cascade_));
    InMux I__10948 (
            .O(N__47176),
            .I(N__47173));
    LocalMux I__10947 (
            .O(N__47173),
            .I(N__47169));
    InMux I__10946 (
            .O(N__47172),
            .I(N__47166));
    Sp12to4 I__10945 (
            .O(N__47169),
            .I(N__47163));
    LocalMux I__10944 (
            .O(N__47166),
            .I(comm_buf_6_1));
    Odrv12 I__10943 (
            .O(N__47163),
            .I(comm_buf_6_1));
    CascadeMux I__10942 (
            .O(N__47158),
            .I(n20792_cascade_));
    InMux I__10941 (
            .O(N__47155),
            .I(N__47152));
    LocalMux I__10940 (
            .O(N__47152),
            .I(N__47149));
    Span4Mux_v I__10939 (
            .O(N__47149),
            .I(N__47146));
    Span4Mux_h I__10938 (
            .O(N__47146),
            .I(N__47143));
    Odrv4 I__10937 (
            .O(N__47143),
            .I(n21994));
    CEMux I__10936 (
            .O(N__47140),
            .I(N__47137));
    LocalMux I__10935 (
            .O(N__47137),
            .I(N__47132));
    CEMux I__10934 (
            .O(N__47136),
            .I(N__47129));
    CEMux I__10933 (
            .O(N__47135),
            .I(N__47125));
    Span4Mux_v I__10932 (
            .O(N__47132),
            .I(N__47119));
    LocalMux I__10931 (
            .O(N__47129),
            .I(N__47119));
    CEMux I__10930 (
            .O(N__47128),
            .I(N__47116));
    LocalMux I__10929 (
            .O(N__47125),
            .I(N__47113));
    CEMux I__10928 (
            .O(N__47124),
            .I(N__47110));
    Span4Mux_v I__10927 (
            .O(N__47119),
            .I(N__47105));
    LocalMux I__10926 (
            .O(N__47116),
            .I(N__47105));
    Span4Mux_v I__10925 (
            .O(N__47113),
            .I(N__47101));
    LocalMux I__10924 (
            .O(N__47110),
            .I(N__47098));
    Span4Mux_v I__10923 (
            .O(N__47105),
            .I(N__47095));
    CEMux I__10922 (
            .O(N__47104),
            .I(N__47092));
    Span4Mux_h I__10921 (
            .O(N__47101),
            .I(N__47085));
    Span4Mux_v I__10920 (
            .O(N__47098),
            .I(N__47085));
    Span4Mux_h I__10919 (
            .O(N__47095),
            .I(N__47085));
    LocalMux I__10918 (
            .O(N__47092),
            .I(N__47082));
    Sp12to4 I__10917 (
            .O(N__47085),
            .I(N__47078));
    Span4Mux_h I__10916 (
            .O(N__47082),
            .I(N__47075));
    InMux I__10915 (
            .O(N__47081),
            .I(N__47072));
    Odrv12 I__10914 (
            .O(N__47078),
            .I(n12322));
    Odrv4 I__10913 (
            .O(N__47075),
            .I(n12322));
    LocalMux I__10912 (
            .O(N__47072),
            .I(n12322));
    SRMux I__10911 (
            .O(N__47065),
            .I(N__47062));
    LocalMux I__10910 (
            .O(N__47062),
            .I(N__47058));
    SRMux I__10909 (
            .O(N__47061),
            .I(N__47053));
    Span4Mux_v I__10908 (
            .O(N__47058),
            .I(N__47049));
    SRMux I__10907 (
            .O(N__47057),
            .I(N__47045));
    SRMux I__10906 (
            .O(N__47056),
            .I(N__47042));
    LocalMux I__10905 (
            .O(N__47053),
            .I(N__47039));
    SRMux I__10904 (
            .O(N__47052),
            .I(N__47036));
    Span4Mux_h I__10903 (
            .O(N__47049),
            .I(N__47033));
    SRMux I__10902 (
            .O(N__47048),
            .I(N__47030));
    LocalMux I__10901 (
            .O(N__47045),
            .I(N__47027));
    LocalMux I__10900 (
            .O(N__47042),
            .I(N__47024));
    Span4Mux_h I__10899 (
            .O(N__47039),
            .I(N__47019));
    LocalMux I__10898 (
            .O(N__47036),
            .I(N__47019));
    Span4Mux_v I__10897 (
            .O(N__47033),
            .I(N__47014));
    LocalMux I__10896 (
            .O(N__47030),
            .I(N__47014));
    Span4Mux_v I__10895 (
            .O(N__47027),
            .I(N__47011));
    Span4Mux_h I__10894 (
            .O(N__47024),
            .I(N__47006));
    Span4Mux_h I__10893 (
            .O(N__47019),
            .I(N__47006));
    Span4Mux_h I__10892 (
            .O(N__47014),
            .I(N__47003));
    Odrv4 I__10891 (
            .O(N__47011),
            .I(n14784));
    Odrv4 I__10890 (
            .O(N__47006),
            .I(n14784));
    Odrv4 I__10889 (
            .O(N__47003),
            .I(n14784));
    InMux I__10888 (
            .O(N__46996),
            .I(N__46993));
    LocalMux I__10887 (
            .O(N__46993),
            .I(N__46990));
    Odrv4 I__10886 (
            .O(N__46990),
            .I(n21069));
    CascadeMux I__10885 (
            .O(N__46987),
            .I(N__46983));
    InMux I__10884 (
            .O(N__46986),
            .I(N__46980));
    InMux I__10883 (
            .O(N__46983),
            .I(N__46977));
    LocalMux I__10882 (
            .O(N__46980),
            .I(N__46972));
    LocalMux I__10881 (
            .O(N__46977),
            .I(N__46969));
    InMux I__10880 (
            .O(N__46976),
            .I(N__46963));
    InMux I__10879 (
            .O(N__46975),
            .I(N__46963));
    Span4Mux_v I__10878 (
            .O(N__46972),
            .I(N__46960));
    Span4Mux_h I__10877 (
            .O(N__46969),
            .I(N__46957));
    InMux I__10876 (
            .O(N__46968),
            .I(N__46953));
    LocalMux I__10875 (
            .O(N__46963),
            .I(N__46946));
    Span4Mux_h I__10874 (
            .O(N__46960),
            .I(N__46946));
    Span4Mux_h I__10873 (
            .O(N__46957),
            .I(N__46946));
    InMux I__10872 (
            .O(N__46956),
            .I(N__46943));
    LocalMux I__10871 (
            .O(N__46953),
            .I(iac_raw_buf_N_728));
    Odrv4 I__10870 (
            .O(N__46946),
            .I(iac_raw_buf_N_728));
    LocalMux I__10869 (
            .O(N__46943),
            .I(iac_raw_buf_N_728));
    InMux I__10868 (
            .O(N__46936),
            .I(N__46932));
    InMux I__10867 (
            .O(N__46935),
            .I(N__46929));
    LocalMux I__10866 (
            .O(N__46932),
            .I(N__46923));
    LocalMux I__10865 (
            .O(N__46929),
            .I(N__46923));
    InMux I__10864 (
            .O(N__46928),
            .I(N__46920));
    Span4Mux_h I__10863 (
            .O(N__46923),
            .I(N__46917));
    LocalMux I__10862 (
            .O(N__46920),
            .I(data_cntvec_0));
    Odrv4 I__10861 (
            .O(N__46917),
            .I(data_cntvec_0));
    InMux I__10860 (
            .O(N__46912),
            .I(N__46909));
    LocalMux I__10859 (
            .O(N__46909),
            .I(N__46904));
    InMux I__10858 (
            .O(N__46908),
            .I(N__46901));
    InMux I__10857 (
            .O(N__46907),
            .I(N__46898));
    Span4Mux_h I__10856 (
            .O(N__46904),
            .I(N__46895));
    LocalMux I__10855 (
            .O(N__46901),
            .I(N__46892));
    LocalMux I__10854 (
            .O(N__46898),
            .I(data_cntvec_1));
    Odrv4 I__10853 (
            .O(N__46895),
            .I(data_cntvec_1));
    Odrv12 I__10852 (
            .O(N__46892),
            .I(data_cntvec_1));
    InMux I__10851 (
            .O(N__46885),
            .I(n19296));
    InMux I__10850 (
            .O(N__46882),
            .I(N__46878));
    InMux I__10849 (
            .O(N__46881),
            .I(N__46875));
    LocalMux I__10848 (
            .O(N__46878),
            .I(N__46872));
    LocalMux I__10847 (
            .O(N__46875),
            .I(N__46866));
    Span4Mux_h I__10846 (
            .O(N__46872),
            .I(N__46866));
    InMux I__10845 (
            .O(N__46871),
            .I(N__46863));
    Span4Mux_h I__10844 (
            .O(N__46866),
            .I(N__46860));
    LocalMux I__10843 (
            .O(N__46863),
            .I(data_cntvec_2));
    Odrv4 I__10842 (
            .O(N__46860),
            .I(data_cntvec_2));
    InMux I__10841 (
            .O(N__46855),
            .I(n19297));
    InMux I__10840 (
            .O(N__46852),
            .I(N__46848));
    InMux I__10839 (
            .O(N__46851),
            .I(N__46845));
    LocalMux I__10838 (
            .O(N__46848),
            .I(N__46842));
    LocalMux I__10837 (
            .O(N__46845),
            .I(N__46839));
    Span4Mux_v I__10836 (
            .O(N__46842),
            .I(N__46835));
    Span4Mux_h I__10835 (
            .O(N__46839),
            .I(N__46832));
    InMux I__10834 (
            .O(N__46838),
            .I(N__46829));
    Span4Mux_h I__10833 (
            .O(N__46835),
            .I(N__46826));
    Span4Mux_h I__10832 (
            .O(N__46832),
            .I(N__46823));
    LocalMux I__10831 (
            .O(N__46829),
            .I(data_cntvec_3));
    Odrv4 I__10830 (
            .O(N__46826),
            .I(data_cntvec_3));
    Odrv4 I__10829 (
            .O(N__46823),
            .I(data_cntvec_3));
    InMux I__10828 (
            .O(N__46816),
            .I(n19298));
    InMux I__10827 (
            .O(N__46813),
            .I(N__46809));
    InMux I__10826 (
            .O(N__46812),
            .I(N__46806));
    LocalMux I__10825 (
            .O(N__46809),
            .I(N__46803));
    LocalMux I__10824 (
            .O(N__46806),
            .I(N__46797));
    Span4Mux_h I__10823 (
            .O(N__46803),
            .I(N__46797));
    InMux I__10822 (
            .O(N__46802),
            .I(N__46794));
    Span4Mux_h I__10821 (
            .O(N__46797),
            .I(N__46791));
    LocalMux I__10820 (
            .O(N__46794),
            .I(data_cntvec_4));
    Odrv4 I__10819 (
            .O(N__46791),
            .I(data_cntvec_4));
    InMux I__10818 (
            .O(N__46786),
            .I(n19299));
    InMux I__10817 (
            .O(N__46783),
            .I(N__46779));
    InMux I__10816 (
            .O(N__46782),
            .I(N__46776));
    LocalMux I__10815 (
            .O(N__46779),
            .I(N__46773));
    LocalMux I__10814 (
            .O(N__46776),
            .I(N__46767));
    Span4Mux_h I__10813 (
            .O(N__46773),
            .I(N__46767));
    InMux I__10812 (
            .O(N__46772),
            .I(N__46764));
    Span4Mux_h I__10811 (
            .O(N__46767),
            .I(N__46761));
    LocalMux I__10810 (
            .O(N__46764),
            .I(data_cntvec_5));
    Odrv4 I__10809 (
            .O(N__46761),
            .I(data_cntvec_5));
    InMux I__10808 (
            .O(N__46756),
            .I(n19300));
    InMux I__10807 (
            .O(N__46753),
            .I(N__46750));
    LocalMux I__10806 (
            .O(N__46750),
            .I(N__46747));
    Span4Mux_h I__10805 (
            .O(N__46747),
            .I(N__46744));
    Odrv4 I__10804 (
            .O(N__46744),
            .I(n4_adj_1566));
    CascadeMux I__10803 (
            .O(N__46741),
            .I(n22063_cascade_));
    InMux I__10802 (
            .O(N__46738),
            .I(N__46735));
    LocalMux I__10801 (
            .O(N__46735),
            .I(N__46731));
    InMux I__10800 (
            .O(N__46734),
            .I(N__46728));
    Span4Mux_h I__10799 (
            .O(N__46731),
            .I(N__46725));
    LocalMux I__10798 (
            .O(N__46728),
            .I(N__46720));
    Span4Mux_h I__10797 (
            .O(N__46725),
            .I(N__46720));
    Odrv4 I__10796 (
            .O(N__46720),
            .I(comm_buf_6_4));
    CascadeMux I__10795 (
            .O(N__46717),
            .I(N__46714));
    InMux I__10794 (
            .O(N__46714),
            .I(N__46711));
    LocalMux I__10793 (
            .O(N__46711),
            .I(n21081));
    CascadeMux I__10792 (
            .O(N__46708),
            .I(N__46704));
    InMux I__10791 (
            .O(N__46707),
            .I(N__46701));
    InMux I__10790 (
            .O(N__46704),
            .I(N__46697));
    LocalMux I__10789 (
            .O(N__46701),
            .I(N__46694));
    InMux I__10788 (
            .O(N__46700),
            .I(N__46691));
    LocalMux I__10787 (
            .O(N__46697),
            .I(N__46688));
    Span4Mux_v I__10786 (
            .O(N__46694),
            .I(N__46683));
    LocalMux I__10785 (
            .O(N__46691),
            .I(N__46683));
    Span4Mux_v I__10784 (
            .O(N__46688),
            .I(N__46680));
    Sp12to4 I__10783 (
            .O(N__46683),
            .I(N__46677));
    Span4Mux_h I__10782 (
            .O(N__46680),
            .I(N__46674));
    Span12Mux_h I__10781 (
            .O(N__46677),
            .I(N__46671));
    Odrv4 I__10780 (
            .O(N__46674),
            .I(comm_buf_0_4));
    Odrv12 I__10779 (
            .O(N__46671),
            .I(comm_buf_0_4));
    InMux I__10778 (
            .O(N__46666),
            .I(N__46661));
    CascadeMux I__10777 (
            .O(N__46665),
            .I(N__46658));
    InMux I__10776 (
            .O(N__46664),
            .I(N__46655));
    LocalMux I__10775 (
            .O(N__46661),
            .I(N__46651));
    InMux I__10774 (
            .O(N__46658),
            .I(N__46648));
    LocalMux I__10773 (
            .O(N__46655),
            .I(N__46643));
    InMux I__10772 (
            .O(N__46654),
            .I(N__46640));
    Span4Mux_v I__10771 (
            .O(N__46651),
            .I(N__46637));
    LocalMux I__10770 (
            .O(N__46648),
            .I(N__46634));
    InMux I__10769 (
            .O(N__46647),
            .I(N__46631));
    InMux I__10768 (
            .O(N__46646),
            .I(N__46628));
    Span4Mux_v I__10767 (
            .O(N__46643),
            .I(N__46625));
    LocalMux I__10766 (
            .O(N__46640),
            .I(N__46622));
    Span4Mux_h I__10765 (
            .O(N__46637),
            .I(N__46619));
    Span4Mux_h I__10764 (
            .O(N__46634),
            .I(N__46614));
    LocalMux I__10763 (
            .O(N__46631),
            .I(N__46614));
    LocalMux I__10762 (
            .O(N__46628),
            .I(N__46611));
    Span4Mux_h I__10761 (
            .O(N__46625),
            .I(N__46606));
    Span4Mux_h I__10760 (
            .O(N__46622),
            .I(N__46606));
    Odrv4 I__10759 (
            .O(N__46619),
            .I(comm_buf_1_4));
    Odrv4 I__10758 (
            .O(N__46614),
            .I(comm_buf_1_4));
    Odrv12 I__10757 (
            .O(N__46611),
            .I(comm_buf_1_4));
    Odrv4 I__10756 (
            .O(N__46606),
            .I(comm_buf_1_4));
    InMux I__10755 (
            .O(N__46597),
            .I(N__46594));
    LocalMux I__10754 (
            .O(N__46594),
            .I(n1_adj_1564));
    CascadeMux I__10753 (
            .O(N__46591),
            .I(n18824_cascade_));
    InMux I__10752 (
            .O(N__46588),
            .I(N__46585));
    LocalMux I__10751 (
            .O(N__46585),
            .I(N__46582));
    Span4Mux_v I__10750 (
            .O(N__46582),
            .I(N__46578));
    InMux I__10749 (
            .O(N__46581),
            .I(N__46575));
    Span4Mux_h I__10748 (
            .O(N__46578),
            .I(N__46570));
    LocalMux I__10747 (
            .O(N__46575),
            .I(N__46570));
    Odrv4 I__10746 (
            .O(N__46570),
            .I(n20507));
    CascadeMux I__10745 (
            .O(N__46567),
            .I(N__46564));
    InMux I__10744 (
            .O(N__46564),
            .I(N__46561));
    LocalMux I__10743 (
            .O(N__46561),
            .I(N__46558));
    Span4Mux_h I__10742 (
            .O(N__46558),
            .I(N__46555));
    Odrv4 I__10741 (
            .O(N__46555),
            .I(comm_buf_2_4));
    InMux I__10740 (
            .O(N__46552),
            .I(N__46549));
    LocalMux I__10739 (
            .O(N__46549),
            .I(N__46546));
    Span4Mux_v I__10738 (
            .O(N__46546),
            .I(N__46543));
    Span4Mux_h I__10737 (
            .O(N__46543),
            .I(N__46540));
    Odrv4 I__10736 (
            .O(N__46540),
            .I(comm_buf_3_4));
    InMux I__10735 (
            .O(N__46537),
            .I(N__46534));
    LocalMux I__10734 (
            .O(N__46534),
            .I(n2_adj_1565));
    InMux I__10733 (
            .O(N__46531),
            .I(N__46528));
    LocalMux I__10732 (
            .O(N__46528),
            .I(N__46525));
    Odrv12 I__10731 (
            .O(N__46525),
            .I(comm_buf_5_1));
    InMux I__10730 (
            .O(N__46522),
            .I(N__46519));
    LocalMux I__10729 (
            .O(N__46519),
            .I(N__46516));
    Span4Mux_h I__10728 (
            .O(N__46516),
            .I(N__46513));
    Odrv4 I__10727 (
            .O(N__46513),
            .I(comm_buf_4_1));
    CascadeMux I__10726 (
            .O(N__46510),
            .I(n4_adj_1483_cascade_));
    InMux I__10725 (
            .O(N__46507),
            .I(N__46504));
    LocalMux I__10724 (
            .O(N__46504),
            .I(N__46501));
    Span4Mux_h I__10723 (
            .O(N__46501),
            .I(N__46497));
    InMux I__10722 (
            .O(N__46500),
            .I(N__46494));
    Span4Mux_h I__10721 (
            .O(N__46497),
            .I(N__46491));
    LocalMux I__10720 (
            .O(N__46494),
            .I(N__46488));
    Odrv4 I__10719 (
            .O(N__46491),
            .I(n12205));
    Odrv4 I__10718 (
            .O(N__46488),
            .I(n12205));
    InMux I__10717 (
            .O(N__46483),
            .I(N__46480));
    LocalMux I__10716 (
            .O(N__46480),
            .I(N__46477));
    Span12Mux_v I__10715 (
            .O(N__46477),
            .I(N__46474));
    Odrv12 I__10714 (
            .O(N__46474),
            .I(n4));
    CascadeMux I__10713 (
            .O(N__46471),
            .I(n20510_cascade_));
    InMux I__10712 (
            .O(N__46468),
            .I(N__46462));
    InMux I__10711 (
            .O(N__46467),
            .I(N__46462));
    LocalMux I__10710 (
            .O(N__46462),
            .I(N__46459));
    Span4Mux_v I__10709 (
            .O(N__46459),
            .I(N__46456));
    Odrv4 I__10708 (
            .O(N__46456),
            .I(n3));
    CEMux I__10707 (
            .O(N__46453),
            .I(N__46450));
    LocalMux I__10706 (
            .O(N__46450),
            .I(N__46447));
    Span4Mux_h I__10705 (
            .O(N__46447),
            .I(N__46444));
    Span4Mux_h I__10704 (
            .O(N__46444),
            .I(N__46441));
    Odrv4 I__10703 (
            .O(N__46441),
            .I(n20534));
    InMux I__10702 (
            .O(N__46438),
            .I(N__46435));
    LocalMux I__10701 (
            .O(N__46435),
            .I(n11810));
    CascadeMux I__10700 (
            .O(N__46432),
            .I(n11810_cascade_));
    InMux I__10699 (
            .O(N__46429),
            .I(N__46426));
    LocalMux I__10698 (
            .O(N__46426),
            .I(N__46423));
    Span4Mux_v I__10697 (
            .O(N__46423),
            .I(N__46419));
    InMux I__10696 (
            .O(N__46422),
            .I(N__46416));
    Span4Mux_h I__10695 (
            .O(N__46419),
            .I(N__46413));
    LocalMux I__10694 (
            .O(N__46416),
            .I(n20650));
    Odrv4 I__10693 (
            .O(N__46413),
            .I(n20650));
    CascadeMux I__10692 (
            .O(N__46408),
            .I(n20672_cascade_));
    InMux I__10691 (
            .O(N__46405),
            .I(N__46402));
    LocalMux I__10690 (
            .O(N__46402),
            .I(n20510));
    InMux I__10689 (
            .O(N__46399),
            .I(N__46395));
    InMux I__10688 (
            .O(N__46398),
            .I(N__46392));
    LocalMux I__10687 (
            .O(N__46395),
            .I(n20585));
    LocalMux I__10686 (
            .O(N__46392),
            .I(n20585));
    InMux I__10685 (
            .O(N__46387),
            .I(N__46384));
    LocalMux I__10684 (
            .O(N__46384),
            .I(n11824));
    InMux I__10683 (
            .O(N__46381),
            .I(N__46378));
    LocalMux I__10682 (
            .O(N__46378),
            .I(N__46367));
    InMux I__10681 (
            .O(N__46377),
            .I(N__46364));
    InMux I__10680 (
            .O(N__46376),
            .I(N__46349));
    InMux I__10679 (
            .O(N__46375),
            .I(N__46349));
    InMux I__10678 (
            .O(N__46374),
            .I(N__46349));
    InMux I__10677 (
            .O(N__46373),
            .I(N__46349));
    InMux I__10676 (
            .O(N__46372),
            .I(N__46349));
    InMux I__10675 (
            .O(N__46371),
            .I(N__46349));
    InMux I__10674 (
            .O(N__46370),
            .I(N__46349));
    Odrv12 I__10673 (
            .O(N__46367),
            .I(\comm_spi.bit_cnt_3 ));
    LocalMux I__10672 (
            .O(N__46364),
            .I(\comm_spi.bit_cnt_3 ));
    LocalMux I__10671 (
            .O(N__46349),
            .I(\comm_spi.bit_cnt_3 ));
    InMux I__10670 (
            .O(N__46342),
            .I(N__46339));
    LocalMux I__10669 (
            .O(N__46339),
            .I(N__46336));
    Span4Mux_h I__10668 (
            .O(N__46336),
            .I(N__46333));
    Span4Mux_h I__10667 (
            .O(N__46333),
            .I(N__46323));
    InMux I__10666 (
            .O(N__46332),
            .I(N__46308));
    InMux I__10665 (
            .O(N__46331),
            .I(N__46308));
    InMux I__10664 (
            .O(N__46330),
            .I(N__46308));
    InMux I__10663 (
            .O(N__46329),
            .I(N__46308));
    InMux I__10662 (
            .O(N__46328),
            .I(N__46308));
    InMux I__10661 (
            .O(N__46327),
            .I(N__46308));
    InMux I__10660 (
            .O(N__46326),
            .I(N__46308));
    Odrv4 I__10659 (
            .O(N__46323),
            .I(\comm_spi.n16858 ));
    LocalMux I__10658 (
            .O(N__46308),
            .I(\comm_spi.n16858 ));
    InMux I__10657 (
            .O(N__46303),
            .I(N__46300));
    LocalMux I__10656 (
            .O(N__46300),
            .I(N__46297));
    Odrv4 I__10655 (
            .O(N__46297),
            .I(n21087));
    InMux I__10654 (
            .O(N__46294),
            .I(N__46290));
    InMux I__10653 (
            .O(N__46293),
            .I(N__46287));
    LocalMux I__10652 (
            .O(N__46290),
            .I(\comm_spi.n14620 ));
    LocalMux I__10651 (
            .O(N__46287),
            .I(\comm_spi.n14620 ));
    SRMux I__10650 (
            .O(N__46282),
            .I(N__46279));
    LocalMux I__10649 (
            .O(N__46279),
            .I(N__46276));
    Odrv12 I__10648 (
            .O(N__46276),
            .I(\comm_spi.data_tx_7__N_772 ));
    InMux I__10647 (
            .O(N__46273),
            .I(N__46270));
    LocalMux I__10646 (
            .O(N__46270),
            .I(N__46266));
    InMux I__10645 (
            .O(N__46269),
            .I(N__46263));
    Span4Mux_v I__10644 (
            .O(N__46266),
            .I(N__46258));
    LocalMux I__10643 (
            .O(N__46263),
            .I(N__46258));
    Span4Mux_h I__10642 (
            .O(N__46258),
            .I(N__46254));
    InMux I__10641 (
            .O(N__46257),
            .I(N__46251));
    Odrv4 I__10640 (
            .O(N__46254),
            .I(\comm_spi.n22638 ));
    LocalMux I__10639 (
            .O(N__46251),
            .I(\comm_spi.n22638 ));
    InMux I__10638 (
            .O(N__46246),
            .I(N__46243));
    LocalMux I__10637 (
            .O(N__46243),
            .I(N__46239));
    InMux I__10636 (
            .O(N__46242),
            .I(N__46236));
    Odrv4 I__10635 (
            .O(N__46239),
            .I(\comm_spi.n14619 ));
    LocalMux I__10634 (
            .O(N__46236),
            .I(\comm_spi.n14619 ));
    InMux I__10633 (
            .O(N__46231),
            .I(N__46228));
    LocalMux I__10632 (
            .O(N__46228),
            .I(N__46224));
    InMux I__10631 (
            .O(N__46227),
            .I(N__46221));
    Odrv4 I__10630 (
            .O(N__46224),
            .I(\comm_spi.n14615 ));
    LocalMux I__10629 (
            .O(N__46221),
            .I(\comm_spi.n14615 ));
    SRMux I__10628 (
            .O(N__46216),
            .I(N__46213));
    LocalMux I__10627 (
            .O(N__46213),
            .I(N__46210));
    Odrv12 I__10626 (
            .O(N__46210),
            .I(\comm_spi.data_tx_7__N_761 ));
    InMux I__10625 (
            .O(N__46207),
            .I(N__46203));
    InMux I__10624 (
            .O(N__46206),
            .I(N__46200));
    LocalMux I__10623 (
            .O(N__46203),
            .I(N__46195));
    LocalMux I__10622 (
            .O(N__46200),
            .I(N__46195));
    Span4Mux_v I__10621 (
            .O(N__46195),
            .I(N__46192));
    Sp12to4 I__10620 (
            .O(N__46192),
            .I(N__46188));
    InMux I__10619 (
            .O(N__46191),
            .I(N__46185));
    Odrv12 I__10618 (
            .O(N__46188),
            .I(\comm_spi.n22641 ));
    LocalMux I__10617 (
            .O(N__46185),
            .I(\comm_spi.n22641 ));
    InMux I__10616 (
            .O(N__46180),
            .I(N__46176));
    InMux I__10615 (
            .O(N__46179),
            .I(N__46173));
    LocalMux I__10614 (
            .O(N__46176),
            .I(N__46168));
    LocalMux I__10613 (
            .O(N__46173),
            .I(N__46168));
    Span4Mux_v I__10612 (
            .O(N__46168),
            .I(N__46165));
    Sp12to4 I__10611 (
            .O(N__46165),
            .I(N__46162));
    Odrv12 I__10610 (
            .O(N__46162),
            .I(\comm_spi.n14611 ));
    InMux I__10609 (
            .O(N__46159),
            .I(N__46156));
    LocalMux I__10608 (
            .O(N__46156),
            .I(N__46152));
    InMux I__10607 (
            .O(N__46155),
            .I(N__46149));
    Span4Mux_v I__10606 (
            .O(N__46152),
            .I(N__46146));
    LocalMux I__10605 (
            .O(N__46149),
            .I(N__46143));
    Odrv4 I__10604 (
            .O(N__46146),
            .I(\comm_spi.n14612 ));
    Odrv12 I__10603 (
            .O(N__46143),
            .I(\comm_spi.n14612 ));
    InMux I__10602 (
            .O(N__46138),
            .I(N__46134));
    InMux I__10601 (
            .O(N__46137),
            .I(N__46131));
    LocalMux I__10600 (
            .O(N__46134),
            .I(N__46128));
    LocalMux I__10599 (
            .O(N__46131),
            .I(N__46125));
    Odrv4 I__10598 (
            .O(N__46128),
            .I(\comm_spi.n14616 ));
    Odrv4 I__10597 (
            .O(N__46125),
            .I(\comm_spi.n14616 ));
    InMux I__10596 (
            .O(N__46120),
            .I(N__46117));
    LocalMux I__10595 (
            .O(N__46117),
            .I(N__46114));
    Odrv4 I__10594 (
            .O(N__46114),
            .I(n20641));
    CascadeMux I__10593 (
            .O(N__46111),
            .I(N__46108));
    InMux I__10592 (
            .O(N__46108),
            .I(N__46105));
    LocalMux I__10591 (
            .O(N__46105),
            .I(N__46102));
    Span4Mux_h I__10590 (
            .O(N__46102),
            .I(N__46099));
    Odrv4 I__10589 (
            .O(N__46099),
            .I(n17656));
    InMux I__10588 (
            .O(N__46096),
            .I(N__46093));
    LocalMux I__10587 (
            .O(N__46093),
            .I(N__46090));
    Odrv4 I__10586 (
            .O(N__46090),
            .I(n21162));
    CascadeMux I__10585 (
            .O(N__46087),
            .I(n17658_cascade_));
    InMux I__10584 (
            .O(N__46084),
            .I(N__46081));
    LocalMux I__10583 (
            .O(N__46081),
            .I(N__46078));
    Span4Mux_v I__10582 (
            .O(N__46078),
            .I(N__46074));
    InMux I__10581 (
            .O(N__46077),
            .I(N__46071));
    Sp12to4 I__10580 (
            .O(N__46074),
            .I(N__46066));
    LocalMux I__10579 (
            .O(N__46071),
            .I(N__46066));
    Odrv12 I__10578 (
            .O(N__46066),
            .I(n20653));
    CascadeMux I__10577 (
            .O(N__46063),
            .I(n12220_cascade_));
    InMux I__10576 (
            .O(N__46060),
            .I(N__46057));
    LocalMux I__10575 (
            .O(N__46057),
            .I(n17338));
    InMux I__10574 (
            .O(N__46054),
            .I(N__46050));
    InMux I__10573 (
            .O(N__46053),
            .I(N__46047));
    LocalMux I__10572 (
            .O(N__46050),
            .I(n17336));
    LocalMux I__10571 (
            .O(N__46047),
            .I(n17336));
    InMux I__10570 (
            .O(N__46042),
            .I(N__46039));
    LocalMux I__10569 (
            .O(N__46039),
            .I(N__46034));
    InMux I__10568 (
            .O(N__46038),
            .I(N__46031));
    InMux I__10567 (
            .O(N__46037),
            .I(N__46028));
    Odrv4 I__10566 (
            .O(N__46034),
            .I(data_index_5));
    LocalMux I__10565 (
            .O(N__46031),
            .I(data_index_5));
    LocalMux I__10564 (
            .O(N__46028),
            .I(data_index_5));
    InMux I__10563 (
            .O(N__46021),
            .I(N__46010));
    InMux I__10562 (
            .O(N__46020),
            .I(N__46007));
    InMux I__10561 (
            .O(N__46019),
            .I(N__45994));
    InMux I__10560 (
            .O(N__46018),
            .I(N__45994));
    InMux I__10559 (
            .O(N__46017),
            .I(N__45994));
    InMux I__10558 (
            .O(N__46016),
            .I(N__45994));
    InMux I__10557 (
            .O(N__46015),
            .I(N__45994));
    InMux I__10556 (
            .O(N__46014),
            .I(N__45991));
    InMux I__10555 (
            .O(N__46013),
            .I(N__45988));
    LocalMux I__10554 (
            .O(N__46010),
            .I(N__45982));
    LocalMux I__10553 (
            .O(N__46007),
            .I(N__45982));
    InMux I__10552 (
            .O(N__46006),
            .I(N__45977));
    InMux I__10551 (
            .O(N__46005),
            .I(N__45977));
    LocalMux I__10550 (
            .O(N__45994),
            .I(N__45974));
    LocalMux I__10549 (
            .O(N__45991),
            .I(N__45969));
    LocalMux I__10548 (
            .O(N__45988),
            .I(N__45969));
    InMux I__10547 (
            .O(N__45987),
            .I(N__45966));
    Span4Mux_v I__10546 (
            .O(N__45982),
            .I(N__45960));
    LocalMux I__10545 (
            .O(N__45977),
            .I(N__45960));
    Span4Mux_h I__10544 (
            .O(N__45974),
            .I(N__45953));
    Span4Mux_v I__10543 (
            .O(N__45969),
            .I(N__45953));
    LocalMux I__10542 (
            .O(N__45966),
            .I(N__45953));
    InMux I__10541 (
            .O(N__45965),
            .I(N__45950));
    Sp12to4 I__10540 (
            .O(N__45960),
            .I(N__45947));
    Span4Mux_h I__10539 (
            .O(N__45953),
            .I(N__45942));
    LocalMux I__10538 (
            .O(N__45950),
            .I(N__45942));
    Odrv12 I__10537 (
            .O(N__45947),
            .I(n16708));
    Odrv4 I__10536 (
            .O(N__45942),
            .I(n16708));
    InMux I__10535 (
            .O(N__45937),
            .I(N__45934));
    LocalMux I__10534 (
            .O(N__45934),
            .I(N__45930));
    InMux I__10533 (
            .O(N__45933),
            .I(N__45927));
    Span4Mux_h I__10532 (
            .O(N__45930),
            .I(N__45924));
    LocalMux I__10531 (
            .O(N__45927),
            .I(N__45921));
    Odrv4 I__10530 (
            .O(N__45924),
            .I(n20626));
    Odrv12 I__10529 (
            .O(N__45921),
            .I(n20626));
    CascadeMux I__10528 (
            .O(N__45916),
            .I(N__45908));
    CascadeMux I__10527 (
            .O(N__45915),
            .I(N__45905));
    CascadeMux I__10526 (
            .O(N__45914),
            .I(N__45902));
    CascadeMux I__10525 (
            .O(N__45913),
            .I(N__45897));
    InMux I__10524 (
            .O(N__45912),
            .I(N__45892));
    InMux I__10523 (
            .O(N__45911),
            .I(N__45888));
    InMux I__10522 (
            .O(N__45908),
            .I(N__45877));
    InMux I__10521 (
            .O(N__45905),
            .I(N__45877));
    InMux I__10520 (
            .O(N__45902),
            .I(N__45877));
    InMux I__10519 (
            .O(N__45901),
            .I(N__45877));
    InMux I__10518 (
            .O(N__45900),
            .I(N__45877));
    InMux I__10517 (
            .O(N__45897),
            .I(N__45871));
    InMux I__10516 (
            .O(N__45896),
            .I(N__45871));
    InMux I__10515 (
            .O(N__45895),
            .I(N__45868));
    LocalMux I__10514 (
            .O(N__45892),
            .I(N__45865));
    InMux I__10513 (
            .O(N__45891),
            .I(N__45862));
    LocalMux I__10512 (
            .O(N__45888),
            .I(N__45859));
    LocalMux I__10511 (
            .O(N__45877),
            .I(N__45856));
    InMux I__10510 (
            .O(N__45876),
            .I(N__45853));
    LocalMux I__10509 (
            .O(N__45871),
            .I(N__45850));
    LocalMux I__10508 (
            .O(N__45868),
            .I(N__45847));
    Span4Mux_h I__10507 (
            .O(N__45865),
            .I(N__45844));
    LocalMux I__10506 (
            .O(N__45862),
            .I(N__45841));
    Span4Mux_v I__10505 (
            .O(N__45859),
            .I(N__45835));
    Span4Mux_h I__10504 (
            .O(N__45856),
            .I(N__45830));
    LocalMux I__10503 (
            .O(N__45853),
            .I(N__45830));
    Span4Mux_h I__10502 (
            .O(N__45850),
            .I(N__45822));
    Span4Mux_v I__10501 (
            .O(N__45847),
            .I(N__45822));
    Span4Mux_v I__10500 (
            .O(N__45844),
            .I(N__45822));
    Span4Mux_h I__10499 (
            .O(N__45841),
            .I(N__45819));
    InMux I__10498 (
            .O(N__45840),
            .I(N__45816));
    InMux I__10497 (
            .O(N__45839),
            .I(N__45811));
    InMux I__10496 (
            .O(N__45838),
            .I(N__45811));
    Span4Mux_h I__10495 (
            .O(N__45835),
            .I(N__45807));
    Span4Mux_h I__10494 (
            .O(N__45830),
            .I(N__45804));
    InMux I__10493 (
            .O(N__45829),
            .I(N__45801));
    Span4Mux_h I__10492 (
            .O(N__45822),
            .I(N__45798));
    Span4Mux_h I__10491 (
            .O(N__45819),
            .I(N__45795));
    LocalMux I__10490 (
            .O(N__45816),
            .I(N__45790));
    LocalMux I__10489 (
            .O(N__45811),
            .I(N__45790));
    InMux I__10488 (
            .O(N__45810),
            .I(N__45787));
    Odrv4 I__10487 (
            .O(N__45807),
            .I(n11805));
    Odrv4 I__10486 (
            .O(N__45804),
            .I(n11805));
    LocalMux I__10485 (
            .O(N__45801),
            .I(n11805));
    Odrv4 I__10484 (
            .O(N__45798),
            .I(n11805));
    Odrv4 I__10483 (
            .O(N__45795),
            .I(n11805));
    Odrv12 I__10482 (
            .O(N__45790),
            .I(n11805));
    LocalMux I__10481 (
            .O(N__45787),
            .I(n11805));
    CascadeMux I__10480 (
            .O(N__45772),
            .I(N__45769));
    InMux I__10479 (
            .O(N__45769),
            .I(N__45762));
    CascadeMux I__10478 (
            .O(N__45768),
            .I(N__45759));
    InMux I__10477 (
            .O(N__45767),
            .I(N__45756));
    InMux I__10476 (
            .O(N__45766),
            .I(N__45753));
    InMux I__10475 (
            .O(N__45765),
            .I(N__45750));
    LocalMux I__10474 (
            .O(N__45762),
            .I(N__45747));
    InMux I__10473 (
            .O(N__45759),
            .I(N__45744));
    LocalMux I__10472 (
            .O(N__45756),
            .I(N__45741));
    LocalMux I__10471 (
            .O(N__45753),
            .I(N__45738));
    LocalMux I__10470 (
            .O(N__45750),
            .I(N__45735));
    Span4Mux_h I__10469 (
            .O(N__45747),
            .I(N__45728));
    LocalMux I__10468 (
            .O(N__45744),
            .I(N__45728));
    Span4Mux_v I__10467 (
            .O(N__45741),
            .I(N__45728));
    Span4Mux_h I__10466 (
            .O(N__45738),
            .I(N__45724));
    Span4Mux_v I__10465 (
            .O(N__45735),
            .I(N__45721));
    Span4Mux_h I__10464 (
            .O(N__45728),
            .I(N__45718));
    InMux I__10463 (
            .O(N__45727),
            .I(N__45715));
    Span4Mux_v I__10462 (
            .O(N__45724),
            .I(N__45712));
    Span4Mux_v I__10461 (
            .O(N__45721),
            .I(N__45709));
    Span4Mux_h I__10460 (
            .O(N__45718),
            .I(N__45706));
    LocalMux I__10459 (
            .O(N__45715),
            .I(n14_adj_1523));
    Odrv4 I__10458 (
            .O(N__45712),
            .I(n14_adj_1523));
    Odrv4 I__10457 (
            .O(N__45709),
            .I(n14_adj_1523));
    Odrv4 I__10456 (
            .O(N__45706),
            .I(n14_adj_1523));
    InMux I__10455 (
            .O(N__45697),
            .I(N__45688));
    InMux I__10454 (
            .O(N__45696),
            .I(N__45681));
    InMux I__10453 (
            .O(N__45695),
            .I(N__45681));
    InMux I__10452 (
            .O(N__45694),
            .I(N__45681));
    InMux I__10451 (
            .O(N__45693),
            .I(N__45678));
    InMux I__10450 (
            .O(N__45692),
            .I(N__45668));
    InMux I__10449 (
            .O(N__45691),
            .I(N__45668));
    LocalMux I__10448 (
            .O(N__45688),
            .I(N__45661));
    LocalMux I__10447 (
            .O(N__45681),
            .I(N__45661));
    LocalMux I__10446 (
            .O(N__45678),
            .I(N__45661));
    InMux I__10445 (
            .O(N__45677),
            .I(N__45658));
    InMux I__10444 (
            .O(N__45676),
            .I(N__45650));
    InMux I__10443 (
            .O(N__45675),
            .I(N__45650));
    InMux I__10442 (
            .O(N__45674),
            .I(N__45647));
    InMux I__10441 (
            .O(N__45673),
            .I(N__45644));
    LocalMux I__10440 (
            .O(N__45668),
            .I(N__45641));
    Span4Mux_v I__10439 (
            .O(N__45661),
            .I(N__45638));
    LocalMux I__10438 (
            .O(N__45658),
            .I(N__45635));
    InMux I__10437 (
            .O(N__45657),
            .I(N__45632));
    InMux I__10436 (
            .O(N__45656),
            .I(N__45629));
    InMux I__10435 (
            .O(N__45655),
            .I(N__45626));
    LocalMux I__10434 (
            .O(N__45650),
            .I(N__45621));
    LocalMux I__10433 (
            .O(N__45647),
            .I(N__45621));
    LocalMux I__10432 (
            .O(N__45644),
            .I(N__45616));
    Span4Mux_v I__10431 (
            .O(N__45641),
            .I(N__45616));
    Span4Mux_h I__10430 (
            .O(N__45638),
            .I(N__45611));
    Span4Mux_h I__10429 (
            .O(N__45635),
            .I(N__45611));
    LocalMux I__10428 (
            .O(N__45632),
            .I(N__45608));
    LocalMux I__10427 (
            .O(N__45629),
            .I(n12353));
    LocalMux I__10426 (
            .O(N__45626),
            .I(n12353));
    Odrv12 I__10425 (
            .O(N__45621),
            .I(n12353));
    Odrv4 I__10424 (
            .O(N__45616),
            .I(n12353));
    Odrv4 I__10423 (
            .O(N__45611),
            .I(n12353));
    Odrv4 I__10422 (
            .O(N__45608),
            .I(n12353));
    CascadeMux I__10421 (
            .O(N__45595),
            .I(N__45592));
    InMux I__10420 (
            .O(N__45592),
            .I(N__45588));
    InMux I__10419 (
            .O(N__45591),
            .I(N__45585));
    LocalMux I__10418 (
            .O(N__45588),
            .I(N__45582));
    LocalMux I__10417 (
            .O(N__45585),
            .I(N__45578));
    Span4Mux_v I__10416 (
            .O(N__45582),
            .I(N__45575));
    InMux I__10415 (
            .O(N__45581),
            .I(N__45572));
    Span4Mux_v I__10414 (
            .O(N__45578),
            .I(N__45567));
    Span4Mux_h I__10413 (
            .O(N__45575),
            .I(N__45567));
    LocalMux I__10412 (
            .O(N__45572),
            .I(buf_dds0_15));
    Odrv4 I__10411 (
            .O(N__45567),
            .I(buf_dds0_15));
    InMux I__10410 (
            .O(N__45562),
            .I(N__45558));
    InMux I__10409 (
            .O(N__45561),
            .I(N__45555));
    LocalMux I__10408 (
            .O(N__45558),
            .I(N__45552));
    LocalMux I__10407 (
            .O(N__45555),
            .I(N__45549));
    Span4Mux_v I__10406 (
            .O(N__45552),
            .I(N__45546));
    Span4Mux_h I__10405 (
            .O(N__45549),
            .I(N__45543));
    Odrv4 I__10404 (
            .O(N__45546),
            .I(n9));
    Odrv4 I__10403 (
            .O(N__45543),
            .I(n9));
    CEMux I__10402 (
            .O(N__45538),
            .I(N__45535));
    LocalMux I__10401 (
            .O(N__45535),
            .I(N__45531));
    CEMux I__10400 (
            .O(N__45534),
            .I(N__45528));
    Span4Mux_v I__10399 (
            .O(N__45531),
            .I(N__45525));
    LocalMux I__10398 (
            .O(N__45528),
            .I(N__45522));
    Span4Mux_h I__10397 (
            .O(N__45525),
            .I(N__45519));
    Span4Mux_h I__10396 (
            .O(N__45522),
            .I(N__45516));
    Odrv4 I__10395 (
            .O(N__45519),
            .I(\SIG_DDS.n9 ));
    Odrv4 I__10394 (
            .O(N__45516),
            .I(\SIG_DDS.n9 ));
    IoInMux I__10393 (
            .O(N__45511),
            .I(N__45507));
    InMux I__10392 (
            .O(N__45510),
            .I(N__45504));
    LocalMux I__10391 (
            .O(N__45507),
            .I(N__45501));
    LocalMux I__10390 (
            .O(N__45504),
            .I(N__45498));
    Span4Mux_s1_v I__10389 (
            .O(N__45501),
            .I(N__45494));
    Span4Mux_h I__10388 (
            .O(N__45498),
            .I(N__45491));
    InMux I__10387 (
            .O(N__45497),
            .I(N__45488));
    Span4Mux_v I__10386 (
            .O(N__45494),
            .I(N__45483));
    Span4Mux_v I__10385 (
            .O(N__45491),
            .I(N__45483));
    LocalMux I__10384 (
            .O(N__45488),
            .I(SELIRNG1));
    Odrv4 I__10383 (
            .O(N__45483),
            .I(SELIRNG1));
    InMux I__10382 (
            .O(N__45478),
            .I(N__45474));
    CascadeMux I__10381 (
            .O(N__45477),
            .I(N__45471));
    LocalMux I__10380 (
            .O(N__45474),
            .I(N__45467));
    InMux I__10379 (
            .O(N__45471),
            .I(N__45464));
    InMux I__10378 (
            .O(N__45470),
            .I(N__45461));
    Span4Mux_h I__10377 (
            .O(N__45467),
            .I(N__45456));
    LocalMux I__10376 (
            .O(N__45464),
            .I(N__45456));
    LocalMux I__10375 (
            .O(N__45461),
            .I(acadc_skipCount_11));
    Odrv4 I__10374 (
            .O(N__45456),
            .I(acadc_skipCount_11));
    InMux I__10373 (
            .O(N__45451),
            .I(N__45448));
    LocalMux I__10372 (
            .O(N__45448),
            .I(n23_adj_1518));
    InMux I__10371 (
            .O(N__45445),
            .I(N__45442));
    LocalMux I__10370 (
            .O(N__45442),
            .I(comm_length_0));
    CEMux I__10369 (
            .O(N__45439),
            .I(N__45436));
    LocalMux I__10368 (
            .O(N__45436),
            .I(N__45433));
    Span4Mux_v I__10367 (
            .O(N__45433),
            .I(N__45428));
    InMux I__10366 (
            .O(N__45432),
            .I(N__45425));
    InMux I__10365 (
            .O(N__45431),
            .I(N__45422));
    Span4Mux_h I__10364 (
            .O(N__45428),
            .I(N__45419));
    LocalMux I__10363 (
            .O(N__45425),
            .I(N__45414));
    LocalMux I__10362 (
            .O(N__45422),
            .I(N__45414));
    Span4Mux_h I__10361 (
            .O(N__45419),
            .I(N__45411));
    Span4Mux_h I__10360 (
            .O(N__45414),
            .I(N__45408));
    Odrv4 I__10359 (
            .O(N__45411),
            .I(n11846));
    Odrv4 I__10358 (
            .O(N__45408),
            .I(n11846));
    SRMux I__10357 (
            .O(N__45403),
            .I(N__45400));
    LocalMux I__10356 (
            .O(N__45400),
            .I(N__45397));
    Odrv12 I__10355 (
            .O(N__45397),
            .I(n14652));
    CascadeMux I__10354 (
            .O(N__45394),
            .I(N__45391));
    InMux I__10353 (
            .O(N__45391),
            .I(N__45388));
    LocalMux I__10352 (
            .O(N__45388),
            .I(N__45385));
    Odrv4 I__10351 (
            .O(N__45385),
            .I(n10553));
    CascadeMux I__10350 (
            .O(N__45382),
            .I(N__45377));
    CascadeMux I__10349 (
            .O(N__45381),
            .I(N__45373));
    InMux I__10348 (
            .O(N__45380),
            .I(N__45370));
    InMux I__10347 (
            .O(N__45377),
            .I(N__45367));
    InMux I__10346 (
            .O(N__45376),
            .I(N__45364));
    InMux I__10345 (
            .O(N__45373),
            .I(N__45361));
    LocalMux I__10344 (
            .O(N__45370),
            .I(N__45356));
    LocalMux I__10343 (
            .O(N__45367),
            .I(N__45356));
    LocalMux I__10342 (
            .O(N__45364),
            .I(N__45353));
    LocalMux I__10341 (
            .O(N__45361),
            .I(N__45350));
    Span4Mux_h I__10340 (
            .O(N__45356),
            .I(N__45347));
    Span12Mux_h I__10339 (
            .O(N__45353),
            .I(N__45344));
    Span4Mux_h I__10338 (
            .O(N__45350),
            .I(N__45341));
    Span4Mux_v I__10337 (
            .O(N__45347),
            .I(N__45338));
    Odrv12 I__10336 (
            .O(N__45344),
            .I(n20622));
    Odrv4 I__10335 (
            .O(N__45341),
            .I(n20622));
    Odrv4 I__10334 (
            .O(N__45338),
            .I(n20622));
    InMux I__10333 (
            .O(N__45331),
            .I(N__45324));
    InMux I__10332 (
            .O(N__45330),
            .I(N__45317));
    InMux I__10331 (
            .O(N__45329),
            .I(N__45317));
    InMux I__10330 (
            .O(N__45328),
            .I(N__45317));
    InMux I__10329 (
            .O(N__45327),
            .I(N__45314));
    LocalMux I__10328 (
            .O(N__45324),
            .I(N__45311));
    LocalMux I__10327 (
            .O(N__45317),
            .I(N__45307));
    LocalMux I__10326 (
            .O(N__45314),
            .I(N__45304));
    Span4Mux_v I__10325 (
            .O(N__45311),
            .I(N__45301));
    InMux I__10324 (
            .O(N__45310),
            .I(N__45298));
    Span4Mux_h I__10323 (
            .O(N__45307),
            .I(N__45293));
    Span4Mux_v I__10322 (
            .O(N__45304),
            .I(N__45293));
    Sp12to4 I__10321 (
            .O(N__45301),
            .I(N__45289));
    LocalMux I__10320 (
            .O(N__45298),
            .I(N__45286));
    Span4Mux_h I__10319 (
            .O(N__45293),
            .I(N__45283));
    InMux I__10318 (
            .O(N__45292),
            .I(N__45280));
    Span12Mux_h I__10317 (
            .O(N__45289),
            .I(N__45276));
    Span12Mux_v I__10316 (
            .O(N__45286),
            .I(N__45273));
    Span4Mux_h I__10315 (
            .O(N__45283),
            .I(N__45268));
    LocalMux I__10314 (
            .O(N__45280),
            .I(N__45268));
    InMux I__10313 (
            .O(N__45279),
            .I(N__45265));
    Odrv12 I__10312 (
            .O(N__45276),
            .I(n12381));
    Odrv12 I__10311 (
            .O(N__45273),
            .I(n12381));
    Odrv4 I__10310 (
            .O(N__45268),
            .I(n12381));
    LocalMux I__10309 (
            .O(N__45265),
            .I(n12381));
    CascadeMux I__10308 (
            .O(N__45256),
            .I(N__45251));
    InMux I__10307 (
            .O(N__45255),
            .I(N__45248));
    InMux I__10306 (
            .O(N__45254),
            .I(N__45245));
    InMux I__10305 (
            .O(N__45251),
            .I(N__45242));
    LocalMux I__10304 (
            .O(N__45248),
            .I(req_data_cnt_11));
    LocalMux I__10303 (
            .O(N__45245),
            .I(req_data_cnt_11));
    LocalMux I__10302 (
            .O(N__45242),
            .I(req_data_cnt_11));
    InMux I__10301 (
            .O(N__45235),
            .I(N__45232));
    LocalMux I__10300 (
            .O(N__45232),
            .I(N__45228));
    InMux I__10299 (
            .O(N__45231),
            .I(N__45224));
    Span12Mux_h I__10298 (
            .O(N__45228),
            .I(N__45221));
    InMux I__10297 (
            .O(N__45227),
            .I(N__45218));
    LocalMux I__10296 (
            .O(N__45224),
            .I(req_data_cnt_14));
    Odrv12 I__10295 (
            .O(N__45221),
            .I(req_data_cnt_14));
    LocalMux I__10294 (
            .O(N__45218),
            .I(req_data_cnt_14));
    InMux I__10293 (
            .O(N__45211),
            .I(N__45208));
    LocalMux I__10292 (
            .O(N__45208),
            .I(n23_adj_1491));
    CascadeMux I__10291 (
            .O(N__45205),
            .I(N__45202));
    InMux I__10290 (
            .O(N__45202),
            .I(N__45198));
    CascadeMux I__10289 (
            .O(N__45201),
            .I(N__45195));
    LocalMux I__10288 (
            .O(N__45198),
            .I(N__45192));
    InMux I__10287 (
            .O(N__45195),
            .I(N__45189));
    Span4Mux_v I__10286 (
            .O(N__45192),
            .I(N__45186));
    LocalMux I__10285 (
            .O(N__45189),
            .I(N__45183));
    Span4Mux_h I__10284 (
            .O(N__45186),
            .I(N__45180));
    Span4Mux_v I__10283 (
            .O(N__45183),
            .I(N__45176));
    Span4Mux_h I__10282 (
            .O(N__45180),
            .I(N__45173));
    InMux I__10281 (
            .O(N__45179),
            .I(N__45170));
    Odrv4 I__10280 (
            .O(N__45176),
            .I(cmd_rdadctmp_15_adj_1428));
    Odrv4 I__10279 (
            .O(N__45173),
            .I(cmd_rdadctmp_15_adj_1428));
    LocalMux I__10278 (
            .O(N__45170),
            .I(cmd_rdadctmp_15_adj_1428));
    CascadeMux I__10277 (
            .O(N__45163),
            .I(N__45160));
    InMux I__10276 (
            .O(N__45160),
            .I(N__45156));
    CascadeMux I__10275 (
            .O(N__45159),
            .I(N__45152));
    LocalMux I__10274 (
            .O(N__45156),
            .I(N__45149));
    InMux I__10273 (
            .O(N__45155),
            .I(N__45144));
    InMux I__10272 (
            .O(N__45152),
            .I(N__45144));
    Odrv4 I__10271 (
            .O(N__45149),
            .I(cmd_rdadctmp_15));
    LocalMux I__10270 (
            .O(N__45144),
            .I(cmd_rdadctmp_15));
    CascadeMux I__10269 (
            .O(N__45139),
            .I(N__45135));
    CascadeMux I__10268 (
            .O(N__45138),
            .I(N__45132));
    InMux I__10267 (
            .O(N__45135),
            .I(N__45129));
    InMux I__10266 (
            .O(N__45132),
            .I(N__45126));
    LocalMux I__10265 (
            .O(N__45129),
            .I(N__45123));
    LocalMux I__10264 (
            .O(N__45126),
            .I(N__45120));
    Span4Mux_h I__10263 (
            .O(N__45123),
            .I(N__45117));
    Span4Mux_v I__10262 (
            .O(N__45120),
            .I(N__45114));
    Span4Mux_h I__10261 (
            .O(N__45117),
            .I(N__45110));
    Sp12to4 I__10260 (
            .O(N__45114),
            .I(N__45107));
    InMux I__10259 (
            .O(N__45113),
            .I(N__45104));
    Span4Mux_h I__10258 (
            .O(N__45110),
            .I(N__45101));
    Span12Mux_h I__10257 (
            .O(N__45107),
            .I(N__45098));
    LocalMux I__10256 (
            .O(N__45104),
            .I(cmd_rdadctmp_16));
    Odrv4 I__10255 (
            .O(N__45101),
            .I(cmd_rdadctmp_16));
    Odrv12 I__10254 (
            .O(N__45098),
            .I(cmd_rdadctmp_16));
    CascadeMux I__10253 (
            .O(N__45091),
            .I(N__45088));
    InMux I__10252 (
            .O(N__45088),
            .I(N__45083));
    InMux I__10251 (
            .O(N__45087),
            .I(N__45080));
    InMux I__10250 (
            .O(N__45086),
            .I(N__45077));
    LocalMux I__10249 (
            .O(N__45083),
            .I(N__45074));
    LocalMux I__10248 (
            .O(N__45080),
            .I(req_data_cnt_13));
    LocalMux I__10247 (
            .O(N__45077),
            .I(req_data_cnt_13));
    Odrv4 I__10246 (
            .O(N__45074),
            .I(req_data_cnt_13));
    InMux I__10245 (
            .O(N__45067),
            .I(N__45064));
    LocalMux I__10244 (
            .O(N__45064),
            .I(N__45061));
    Odrv12 I__10243 (
            .O(N__45061),
            .I(n21022));
    CascadeMux I__10242 (
            .O(N__45058),
            .I(N__45055));
    InMux I__10241 (
            .O(N__45055),
            .I(N__45052));
    LocalMux I__10240 (
            .O(N__45052),
            .I(N__45049));
    Span4Mux_v I__10239 (
            .O(N__45049),
            .I(N__45046));
    Span4Mux_h I__10238 (
            .O(N__45046),
            .I(N__45043));
    Odrv4 I__10237 (
            .O(N__45043),
            .I(n21049));
    InMux I__10236 (
            .O(N__45040),
            .I(N__45034));
    InMux I__10235 (
            .O(N__45039),
            .I(N__45034));
    LocalMux I__10234 (
            .O(N__45034),
            .I(comm_length_2));
    CascadeMux I__10233 (
            .O(N__45031),
            .I(n21955_cascade_));
    InMux I__10232 (
            .O(N__45028),
            .I(N__45025));
    LocalMux I__10231 (
            .O(N__45025),
            .I(n21958));
    InMux I__10230 (
            .O(N__45022),
            .I(N__45019));
    LocalMux I__10229 (
            .O(N__45019),
            .I(n21024));
    InMux I__10228 (
            .O(N__45016),
            .I(N__45013));
    LocalMux I__10227 (
            .O(N__45013),
            .I(N__45010));
    Span4Mux_v I__10226 (
            .O(N__45010),
            .I(N__45007));
    Sp12to4 I__10225 (
            .O(N__45007),
            .I(N__45004));
    Span12Mux_h I__10224 (
            .O(N__45004),
            .I(N__45001));
    Odrv12 I__10223 (
            .O(N__45001),
            .I(buf_data_iac_19));
    InMux I__10222 (
            .O(N__44998),
            .I(N__44995));
    LocalMux I__10221 (
            .O(N__44995),
            .I(n20950));
    InMux I__10220 (
            .O(N__44992),
            .I(N__44989));
    LocalMux I__10219 (
            .O(N__44989),
            .I(N__44985));
    InMux I__10218 (
            .O(N__44988),
            .I(N__44982));
    Span4Mux_h I__10217 (
            .O(N__44985),
            .I(N__44979));
    LocalMux I__10216 (
            .O(N__44982),
            .I(data_idxvec_11));
    Odrv4 I__10215 (
            .O(N__44979),
            .I(data_idxvec_11));
    InMux I__10214 (
            .O(N__44974),
            .I(N__44971));
    LocalMux I__10213 (
            .O(N__44971),
            .I(n26_adj_1519));
    InMux I__10212 (
            .O(N__44968),
            .I(N__44964));
    InMux I__10211 (
            .O(N__44967),
            .I(N__44961));
    LocalMux I__10210 (
            .O(N__44964),
            .I(secclk_cnt_17));
    LocalMux I__10209 (
            .O(N__44961),
            .I(secclk_cnt_17));
    InMux I__10208 (
            .O(N__44956),
            .I(n19463));
    InMux I__10207 (
            .O(N__44953),
            .I(N__44949));
    InMux I__10206 (
            .O(N__44952),
            .I(N__44946));
    LocalMux I__10205 (
            .O(N__44949),
            .I(N__44943));
    LocalMux I__10204 (
            .O(N__44946),
            .I(secclk_cnt_18));
    Odrv4 I__10203 (
            .O(N__44943),
            .I(secclk_cnt_18));
    InMux I__10202 (
            .O(N__44938),
            .I(n19464));
    InMux I__10201 (
            .O(N__44935),
            .I(n19465));
    InMux I__10200 (
            .O(N__44932),
            .I(N__44928));
    InMux I__10199 (
            .O(N__44931),
            .I(N__44925));
    LocalMux I__10198 (
            .O(N__44928),
            .I(secclk_cnt_20));
    LocalMux I__10197 (
            .O(N__44925),
            .I(secclk_cnt_20));
    InMux I__10196 (
            .O(N__44920),
            .I(n19466));
    InMux I__10195 (
            .O(N__44917),
            .I(n19467));
    InMux I__10194 (
            .O(N__44914),
            .I(n19468));
    SRMux I__10193 (
            .O(N__44911),
            .I(N__44907));
    SRMux I__10192 (
            .O(N__44910),
            .I(N__44903));
    LocalMux I__10191 (
            .O(N__44907),
            .I(N__44899));
    SRMux I__10190 (
            .O(N__44906),
            .I(N__44896));
    LocalMux I__10189 (
            .O(N__44903),
            .I(N__44893));
    InMux I__10188 (
            .O(N__44902),
            .I(N__44890));
    Span4Mux_v I__10187 (
            .O(N__44899),
            .I(N__44887));
    LocalMux I__10186 (
            .O(N__44896),
            .I(N__44884));
    Span4Mux_h I__10185 (
            .O(N__44893),
            .I(N__44879));
    LocalMux I__10184 (
            .O(N__44890),
            .I(N__44879));
    Odrv4 I__10183 (
            .O(N__44887),
            .I(n14700));
    Odrv4 I__10182 (
            .O(N__44884),
            .I(n14700));
    Odrv4 I__10181 (
            .O(N__44879),
            .I(n14700));
    InMux I__10180 (
            .O(N__44872),
            .I(N__44868));
    InMux I__10179 (
            .O(N__44871),
            .I(N__44865));
    LocalMux I__10178 (
            .O(N__44868),
            .I(N__44862));
    LocalMux I__10177 (
            .O(N__44865),
            .I(N__44857));
    Span4Mux_h I__10176 (
            .O(N__44862),
            .I(N__44857));
    Span4Mux_h I__10175 (
            .O(N__44857),
            .I(N__44854));
    Odrv4 I__10174 (
            .O(N__44854),
            .I(comm_buf_0_5));
    CascadeMux I__10173 (
            .O(N__44851),
            .I(N__44843));
    InMux I__10172 (
            .O(N__44850),
            .I(N__44840));
    InMux I__10171 (
            .O(N__44849),
            .I(N__44837));
    InMux I__10170 (
            .O(N__44848),
            .I(N__44834));
    InMux I__10169 (
            .O(N__44847),
            .I(N__44831));
    InMux I__10168 (
            .O(N__44846),
            .I(N__44828));
    InMux I__10167 (
            .O(N__44843),
            .I(N__44825));
    LocalMux I__10166 (
            .O(N__44840),
            .I(N__44822));
    LocalMux I__10165 (
            .O(N__44837),
            .I(N__44819));
    LocalMux I__10164 (
            .O(N__44834),
            .I(N__44812));
    LocalMux I__10163 (
            .O(N__44831),
            .I(N__44812));
    LocalMux I__10162 (
            .O(N__44828),
            .I(N__44812));
    LocalMux I__10161 (
            .O(N__44825),
            .I(N__44809));
    Span4Mux_h I__10160 (
            .O(N__44822),
            .I(N__44806));
    Span4Mux_v I__10159 (
            .O(N__44819),
            .I(N__44801));
    Span4Mux_h I__10158 (
            .O(N__44812),
            .I(N__44801));
    Span4Mux_v I__10157 (
            .O(N__44809),
            .I(N__44796));
    Sp12to4 I__10156 (
            .O(N__44806),
            .I(N__44793));
    Span4Mux_h I__10155 (
            .O(N__44801),
            .I(N__44790));
    InMux I__10154 (
            .O(N__44800),
            .I(N__44785));
    InMux I__10153 (
            .O(N__44799),
            .I(N__44785));
    Span4Mux_h I__10152 (
            .O(N__44796),
            .I(N__44782));
    Span12Mux_v I__10151 (
            .O(N__44793),
            .I(N__44779));
    Span4Mux_v I__10150 (
            .O(N__44790),
            .I(N__44776));
    LocalMux I__10149 (
            .O(N__44785),
            .I(n14_adj_1556));
    Odrv4 I__10148 (
            .O(N__44782),
            .I(n14_adj_1556));
    Odrv12 I__10147 (
            .O(N__44779),
            .I(n14_adj_1556));
    Odrv4 I__10146 (
            .O(N__44776),
            .I(n14_adj_1556));
    IoInMux I__10145 (
            .O(N__44767),
            .I(N__44764));
    LocalMux I__10144 (
            .O(N__44764),
            .I(N__44761));
    IoSpan4Mux I__10143 (
            .O(N__44761),
            .I(N__44758));
    Span4Mux_s1_h I__10142 (
            .O(N__44758),
            .I(N__44755));
    Sp12to4 I__10141 (
            .O(N__44755),
            .I(N__44751));
    InMux I__10140 (
            .O(N__44754),
            .I(N__44748));
    Span12Mux_v I__10139 (
            .O(N__44751),
            .I(N__44745));
    LocalMux I__10138 (
            .O(N__44748),
            .I(N__44741));
    Span12Mux_h I__10137 (
            .O(N__44745),
            .I(N__44738));
    InMux I__10136 (
            .O(N__44744),
            .I(N__44735));
    Span4Mux_h I__10135 (
            .O(N__44741),
            .I(N__44732));
    Odrv12 I__10134 (
            .O(N__44738),
            .I(VDC_RNG0));
    LocalMux I__10133 (
            .O(N__44735),
            .I(VDC_RNG0));
    Odrv4 I__10132 (
            .O(N__44732),
            .I(VDC_RNG0));
    InMux I__10131 (
            .O(N__44725),
            .I(N__44722));
    LocalMux I__10130 (
            .O(N__44722),
            .I(N__44719));
    Span4Mux_h I__10129 (
            .O(N__44719),
            .I(N__44714));
    InMux I__10128 (
            .O(N__44718),
            .I(N__44709));
    InMux I__10127 (
            .O(N__44717),
            .I(N__44709));
    Odrv4 I__10126 (
            .O(N__44714),
            .I(acadc_skipCount_12));
    LocalMux I__10125 (
            .O(N__44709),
            .I(acadc_skipCount_12));
    InMux I__10124 (
            .O(N__44704),
            .I(N__44700));
    InMux I__10123 (
            .O(N__44703),
            .I(N__44697));
    LocalMux I__10122 (
            .O(N__44700),
            .I(secclk_cnt_9));
    LocalMux I__10121 (
            .O(N__44697),
            .I(secclk_cnt_9));
    InMux I__10120 (
            .O(N__44692),
            .I(n19455));
    CascadeMux I__10119 (
            .O(N__44689),
            .I(N__44685));
    InMux I__10118 (
            .O(N__44688),
            .I(N__44682));
    InMux I__10117 (
            .O(N__44685),
            .I(N__44679));
    LocalMux I__10116 (
            .O(N__44682),
            .I(secclk_cnt_10));
    LocalMux I__10115 (
            .O(N__44679),
            .I(secclk_cnt_10));
    InMux I__10114 (
            .O(N__44674),
            .I(n19456));
    CascadeMux I__10113 (
            .O(N__44671),
            .I(N__44667));
    InMux I__10112 (
            .O(N__44670),
            .I(N__44664));
    InMux I__10111 (
            .O(N__44667),
            .I(N__44661));
    LocalMux I__10110 (
            .O(N__44664),
            .I(secclk_cnt_11));
    LocalMux I__10109 (
            .O(N__44661),
            .I(secclk_cnt_11));
    InMux I__10108 (
            .O(N__44656),
            .I(n19457));
    InMux I__10107 (
            .O(N__44653),
            .I(n19458));
    CascadeMux I__10106 (
            .O(N__44650),
            .I(N__44646));
    InMux I__10105 (
            .O(N__44649),
            .I(N__44643));
    InMux I__10104 (
            .O(N__44646),
            .I(N__44640));
    LocalMux I__10103 (
            .O(N__44643),
            .I(secclk_cnt_13));
    LocalMux I__10102 (
            .O(N__44640),
            .I(secclk_cnt_13));
    InMux I__10101 (
            .O(N__44635),
            .I(n19459));
    InMux I__10100 (
            .O(N__44632),
            .I(N__44628));
    InMux I__10099 (
            .O(N__44631),
            .I(N__44625));
    LocalMux I__10098 (
            .O(N__44628),
            .I(secclk_cnt_14));
    LocalMux I__10097 (
            .O(N__44625),
            .I(secclk_cnt_14));
    InMux I__10096 (
            .O(N__44620),
            .I(n19460));
    InMux I__10095 (
            .O(N__44617),
            .I(N__44613));
    InMux I__10094 (
            .O(N__44616),
            .I(N__44610));
    LocalMux I__10093 (
            .O(N__44613),
            .I(secclk_cnt_15));
    LocalMux I__10092 (
            .O(N__44610),
            .I(secclk_cnt_15));
    InMux I__10091 (
            .O(N__44605),
            .I(n19461));
    InMux I__10090 (
            .O(N__44602),
            .I(N__44598));
    InMux I__10089 (
            .O(N__44601),
            .I(N__44595));
    LocalMux I__10088 (
            .O(N__44598),
            .I(secclk_cnt_16));
    LocalMux I__10087 (
            .O(N__44595),
            .I(secclk_cnt_16));
    InMux I__10086 (
            .O(N__44590),
            .I(bfn_17_11_0_));
    InMux I__10085 (
            .O(N__44587),
            .I(N__44583));
    InMux I__10084 (
            .O(N__44586),
            .I(N__44580));
    LocalMux I__10083 (
            .O(N__44583),
            .I(secclk_cnt_0));
    LocalMux I__10082 (
            .O(N__44580),
            .I(secclk_cnt_0));
    InMux I__10081 (
            .O(N__44575),
            .I(bfn_17_9_0_));
    CascadeMux I__10080 (
            .O(N__44572),
            .I(N__44568));
    InMux I__10079 (
            .O(N__44571),
            .I(N__44565));
    InMux I__10078 (
            .O(N__44568),
            .I(N__44562));
    LocalMux I__10077 (
            .O(N__44565),
            .I(secclk_cnt_1));
    LocalMux I__10076 (
            .O(N__44562),
            .I(secclk_cnt_1));
    InMux I__10075 (
            .O(N__44557),
            .I(n19447));
    InMux I__10074 (
            .O(N__44554),
            .I(N__44550));
    InMux I__10073 (
            .O(N__44553),
            .I(N__44547));
    LocalMux I__10072 (
            .O(N__44550),
            .I(secclk_cnt_2));
    LocalMux I__10071 (
            .O(N__44547),
            .I(secclk_cnt_2));
    InMux I__10070 (
            .O(N__44542),
            .I(n19448));
    InMux I__10069 (
            .O(N__44539),
            .I(N__44536));
    LocalMux I__10068 (
            .O(N__44536),
            .I(N__44532));
    InMux I__10067 (
            .O(N__44535),
            .I(N__44529));
    Odrv4 I__10066 (
            .O(N__44532),
            .I(secclk_cnt_3));
    LocalMux I__10065 (
            .O(N__44529),
            .I(secclk_cnt_3));
    InMux I__10064 (
            .O(N__44524),
            .I(n19449));
    InMux I__10063 (
            .O(N__44521),
            .I(N__44517));
    InMux I__10062 (
            .O(N__44520),
            .I(N__44514));
    LocalMux I__10061 (
            .O(N__44517),
            .I(secclk_cnt_4));
    LocalMux I__10060 (
            .O(N__44514),
            .I(secclk_cnt_4));
    InMux I__10059 (
            .O(N__44509),
            .I(n19450));
    InMux I__10058 (
            .O(N__44506),
            .I(N__44502));
    InMux I__10057 (
            .O(N__44505),
            .I(N__44499));
    LocalMux I__10056 (
            .O(N__44502),
            .I(N__44496));
    LocalMux I__10055 (
            .O(N__44499),
            .I(secclk_cnt_5));
    Odrv4 I__10054 (
            .O(N__44496),
            .I(secclk_cnt_5));
    InMux I__10053 (
            .O(N__44491),
            .I(n19451));
    InMux I__10052 (
            .O(N__44488),
            .I(N__44484));
    InMux I__10051 (
            .O(N__44487),
            .I(N__44481));
    LocalMux I__10050 (
            .O(N__44484),
            .I(secclk_cnt_6));
    LocalMux I__10049 (
            .O(N__44481),
            .I(secclk_cnt_6));
    InMux I__10048 (
            .O(N__44476),
            .I(n19452));
    InMux I__10047 (
            .O(N__44473),
            .I(N__44469));
    InMux I__10046 (
            .O(N__44472),
            .I(N__44466));
    LocalMux I__10045 (
            .O(N__44469),
            .I(N__44463));
    LocalMux I__10044 (
            .O(N__44466),
            .I(secclk_cnt_7));
    Odrv4 I__10043 (
            .O(N__44463),
            .I(secclk_cnt_7));
    InMux I__10042 (
            .O(N__44458),
            .I(n19453));
    InMux I__10041 (
            .O(N__44455),
            .I(N__44451));
    InMux I__10040 (
            .O(N__44454),
            .I(N__44448));
    LocalMux I__10039 (
            .O(N__44451),
            .I(secclk_cnt_8));
    LocalMux I__10038 (
            .O(N__44448),
            .I(secclk_cnt_8));
    InMux I__10037 (
            .O(N__44443),
            .I(bfn_17_10_0_));
    InMux I__10036 (
            .O(N__44440),
            .I(N__44437));
    LocalMux I__10035 (
            .O(N__44437),
            .I(comm_state_3_N_412_3));
    InMux I__10034 (
            .O(N__44434),
            .I(N__44431));
    LocalMux I__10033 (
            .O(N__44431),
            .I(n1252));
    InMux I__10032 (
            .O(N__44428),
            .I(N__44425));
    LocalMux I__10031 (
            .O(N__44425),
            .I(n8_adj_1555));
    CascadeMux I__10030 (
            .O(N__44422),
            .I(n2342_cascade_));
    InMux I__10029 (
            .O(N__44419),
            .I(N__44415));
    InMux I__10028 (
            .O(N__44418),
            .I(N__44412));
    LocalMux I__10027 (
            .O(N__44415),
            .I(N__44408));
    LocalMux I__10026 (
            .O(N__44412),
            .I(N__44405));
    InMux I__10025 (
            .O(N__44411),
            .I(N__44402));
    Span4Mux_v I__10024 (
            .O(N__44408),
            .I(N__44397));
    Span12Mux_v I__10023 (
            .O(N__44405),
            .I(N__44392));
    LocalMux I__10022 (
            .O(N__44402),
            .I(N__44392));
    InMux I__10021 (
            .O(N__44401),
            .I(N__44389));
    InMux I__10020 (
            .O(N__44400),
            .I(N__44386));
    Sp12to4 I__10019 (
            .O(N__44397),
            .I(N__44379));
    Span12Mux_v I__10018 (
            .O(N__44392),
            .I(N__44379));
    LocalMux I__10017 (
            .O(N__44389),
            .I(N__44379));
    LocalMux I__10016 (
            .O(N__44386),
            .I(comm_state_3_N_428_2));
    Odrv12 I__10015 (
            .O(N__44379),
            .I(comm_state_3_N_428_2));
    CascadeMux I__10014 (
            .O(N__44374),
            .I(n15_adj_1602_cascade_));
    InMux I__10013 (
            .O(N__44371),
            .I(N__44368));
    LocalMux I__10012 (
            .O(N__44368),
            .I(n20571));
    CascadeMux I__10011 (
            .O(N__44365),
            .I(n20641_cascade_));
    InMux I__10010 (
            .O(N__44362),
            .I(N__44359));
    LocalMux I__10009 (
            .O(N__44359),
            .I(n12_adj_1603));
    InMux I__10008 (
            .O(N__44356),
            .I(N__44353));
    LocalMux I__10007 (
            .O(N__44353),
            .I(N__44350));
    Span4Mux_h I__10006 (
            .O(N__44350),
            .I(N__44347));
    Span4Mux_h I__10005 (
            .O(N__44347),
            .I(N__44344));
    Odrv4 I__10004 (
            .O(N__44344),
            .I(n7_adj_1588));
    SRMux I__10003 (
            .O(N__44341),
            .I(N__44338));
    LocalMux I__10002 (
            .O(N__44338),
            .I(N__44335));
    Span4Mux_v I__10001 (
            .O(N__44335),
            .I(N__44332));
    Span4Mux_h I__10000 (
            .O(N__44332),
            .I(N__44329));
    Span4Mux_v I__9999 (
            .O(N__44329),
            .I(N__44326));
    Odrv4 I__9998 (
            .O(N__44326),
            .I(\comm_spi.data_tx_7__N_759 ));
    InMux I__9997 (
            .O(N__44323),
            .I(N__44319));
    InMux I__9996 (
            .O(N__44322),
            .I(N__44316));
    LocalMux I__9995 (
            .O(N__44319),
            .I(\comm_spi.n14596 ));
    LocalMux I__9994 (
            .O(N__44316),
            .I(\comm_spi.n14596 ));
    InMux I__9993 (
            .O(N__44311),
            .I(N__44307));
    InMux I__9992 (
            .O(N__44310),
            .I(N__44304));
    LocalMux I__9991 (
            .O(N__44307),
            .I(N__44301));
    LocalMux I__9990 (
            .O(N__44304),
            .I(N__44298));
    Span4Mux_v I__9989 (
            .O(N__44301),
            .I(N__44295));
    Span4Mux_v I__9988 (
            .O(N__44298),
            .I(N__44292));
    Odrv4 I__9987 (
            .O(N__44295),
            .I(\comm_spi.n14595 ));
    Odrv4 I__9986 (
            .O(N__44292),
            .I(\comm_spi.n14595 ));
    InMux I__9985 (
            .O(N__44287),
            .I(N__44284));
    LocalMux I__9984 (
            .O(N__44284),
            .I(N__44279));
    InMux I__9983 (
            .O(N__44283),
            .I(N__44276));
    InMux I__9982 (
            .O(N__44282),
            .I(N__44273));
    Span4Mux_v I__9981 (
            .O(N__44279),
            .I(N__44263));
    LocalMux I__9980 (
            .O(N__44276),
            .I(N__44263));
    LocalMux I__9979 (
            .O(N__44273),
            .I(N__44263));
    InMux I__9978 (
            .O(N__44272),
            .I(N__44260));
    InMux I__9977 (
            .O(N__44271),
            .I(N__44257));
    InMux I__9976 (
            .O(N__44270),
            .I(N__44254));
    Span4Mux_h I__9975 (
            .O(N__44263),
            .I(N__44251));
    LocalMux I__9974 (
            .O(N__44260),
            .I(\comm_spi.n14588 ));
    LocalMux I__9973 (
            .O(N__44257),
            .I(\comm_spi.n14588 ));
    LocalMux I__9972 (
            .O(N__44254),
            .I(\comm_spi.n14588 ));
    Odrv4 I__9971 (
            .O(N__44251),
            .I(\comm_spi.n14588 ));
    InMux I__9970 (
            .O(N__44242),
            .I(N__44239));
    LocalMux I__9969 (
            .O(N__44239),
            .I(N__44236));
    Odrv4 I__9968 (
            .O(N__44236),
            .I(\comm_spi.n14590 ));
    SRMux I__9967 (
            .O(N__44233),
            .I(N__44228));
    SRMux I__9966 (
            .O(N__44232),
            .I(N__44225));
    SRMux I__9965 (
            .O(N__44231),
            .I(N__44222));
    LocalMux I__9964 (
            .O(N__44228),
            .I(N__44219));
    LocalMux I__9963 (
            .O(N__44225),
            .I(N__44216));
    LocalMux I__9962 (
            .O(N__44222),
            .I(N__44213));
    Span4Mux_h I__9961 (
            .O(N__44219),
            .I(N__44210));
    Span4Mux_v I__9960 (
            .O(N__44216),
            .I(N__44207));
    Span4Mux_v I__9959 (
            .O(N__44213),
            .I(N__44204));
    Odrv4 I__9958 (
            .O(N__44210),
            .I(\comm_spi.data_tx_7__N_766 ));
    Odrv4 I__9957 (
            .O(N__44207),
            .I(\comm_spi.data_tx_7__N_766 ));
    Odrv4 I__9956 (
            .O(N__44204),
            .I(\comm_spi.data_tx_7__N_766 ));
    InMux I__9955 (
            .O(N__44197),
            .I(N__44194));
    LocalMux I__9954 (
            .O(N__44194),
            .I(N__44191));
    Span4Mux_h I__9953 (
            .O(N__44191),
            .I(N__44188));
    Span4Mux_h I__9952 (
            .O(N__44188),
            .I(N__44185));
    Odrv4 I__9951 (
            .O(N__44185),
            .I(n20931));
    CascadeMux I__9950 (
            .O(N__44182),
            .I(n21913_cascade_));
    InMux I__9949 (
            .O(N__44179),
            .I(N__44176));
    LocalMux I__9948 (
            .O(N__44176),
            .I(n21916));
    CascadeMux I__9947 (
            .O(N__44173),
            .I(n1252_cascade_));
    InMux I__9946 (
            .O(N__44170),
            .I(N__44167));
    LocalMux I__9945 (
            .O(N__44167),
            .I(n2));
    CascadeMux I__9944 (
            .O(N__44164),
            .I(n21088_cascade_));
    CEMux I__9943 (
            .O(N__44161),
            .I(N__44158));
    LocalMux I__9942 (
            .O(N__44158),
            .I(N__44155));
    Span4Mux_v I__9941 (
            .O(N__44155),
            .I(N__44152));
    Odrv4 I__9940 (
            .O(N__44152),
            .I(n14_adj_1497));
    CascadeMux I__9939 (
            .O(N__44149),
            .I(N__44143));
    CascadeMux I__9938 (
            .O(N__44148),
            .I(N__44140));
    CascadeMux I__9937 (
            .O(N__44147),
            .I(N__44137));
    CascadeMux I__9936 (
            .O(N__44146),
            .I(N__44134));
    InMux I__9935 (
            .O(N__44143),
            .I(N__44131));
    InMux I__9934 (
            .O(N__44140),
            .I(N__44128));
    InMux I__9933 (
            .O(N__44137),
            .I(N__44124));
    InMux I__9932 (
            .O(N__44134),
            .I(N__44121));
    LocalMux I__9931 (
            .O(N__44131),
            .I(N__44116));
    LocalMux I__9930 (
            .O(N__44128),
            .I(N__44116));
    InMux I__9929 (
            .O(N__44127),
            .I(N__44113));
    LocalMux I__9928 (
            .O(N__44124),
            .I(N__44109));
    LocalMux I__9927 (
            .O(N__44121),
            .I(N__44104));
    Span4Mux_v I__9926 (
            .O(N__44116),
            .I(N__44101));
    LocalMux I__9925 (
            .O(N__44113),
            .I(N__44098));
    InMux I__9924 (
            .O(N__44112),
            .I(N__44095));
    Span4Mux_v I__9923 (
            .O(N__44109),
            .I(N__44092));
    InMux I__9922 (
            .O(N__44108),
            .I(N__44089));
    InMux I__9921 (
            .O(N__44107),
            .I(N__44086));
    Span4Mux_v I__9920 (
            .O(N__44104),
            .I(N__44081));
    Span4Mux_h I__9919 (
            .O(N__44101),
            .I(N__44076));
    Span4Mux_v I__9918 (
            .O(N__44098),
            .I(N__44076));
    LocalMux I__9917 (
            .O(N__44095),
            .I(N__44073));
    Span4Mux_h I__9916 (
            .O(N__44092),
            .I(N__44066));
    LocalMux I__9915 (
            .O(N__44089),
            .I(N__44066));
    LocalMux I__9914 (
            .O(N__44086),
            .I(N__44066));
    InMux I__9913 (
            .O(N__44085),
            .I(N__44061));
    InMux I__9912 (
            .O(N__44084),
            .I(N__44061));
    Sp12to4 I__9911 (
            .O(N__44081),
            .I(N__44058));
    Span4Mux_v I__9910 (
            .O(N__44076),
            .I(N__44053));
    Span4Mux_v I__9909 (
            .O(N__44073),
            .I(N__44053));
    Span4Mux_v I__9908 (
            .O(N__44066),
            .I(N__44050));
    LocalMux I__9907 (
            .O(N__44061),
            .I(N__44047));
    Span12Mux_v I__9906 (
            .O(N__44058),
            .I(N__44040));
    Sp12to4 I__9905 (
            .O(N__44053),
            .I(N__44040));
    Sp12to4 I__9904 (
            .O(N__44050),
            .I(N__44040));
    Odrv4 I__9903 (
            .O(N__44047),
            .I(comm_buf_0_1));
    Odrv12 I__9902 (
            .O(N__44040),
            .I(comm_buf_0_1));
    IoInMux I__9901 (
            .O(N__44035),
            .I(N__44032));
    LocalMux I__9900 (
            .O(N__44032),
            .I(N__44028));
    InMux I__9899 (
            .O(N__44031),
            .I(N__44025));
    IoSpan4Mux I__9898 (
            .O(N__44028),
            .I(N__44022));
    LocalMux I__9897 (
            .O(N__44025),
            .I(N__44019));
    IoSpan4Mux I__9896 (
            .O(N__44022),
            .I(N__44016));
    Span4Mux_h I__9895 (
            .O(N__44019),
            .I(N__44013));
    Span4Mux_s3_v I__9894 (
            .O(N__44016),
            .I(N__44010));
    Span4Mux_v I__9893 (
            .O(N__44013),
            .I(N__44006));
    Span4Mux_v I__9892 (
            .O(N__44010),
            .I(N__44003));
    InMux I__9891 (
            .O(N__44009),
            .I(N__44000));
    Span4Mux_h I__9890 (
            .O(N__44006),
            .I(N__43997));
    Odrv4 I__9889 (
            .O(N__44003),
            .I(DDS_RNG_0));
    LocalMux I__9888 (
            .O(N__44000),
            .I(DDS_RNG_0));
    Odrv4 I__9887 (
            .O(N__43997),
            .I(DDS_RNG_0));
    InMux I__9886 (
            .O(N__43990),
            .I(N__43987));
    LocalMux I__9885 (
            .O(N__43987),
            .I(N__43984));
    Odrv4 I__9884 (
            .O(N__43984),
            .I(n8_adj_1538));
    InMux I__9883 (
            .O(N__43981),
            .I(N__43977));
    InMux I__9882 (
            .O(N__43980),
            .I(N__43974));
    LocalMux I__9881 (
            .O(N__43977),
            .I(N__43969));
    LocalMux I__9880 (
            .O(N__43974),
            .I(N__43969));
    Odrv12 I__9879 (
            .O(N__43969),
            .I(n7_adj_1537));
    CascadeMux I__9878 (
            .O(N__43966),
            .I(N__43963));
    CascadeBuf I__9877 (
            .O(N__43963),
            .I(N__43960));
    CascadeMux I__9876 (
            .O(N__43960),
            .I(N__43957));
    CascadeBuf I__9875 (
            .O(N__43957),
            .I(N__43954));
    CascadeMux I__9874 (
            .O(N__43954),
            .I(N__43951));
    CascadeBuf I__9873 (
            .O(N__43951),
            .I(N__43948));
    CascadeMux I__9872 (
            .O(N__43948),
            .I(N__43945));
    CascadeBuf I__9871 (
            .O(N__43945),
            .I(N__43942));
    CascadeMux I__9870 (
            .O(N__43942),
            .I(N__43939));
    CascadeBuf I__9869 (
            .O(N__43939),
            .I(N__43936));
    CascadeMux I__9868 (
            .O(N__43936),
            .I(N__43933));
    CascadeBuf I__9867 (
            .O(N__43933),
            .I(N__43930));
    CascadeMux I__9866 (
            .O(N__43930),
            .I(N__43927));
    CascadeBuf I__9865 (
            .O(N__43927),
            .I(N__43924));
    CascadeMux I__9864 (
            .O(N__43924),
            .I(N__43920));
    CascadeMux I__9863 (
            .O(N__43923),
            .I(N__43917));
    CascadeBuf I__9862 (
            .O(N__43920),
            .I(N__43914));
    CascadeBuf I__9861 (
            .O(N__43917),
            .I(N__43911));
    CascadeMux I__9860 (
            .O(N__43914),
            .I(N__43908));
    CascadeMux I__9859 (
            .O(N__43911),
            .I(N__43905));
    CascadeBuf I__9858 (
            .O(N__43908),
            .I(N__43902));
    InMux I__9857 (
            .O(N__43905),
            .I(N__43899));
    CascadeMux I__9856 (
            .O(N__43902),
            .I(N__43896));
    LocalMux I__9855 (
            .O(N__43899),
            .I(N__43893));
    InMux I__9854 (
            .O(N__43896),
            .I(N__43890));
    Span4Mux_v I__9853 (
            .O(N__43893),
            .I(N__43887));
    LocalMux I__9852 (
            .O(N__43890),
            .I(N__43884));
    Span4Mux_h I__9851 (
            .O(N__43887),
            .I(N__43881));
    Span12Mux_h I__9850 (
            .O(N__43884),
            .I(N__43878));
    Odrv4 I__9849 (
            .O(N__43881),
            .I(data_index_9_N_212_6));
    Odrv12 I__9848 (
            .O(N__43878),
            .I(data_index_9_N_212_6));
    InMux I__9847 (
            .O(N__43873),
            .I(N__43866));
    InMux I__9846 (
            .O(N__43872),
            .I(N__43866));
    InMux I__9845 (
            .O(N__43871),
            .I(N__43861));
    LocalMux I__9844 (
            .O(N__43866),
            .I(N__43858));
    InMux I__9843 (
            .O(N__43865),
            .I(N__43855));
    InMux I__9842 (
            .O(N__43864),
            .I(N__43852));
    LocalMux I__9841 (
            .O(N__43861),
            .I(N__43849));
    Span4Mux_v I__9840 (
            .O(N__43858),
            .I(N__43842));
    LocalMux I__9839 (
            .O(N__43855),
            .I(N__43842));
    LocalMux I__9838 (
            .O(N__43852),
            .I(N__43837));
    Span4Mux_h I__9837 (
            .O(N__43849),
            .I(N__43837));
    InMux I__9836 (
            .O(N__43848),
            .I(N__43834));
    InMux I__9835 (
            .O(N__43847),
            .I(N__43831));
    Odrv4 I__9834 (
            .O(N__43842),
            .I(n11901));
    Odrv4 I__9833 (
            .O(N__43837),
            .I(n11901));
    LocalMux I__9832 (
            .O(N__43834),
            .I(n11901));
    LocalMux I__9831 (
            .O(N__43831),
            .I(n11901));
    CascadeMux I__9830 (
            .O(N__43822),
            .I(N__43818));
    InMux I__9829 (
            .O(N__43821),
            .I(N__43813));
    InMux I__9828 (
            .O(N__43818),
            .I(N__43810));
    InMux I__9827 (
            .O(N__43817),
            .I(N__43807));
    CascadeMux I__9826 (
            .O(N__43816),
            .I(N__43803));
    LocalMux I__9825 (
            .O(N__43813),
            .I(N__43797));
    LocalMux I__9824 (
            .O(N__43810),
            .I(N__43797));
    LocalMux I__9823 (
            .O(N__43807),
            .I(N__43793));
    CascadeMux I__9822 (
            .O(N__43806),
            .I(N__43790));
    InMux I__9821 (
            .O(N__43803),
            .I(N__43787));
    InMux I__9820 (
            .O(N__43802),
            .I(N__43784));
    Span4Mux_v I__9819 (
            .O(N__43797),
            .I(N__43781));
    InMux I__9818 (
            .O(N__43796),
            .I(N__43778));
    Span4Mux_h I__9817 (
            .O(N__43793),
            .I(N__43775));
    InMux I__9816 (
            .O(N__43790),
            .I(N__43772));
    LocalMux I__9815 (
            .O(N__43787),
            .I(N__43769));
    LocalMux I__9814 (
            .O(N__43784),
            .I(N__43761));
    Span4Mux_v I__9813 (
            .O(N__43781),
            .I(N__43761));
    LocalMux I__9812 (
            .O(N__43778),
            .I(N__43761));
    Span4Mux_v I__9811 (
            .O(N__43775),
            .I(N__43755));
    LocalMux I__9810 (
            .O(N__43772),
            .I(N__43755));
    Span4Mux_h I__9809 (
            .O(N__43769),
            .I(N__43752));
    InMux I__9808 (
            .O(N__43768),
            .I(N__43749));
    Span4Mux_h I__9807 (
            .O(N__43761),
            .I(N__43746));
    CascadeMux I__9806 (
            .O(N__43760),
            .I(N__43743));
    Span4Mux_h I__9805 (
            .O(N__43755),
            .I(N__43740));
    Span4Mux_v I__9804 (
            .O(N__43752),
            .I(N__43735));
    LocalMux I__9803 (
            .O(N__43749),
            .I(N__43735));
    Span4Mux_h I__9802 (
            .O(N__43746),
            .I(N__43732));
    InMux I__9801 (
            .O(N__43743),
            .I(N__43729));
    Span4Mux_h I__9800 (
            .O(N__43740),
            .I(N__43726));
    Span4Mux_h I__9799 (
            .O(N__43735),
            .I(N__43723));
    Sp12to4 I__9798 (
            .O(N__43732),
            .I(N__43720));
    LocalMux I__9797 (
            .O(N__43729),
            .I(comm_buf_0_3));
    Odrv4 I__9796 (
            .O(N__43726),
            .I(comm_buf_0_3));
    Odrv4 I__9795 (
            .O(N__43723),
            .I(comm_buf_0_3));
    Odrv12 I__9794 (
            .O(N__43720),
            .I(comm_buf_0_3));
    SRMux I__9793 (
            .O(N__43711),
            .I(N__43707));
    InMux I__9792 (
            .O(N__43710),
            .I(N__43704));
    LocalMux I__9791 (
            .O(N__43707),
            .I(N__43701));
    LocalMux I__9790 (
            .O(N__43704),
            .I(N__43698));
    Span4Mux_h I__9789 (
            .O(N__43701),
            .I(N__43695));
    Span4Mux_v I__9788 (
            .O(N__43698),
            .I(N__43692));
    Odrv4 I__9787 (
            .O(N__43695),
            .I(n14869));
    Odrv4 I__9786 (
            .O(N__43692),
            .I(n14869));
    InMux I__9785 (
            .O(N__43687),
            .I(N__43678));
    InMux I__9784 (
            .O(N__43686),
            .I(N__43678));
    InMux I__9783 (
            .O(N__43685),
            .I(N__43678));
    LocalMux I__9782 (
            .O(N__43678),
            .I(N__43674));
    InMux I__9781 (
            .O(N__43677),
            .I(N__43670));
    Span4Mux_h I__9780 (
            .O(N__43674),
            .I(N__43667));
    CascadeMux I__9779 (
            .O(N__43673),
            .I(N__43664));
    LocalMux I__9778 (
            .O(N__43670),
            .I(N__43661));
    Span4Mux_v I__9777 (
            .O(N__43667),
            .I(N__43658));
    InMux I__9776 (
            .O(N__43664),
            .I(N__43655));
    Span12Mux_h I__9775 (
            .O(N__43661),
            .I(N__43652));
    Odrv4 I__9774 (
            .O(N__43658),
            .I(bit_cnt_0));
    LocalMux I__9773 (
            .O(N__43655),
            .I(bit_cnt_0));
    Odrv12 I__9772 (
            .O(N__43652),
            .I(bit_cnt_0));
    InMux I__9771 (
            .O(N__43645),
            .I(N__43642));
    LocalMux I__9770 (
            .O(N__43642),
            .I(N__43638));
    InMux I__9769 (
            .O(N__43641),
            .I(N__43635));
    Odrv4 I__9768 (
            .O(N__43638),
            .I(\comm_spi.n14624 ));
    LocalMux I__9767 (
            .O(N__43635),
            .I(\comm_spi.n14624 ));
    SRMux I__9766 (
            .O(N__43630),
            .I(N__43627));
    LocalMux I__9765 (
            .O(N__43627),
            .I(N__43624));
    Span4Mux_v I__9764 (
            .O(N__43624),
            .I(N__43621));
    Span4Mux_h I__9763 (
            .O(N__43621),
            .I(N__43618));
    Span4Mux_v I__9762 (
            .O(N__43618),
            .I(N__43615));
    Odrv4 I__9761 (
            .O(N__43615),
            .I(\comm_spi.data_tx_7__N_769 ));
    InMux I__9760 (
            .O(N__43612),
            .I(N__43609));
    LocalMux I__9759 (
            .O(N__43609),
            .I(\comm_spi.n22626 ));
    CascadeMux I__9758 (
            .O(N__43606),
            .I(\comm_spi.n22626_cascade_ ));
    InMux I__9757 (
            .O(N__43603),
            .I(N__43600));
    LocalMux I__9756 (
            .O(N__43600),
            .I(N__43597));
    Span4Mux_v I__9755 (
            .O(N__43597),
            .I(N__43594));
    Odrv4 I__9754 (
            .O(N__43594),
            .I(\comm_spi.n14589 ));
    IoInMux I__9753 (
            .O(N__43591),
            .I(N__43588));
    LocalMux I__9752 (
            .O(N__43588),
            .I(N__43585));
    Span4Mux_s1_h I__9751 (
            .O(N__43585),
            .I(N__43582));
    Sp12to4 I__9750 (
            .O(N__43582),
            .I(N__43579));
    Span12Mux_s9_v I__9749 (
            .O(N__43579),
            .I(N__43576));
    Odrv12 I__9748 (
            .O(N__43576),
            .I(ICE_SPI_MISO));
    InMux I__9747 (
            .O(N__43573),
            .I(N__43570));
    LocalMux I__9746 (
            .O(N__43570),
            .I(N__43566));
    InMux I__9745 (
            .O(N__43569),
            .I(N__43563));
    Span4Mux_v I__9744 (
            .O(N__43566),
            .I(N__43559));
    LocalMux I__9743 (
            .O(N__43563),
            .I(N__43556));
    InMux I__9742 (
            .O(N__43562),
            .I(N__43553));
    Odrv4 I__9741 (
            .O(N__43559),
            .I(\comm_spi.n22635 ));
    Odrv12 I__9740 (
            .O(N__43556),
            .I(\comm_spi.n22635 ));
    LocalMux I__9739 (
            .O(N__43553),
            .I(\comm_spi.n22635 ));
    InMux I__9738 (
            .O(N__43546),
            .I(N__43542));
    InMux I__9737 (
            .O(N__43545),
            .I(N__43539));
    LocalMux I__9736 (
            .O(N__43542),
            .I(\comm_spi.n14623 ));
    LocalMux I__9735 (
            .O(N__43539),
            .I(\comm_spi.n14623 ));
    CascadeMux I__9734 (
            .O(N__43534),
            .I(N__43529));
    CascadeMux I__9733 (
            .O(N__43533),
            .I(N__43526));
    CascadeMux I__9732 (
            .O(N__43532),
            .I(N__43521));
    InMux I__9731 (
            .O(N__43529),
            .I(N__43517));
    InMux I__9730 (
            .O(N__43526),
            .I(N__43514));
    CascadeMux I__9729 (
            .O(N__43525),
            .I(N__43511));
    InMux I__9728 (
            .O(N__43524),
            .I(N__43508));
    InMux I__9727 (
            .O(N__43521),
            .I(N__43505));
    InMux I__9726 (
            .O(N__43520),
            .I(N__43501));
    LocalMux I__9725 (
            .O(N__43517),
            .I(N__43496));
    LocalMux I__9724 (
            .O(N__43514),
            .I(N__43496));
    InMux I__9723 (
            .O(N__43511),
            .I(N__43493));
    LocalMux I__9722 (
            .O(N__43508),
            .I(N__43488));
    LocalMux I__9721 (
            .O(N__43505),
            .I(N__43488));
    CascadeMux I__9720 (
            .O(N__43504),
            .I(N__43484));
    LocalMux I__9719 (
            .O(N__43501),
            .I(N__43481));
    Span4Mux_v I__9718 (
            .O(N__43496),
            .I(N__43478));
    LocalMux I__9717 (
            .O(N__43493),
            .I(N__43475));
    Span4Mux_v I__9716 (
            .O(N__43488),
            .I(N__43471));
    InMux I__9715 (
            .O(N__43487),
            .I(N__43468));
    InMux I__9714 (
            .O(N__43484),
            .I(N__43465));
    Span4Mux_h I__9713 (
            .O(N__43481),
            .I(N__43462));
    Span4Mux_v I__9712 (
            .O(N__43478),
            .I(N__43456));
    Span4Mux_h I__9711 (
            .O(N__43475),
            .I(N__43456));
    InMux I__9710 (
            .O(N__43474),
            .I(N__43453));
    Sp12to4 I__9709 (
            .O(N__43471),
            .I(N__43450));
    LocalMux I__9708 (
            .O(N__43468),
            .I(N__43447));
    LocalMux I__9707 (
            .O(N__43465),
            .I(N__43444));
    Span4Mux_v I__9706 (
            .O(N__43462),
            .I(N__43441));
    InMux I__9705 (
            .O(N__43461),
            .I(N__43438));
    Span4Mux_h I__9704 (
            .O(N__43456),
            .I(N__43435));
    LocalMux I__9703 (
            .O(N__43453),
            .I(N__43428));
    Span12Mux_h I__9702 (
            .O(N__43450),
            .I(N__43428));
    Sp12to4 I__9701 (
            .O(N__43447),
            .I(N__43428));
    Odrv4 I__9700 (
            .O(N__43444),
            .I(comm_buf_0_0));
    Odrv4 I__9699 (
            .O(N__43441),
            .I(comm_buf_0_0));
    LocalMux I__9698 (
            .O(N__43438),
            .I(comm_buf_0_0));
    Odrv4 I__9697 (
            .O(N__43435),
            .I(comm_buf_0_0));
    Odrv12 I__9696 (
            .O(N__43428),
            .I(comm_buf_0_0));
    InMux I__9695 (
            .O(N__43417),
            .I(N__43414));
    LocalMux I__9694 (
            .O(N__43414),
            .I(N__43410));
    InMux I__9693 (
            .O(N__43413),
            .I(N__43406));
    Span4Mux_v I__9692 (
            .O(N__43410),
            .I(N__43403));
    InMux I__9691 (
            .O(N__43409),
            .I(N__43400));
    LocalMux I__9690 (
            .O(N__43406),
            .I(N__43397));
    Odrv4 I__9689 (
            .O(N__43403),
            .I(buf_dds0_8));
    LocalMux I__9688 (
            .O(N__43400),
            .I(buf_dds0_8));
    Odrv12 I__9687 (
            .O(N__43397),
            .I(buf_dds0_8));
    InMux I__9686 (
            .O(N__43390),
            .I(N__43387));
    LocalMux I__9685 (
            .O(N__43387),
            .I(N__43384));
    Span4Mux_v I__9684 (
            .O(N__43384),
            .I(N__43379));
    InMux I__9683 (
            .O(N__43383),
            .I(N__43376));
    InMux I__9682 (
            .O(N__43382),
            .I(N__43371));
    Span4Mux_v I__9681 (
            .O(N__43379),
            .I(N__43366));
    LocalMux I__9680 (
            .O(N__43376),
            .I(N__43366));
    InMux I__9679 (
            .O(N__43375),
            .I(N__43363));
    InMux I__9678 (
            .O(N__43374),
            .I(N__43360));
    LocalMux I__9677 (
            .O(N__43371),
            .I(N__43357));
    Span4Mux_v I__9676 (
            .O(N__43366),
            .I(N__43354));
    LocalMux I__9675 (
            .O(N__43363),
            .I(N__43351));
    LocalMux I__9674 (
            .O(N__43360),
            .I(N__43348));
    Span4Mux_h I__9673 (
            .O(N__43357),
            .I(N__43344));
    Span4Mux_h I__9672 (
            .O(N__43354),
            .I(N__43339));
    Span4Mux_v I__9671 (
            .O(N__43351),
            .I(N__43339));
    Span4Mux_v I__9670 (
            .O(N__43348),
            .I(N__43336));
    InMux I__9669 (
            .O(N__43347),
            .I(N__43333));
    Span4Mux_v I__9668 (
            .O(N__43344),
            .I(N__43328));
    Span4Mux_v I__9667 (
            .O(N__43339),
            .I(N__43328));
    Odrv4 I__9666 (
            .O(N__43336),
            .I(comm_buf_1_1));
    LocalMux I__9665 (
            .O(N__43333),
            .I(comm_buf_1_1));
    Odrv4 I__9664 (
            .O(N__43328),
            .I(comm_buf_1_1));
    InMux I__9663 (
            .O(N__43321),
            .I(N__43316));
    InMux I__9662 (
            .O(N__43320),
            .I(N__43313));
    InMux I__9661 (
            .O(N__43319),
            .I(N__43310));
    LocalMux I__9660 (
            .O(N__43316),
            .I(N__43305));
    LocalMux I__9659 (
            .O(N__43313),
            .I(N__43305));
    LocalMux I__9658 (
            .O(N__43310),
            .I(data_index_1));
    Odrv4 I__9657 (
            .O(N__43305),
            .I(data_index_1));
    InMux I__9656 (
            .O(N__43300),
            .I(N__43296));
    InMux I__9655 (
            .O(N__43299),
            .I(N__43292));
    LocalMux I__9654 (
            .O(N__43296),
            .I(N__43288));
    InMux I__9653 (
            .O(N__43295),
            .I(N__43285));
    LocalMux I__9652 (
            .O(N__43292),
            .I(N__43281));
    InMux I__9651 (
            .O(N__43291),
            .I(N__43278));
    Span4Mux_h I__9650 (
            .O(N__43288),
            .I(N__43268));
    LocalMux I__9649 (
            .O(N__43285),
            .I(N__43268));
    InMux I__9648 (
            .O(N__43284),
            .I(N__43265));
    Span4Mux_v I__9647 (
            .O(N__43281),
            .I(N__43260));
    LocalMux I__9646 (
            .O(N__43278),
            .I(N__43260));
    InMux I__9645 (
            .O(N__43277),
            .I(N__43257));
    InMux I__9644 (
            .O(N__43276),
            .I(N__43254));
    InMux I__9643 (
            .O(N__43275),
            .I(N__43249));
    InMux I__9642 (
            .O(N__43274),
            .I(N__43249));
    InMux I__9641 (
            .O(N__43273),
            .I(N__43246));
    Span4Mux_h I__9640 (
            .O(N__43268),
            .I(N__43243));
    LocalMux I__9639 (
            .O(N__43265),
            .I(n8780));
    Odrv4 I__9638 (
            .O(N__43260),
            .I(n8780));
    LocalMux I__9637 (
            .O(N__43257),
            .I(n8780));
    LocalMux I__9636 (
            .O(N__43254),
            .I(n8780));
    LocalMux I__9635 (
            .O(N__43249),
            .I(n8780));
    LocalMux I__9634 (
            .O(N__43246),
            .I(n8780));
    Odrv4 I__9633 (
            .O(N__43243),
            .I(n8780));
    InMux I__9632 (
            .O(N__43228),
            .I(N__43225));
    LocalMux I__9631 (
            .O(N__43225),
            .I(n8_adj_1547));
    CascadeMux I__9630 (
            .O(N__43222),
            .I(n8_adj_1547_cascade_));
    InMux I__9629 (
            .O(N__43219),
            .I(N__43213));
    InMux I__9628 (
            .O(N__43218),
            .I(N__43213));
    LocalMux I__9627 (
            .O(N__43213),
            .I(N__43210));
    Odrv12 I__9626 (
            .O(N__43210),
            .I(n7_adj_1546));
    CascadeMux I__9625 (
            .O(N__43207),
            .I(N__43204));
    CascadeBuf I__9624 (
            .O(N__43204),
            .I(N__43201));
    CascadeMux I__9623 (
            .O(N__43201),
            .I(N__43198));
    CascadeBuf I__9622 (
            .O(N__43198),
            .I(N__43195));
    CascadeMux I__9621 (
            .O(N__43195),
            .I(N__43192));
    CascadeBuf I__9620 (
            .O(N__43192),
            .I(N__43189));
    CascadeMux I__9619 (
            .O(N__43189),
            .I(N__43186));
    CascadeBuf I__9618 (
            .O(N__43186),
            .I(N__43183));
    CascadeMux I__9617 (
            .O(N__43183),
            .I(N__43180));
    CascadeBuf I__9616 (
            .O(N__43180),
            .I(N__43177));
    CascadeMux I__9615 (
            .O(N__43177),
            .I(N__43174));
    CascadeBuf I__9614 (
            .O(N__43174),
            .I(N__43171));
    CascadeMux I__9613 (
            .O(N__43171),
            .I(N__43168));
    CascadeBuf I__9612 (
            .O(N__43168),
            .I(N__43165));
    CascadeMux I__9611 (
            .O(N__43165),
            .I(N__43162));
    CascadeBuf I__9610 (
            .O(N__43162),
            .I(N__43159));
    CascadeMux I__9609 (
            .O(N__43159),
            .I(N__43155));
    CascadeMux I__9608 (
            .O(N__43158),
            .I(N__43152));
    CascadeBuf I__9607 (
            .O(N__43155),
            .I(N__43149));
    CascadeBuf I__9606 (
            .O(N__43152),
            .I(N__43146));
    CascadeMux I__9605 (
            .O(N__43149),
            .I(N__43143));
    CascadeMux I__9604 (
            .O(N__43146),
            .I(N__43140));
    InMux I__9603 (
            .O(N__43143),
            .I(N__43137));
    InMux I__9602 (
            .O(N__43140),
            .I(N__43134));
    LocalMux I__9601 (
            .O(N__43137),
            .I(N__43131));
    LocalMux I__9600 (
            .O(N__43134),
            .I(N__43128));
    Span4Mux_v I__9599 (
            .O(N__43131),
            .I(N__43125));
    Span4Mux_v I__9598 (
            .O(N__43128),
            .I(N__43122));
    Span4Mux_h I__9597 (
            .O(N__43125),
            .I(N__43119));
    Span4Mux_h I__9596 (
            .O(N__43122),
            .I(N__43116));
    Span4Mux_h I__9595 (
            .O(N__43119),
            .I(N__43113));
    Odrv4 I__9594 (
            .O(N__43116),
            .I(data_index_9_N_212_1));
    Odrv4 I__9593 (
            .O(N__43113),
            .I(data_index_9_N_212_1));
    CascadeMux I__9592 (
            .O(N__43108),
            .I(N__43105));
    InMux I__9591 (
            .O(N__43105),
            .I(N__43101));
    CascadeMux I__9590 (
            .O(N__43104),
            .I(N__43098));
    LocalMux I__9589 (
            .O(N__43101),
            .I(N__43094));
    InMux I__9588 (
            .O(N__43098),
            .I(N__43091));
    CascadeMux I__9587 (
            .O(N__43097),
            .I(N__43088));
    Span4Mux_v I__9586 (
            .O(N__43094),
            .I(N__43085));
    LocalMux I__9585 (
            .O(N__43091),
            .I(N__43082));
    InMux I__9584 (
            .O(N__43088),
            .I(N__43079));
    Span4Mux_h I__9583 (
            .O(N__43085),
            .I(N__43076));
    Span12Mux_h I__9582 (
            .O(N__43082),
            .I(N__43073));
    LocalMux I__9581 (
            .O(N__43079),
            .I(buf_dds0_11));
    Odrv4 I__9580 (
            .O(N__43076),
            .I(buf_dds0_11));
    Odrv12 I__9579 (
            .O(N__43073),
            .I(buf_dds0_11));
    InMux I__9578 (
            .O(N__43066),
            .I(N__43062));
    InMux I__9577 (
            .O(N__43065),
            .I(N__43059));
    LocalMux I__9576 (
            .O(N__43062),
            .I(N__43056));
    LocalMux I__9575 (
            .O(N__43059),
            .I(N__43050));
    Span4Mux_h I__9574 (
            .O(N__43056),
            .I(N__43050));
    InMux I__9573 (
            .O(N__43055),
            .I(N__43047));
    Span4Mux_h I__9572 (
            .O(N__43050),
            .I(N__43044));
    LocalMux I__9571 (
            .O(N__43047),
            .I(buf_dds0_5));
    Odrv4 I__9570 (
            .O(N__43044),
            .I(buf_dds0_5));
    InMux I__9569 (
            .O(N__43039),
            .I(N__43035));
    InMux I__9568 (
            .O(N__43038),
            .I(N__43032));
    LocalMux I__9567 (
            .O(N__43035),
            .I(N__43029));
    LocalMux I__9566 (
            .O(N__43032),
            .I(n8_adj_1532));
    Odrv4 I__9565 (
            .O(N__43029),
            .I(n8_adj_1532));
    InMux I__9564 (
            .O(N__43024),
            .I(N__43020));
    InMux I__9563 (
            .O(N__43023),
            .I(N__43017));
    LocalMux I__9562 (
            .O(N__43020),
            .I(N__43014));
    LocalMux I__9561 (
            .O(N__43017),
            .I(n7_adj_1531));
    Odrv12 I__9560 (
            .O(N__43014),
            .I(n7_adj_1531));
    CascadeMux I__9559 (
            .O(N__43009),
            .I(N__43006));
    CascadeBuf I__9558 (
            .O(N__43006),
            .I(N__43003));
    CascadeMux I__9557 (
            .O(N__43003),
            .I(N__43000));
    CascadeBuf I__9556 (
            .O(N__43000),
            .I(N__42997));
    CascadeMux I__9555 (
            .O(N__42997),
            .I(N__42994));
    CascadeBuf I__9554 (
            .O(N__42994),
            .I(N__42991));
    CascadeMux I__9553 (
            .O(N__42991),
            .I(N__42988));
    CascadeBuf I__9552 (
            .O(N__42988),
            .I(N__42985));
    CascadeMux I__9551 (
            .O(N__42985),
            .I(N__42982));
    CascadeBuf I__9550 (
            .O(N__42982),
            .I(N__42979));
    CascadeMux I__9549 (
            .O(N__42979),
            .I(N__42976));
    CascadeBuf I__9548 (
            .O(N__42976),
            .I(N__42973));
    CascadeMux I__9547 (
            .O(N__42973),
            .I(N__42970));
    CascadeBuf I__9546 (
            .O(N__42970),
            .I(N__42967));
    CascadeMux I__9545 (
            .O(N__42967),
            .I(N__42963));
    CascadeMux I__9544 (
            .O(N__42966),
            .I(N__42960));
    CascadeBuf I__9543 (
            .O(N__42963),
            .I(N__42957));
    CascadeBuf I__9542 (
            .O(N__42960),
            .I(N__42954));
    CascadeMux I__9541 (
            .O(N__42957),
            .I(N__42951));
    CascadeMux I__9540 (
            .O(N__42954),
            .I(N__42948));
    CascadeBuf I__9539 (
            .O(N__42951),
            .I(N__42945));
    InMux I__9538 (
            .O(N__42948),
            .I(N__42942));
    CascadeMux I__9537 (
            .O(N__42945),
            .I(N__42939));
    LocalMux I__9536 (
            .O(N__42942),
            .I(N__42936));
    InMux I__9535 (
            .O(N__42939),
            .I(N__42933));
    Span4Mux_v I__9534 (
            .O(N__42936),
            .I(N__42930));
    LocalMux I__9533 (
            .O(N__42933),
            .I(N__42927));
    Span4Mux_h I__9532 (
            .O(N__42930),
            .I(N__42924));
    Span12Mux_h I__9531 (
            .O(N__42927),
            .I(N__42921));
    Odrv4 I__9530 (
            .O(N__42924),
            .I(data_index_9_N_212_9));
    Odrv12 I__9529 (
            .O(N__42921),
            .I(data_index_9_N_212_9));
    CascadeMux I__9528 (
            .O(N__42916),
            .I(N__42912));
    InMux I__9527 (
            .O(N__42915),
            .I(N__42909));
    InMux I__9526 (
            .O(N__42912),
            .I(N__42906));
    LocalMux I__9525 (
            .O(N__42909),
            .I(tmp_buf_15));
    LocalMux I__9524 (
            .O(N__42906),
            .I(tmp_buf_15));
    IoInMux I__9523 (
            .O(N__42901),
            .I(N__42898));
    LocalMux I__9522 (
            .O(N__42898),
            .I(N__42895));
    IoSpan4Mux I__9521 (
            .O(N__42895),
            .I(N__42892));
    Span4Mux_s3_v I__9520 (
            .O(N__42892),
            .I(N__42889));
    Span4Mux_h I__9519 (
            .O(N__42889),
            .I(N__42886));
    Span4Mux_v I__9518 (
            .O(N__42886),
            .I(N__42882));
    InMux I__9517 (
            .O(N__42885),
            .I(N__42879));
    Odrv4 I__9516 (
            .O(N__42882),
            .I(DDS_MOSI));
    LocalMux I__9515 (
            .O(N__42879),
            .I(DDS_MOSI));
    InMux I__9514 (
            .O(N__42874),
            .I(N__42870));
    InMux I__9513 (
            .O(N__42873),
            .I(N__42867));
    LocalMux I__9512 (
            .O(N__42870),
            .I(N__42864));
    LocalMux I__9511 (
            .O(N__42867),
            .I(n7_adj_1515));
    Odrv12 I__9510 (
            .O(N__42864),
            .I(n7_adj_1515));
    InMux I__9509 (
            .O(N__42859),
            .I(N__42856));
    LocalMux I__9508 (
            .O(N__42856),
            .I(N__42852));
    InMux I__9507 (
            .O(N__42855),
            .I(N__42849));
    Span4Mux_h I__9506 (
            .O(N__42852),
            .I(N__42846));
    LocalMux I__9505 (
            .O(N__42849),
            .I(n17314));
    Odrv4 I__9504 (
            .O(N__42846),
            .I(n17314));
    InMux I__9503 (
            .O(N__42841),
            .I(N__42836));
    InMux I__9502 (
            .O(N__42840),
            .I(N__42833));
    InMux I__9501 (
            .O(N__42839),
            .I(N__42830));
    LocalMux I__9500 (
            .O(N__42836),
            .I(data_index_0));
    LocalMux I__9499 (
            .O(N__42833),
            .I(data_index_0));
    LocalMux I__9498 (
            .O(N__42830),
            .I(data_index_0));
    CascadeMux I__9497 (
            .O(N__42823),
            .I(N__42819));
    CascadeMux I__9496 (
            .O(N__42822),
            .I(N__42816));
    InMux I__9495 (
            .O(N__42819),
            .I(N__42812));
    InMux I__9494 (
            .O(N__42816),
            .I(N__42809));
    InMux I__9493 (
            .O(N__42815),
            .I(N__42805));
    LocalMux I__9492 (
            .O(N__42812),
            .I(N__42801));
    LocalMux I__9491 (
            .O(N__42809),
            .I(N__42798));
    CascadeMux I__9490 (
            .O(N__42808),
            .I(N__42795));
    LocalMux I__9489 (
            .O(N__42805),
            .I(N__42792));
    InMux I__9488 (
            .O(N__42804),
            .I(N__42789));
    Span4Mux_v I__9487 (
            .O(N__42801),
            .I(N__42785));
    Span4Mux_h I__9486 (
            .O(N__42798),
            .I(N__42782));
    InMux I__9485 (
            .O(N__42795),
            .I(N__42779));
    Span4Mux_h I__9484 (
            .O(N__42792),
            .I(N__42774));
    LocalMux I__9483 (
            .O(N__42789),
            .I(N__42774));
    InMux I__9482 (
            .O(N__42788),
            .I(N__42771));
    Sp12to4 I__9481 (
            .O(N__42785),
            .I(N__42768));
    Span4Mux_v I__9480 (
            .O(N__42782),
            .I(N__42759));
    LocalMux I__9479 (
            .O(N__42779),
            .I(N__42759));
    Span4Mux_v I__9478 (
            .O(N__42774),
            .I(N__42759));
    LocalMux I__9477 (
            .O(N__42771),
            .I(N__42759));
    Odrv12 I__9476 (
            .O(N__42768),
            .I(comm_buf_1_2));
    Odrv4 I__9475 (
            .O(N__42759),
            .I(comm_buf_1_2));
    InMux I__9474 (
            .O(N__42754),
            .I(N__42750));
    InMux I__9473 (
            .O(N__42753),
            .I(N__42747));
    LocalMux I__9472 (
            .O(N__42750),
            .I(N__42743));
    LocalMux I__9471 (
            .O(N__42747),
            .I(N__42740));
    InMux I__9470 (
            .O(N__42746),
            .I(N__42737));
    Span4Mux_v I__9469 (
            .O(N__42743),
            .I(N__42732));
    Span4Mux_h I__9468 (
            .O(N__42740),
            .I(N__42732));
    LocalMux I__9467 (
            .O(N__42737),
            .I(buf_dds0_2));
    Odrv4 I__9466 (
            .O(N__42732),
            .I(buf_dds0_2));
    InMux I__9465 (
            .O(N__42727),
            .I(N__42720));
    InMux I__9464 (
            .O(N__42726),
            .I(N__42720));
    InMux I__9463 (
            .O(N__42725),
            .I(N__42717));
    LocalMux I__9462 (
            .O(N__42720),
            .I(data_index_9));
    LocalMux I__9461 (
            .O(N__42717),
            .I(data_index_9));
    InMux I__9460 (
            .O(N__42712),
            .I(N__42708));
    InMux I__9459 (
            .O(N__42711),
            .I(N__42705));
    LocalMux I__9458 (
            .O(N__42708),
            .I(N__42702));
    LocalMux I__9457 (
            .O(N__42705),
            .I(N__42698));
    Span4Mux_h I__9456 (
            .O(N__42702),
            .I(N__42695));
    InMux I__9455 (
            .O(N__42701),
            .I(N__42692));
    Span4Mux_h I__9454 (
            .O(N__42698),
            .I(N__42689));
    Odrv4 I__9453 (
            .O(N__42695),
            .I(buf_dds0_4));
    LocalMux I__9452 (
            .O(N__42692),
            .I(buf_dds0_4));
    Odrv4 I__9451 (
            .O(N__42689),
            .I(buf_dds0_4));
    CascadeMux I__9450 (
            .O(N__42682),
            .I(n8_adj_1538_cascade_));
    InMux I__9449 (
            .O(N__42679),
            .I(N__42674));
    InMux I__9448 (
            .O(N__42678),
            .I(N__42671));
    InMux I__9447 (
            .O(N__42677),
            .I(N__42668));
    LocalMux I__9446 (
            .O(N__42674),
            .I(N__42663));
    LocalMux I__9445 (
            .O(N__42671),
            .I(N__42663));
    LocalMux I__9444 (
            .O(N__42668),
            .I(data_index_6));
    Odrv4 I__9443 (
            .O(N__42663),
            .I(data_index_6));
    InMux I__9442 (
            .O(N__42658),
            .I(N__42655));
    LocalMux I__9441 (
            .O(N__42655),
            .I(N__42651));
    InMux I__9440 (
            .O(N__42654),
            .I(N__42648));
    Span4Mux_h I__9439 (
            .O(N__42651),
            .I(N__42645));
    LocalMux I__9438 (
            .O(N__42648),
            .I(N__42641));
    Sp12to4 I__9437 (
            .O(N__42645),
            .I(N__42638));
    InMux I__9436 (
            .O(N__42644),
            .I(N__42635));
    Span4Mux_h I__9435 (
            .O(N__42641),
            .I(N__42632));
    Odrv12 I__9434 (
            .O(N__42638),
            .I(buf_dds0_6));
    LocalMux I__9433 (
            .O(N__42635),
            .I(buf_dds0_6));
    Odrv4 I__9432 (
            .O(N__42632),
            .I(buf_dds0_6));
    CascadeMux I__9431 (
            .O(N__42625),
            .I(N__42620));
    InMux I__9430 (
            .O(N__42624),
            .I(N__42616));
    InMux I__9429 (
            .O(N__42623),
            .I(N__42612));
    InMux I__9428 (
            .O(N__42620),
            .I(N__42609));
    CascadeMux I__9427 (
            .O(N__42619),
            .I(N__42606));
    LocalMux I__9426 (
            .O(N__42616),
            .I(N__42603));
    CascadeMux I__9425 (
            .O(N__42615),
            .I(N__42600));
    LocalMux I__9424 (
            .O(N__42612),
            .I(N__42597));
    LocalMux I__9423 (
            .O(N__42609),
            .I(N__42593));
    InMux I__9422 (
            .O(N__42606),
            .I(N__42590));
    Span4Mux_h I__9421 (
            .O(N__42603),
            .I(N__42587));
    InMux I__9420 (
            .O(N__42600),
            .I(N__42584));
    Span4Mux_v I__9419 (
            .O(N__42597),
            .I(N__42581));
    InMux I__9418 (
            .O(N__42596),
            .I(N__42578));
    Span4Mux_v I__9417 (
            .O(N__42593),
            .I(N__42575));
    LocalMux I__9416 (
            .O(N__42590),
            .I(N__42570));
    Span4Mux_v I__9415 (
            .O(N__42587),
            .I(N__42570));
    LocalMux I__9414 (
            .O(N__42584),
            .I(N__42567));
    Span4Mux_v I__9413 (
            .O(N__42581),
            .I(N__42562));
    LocalMux I__9412 (
            .O(N__42578),
            .I(N__42562));
    Span4Mux_h I__9411 (
            .O(N__42575),
            .I(N__42559));
    Span4Mux_v I__9410 (
            .O(N__42570),
            .I(N__42556));
    Span4Mux_h I__9409 (
            .O(N__42567),
            .I(N__42551));
    Span4Mux_h I__9408 (
            .O(N__42562),
            .I(N__42551));
    Odrv4 I__9407 (
            .O(N__42559),
            .I(comm_buf_1_7));
    Odrv4 I__9406 (
            .O(N__42556),
            .I(comm_buf_1_7));
    Odrv4 I__9405 (
            .O(N__42551),
            .I(comm_buf_1_7));
    InMux I__9404 (
            .O(N__42544),
            .I(N__42540));
    InMux I__9403 (
            .O(N__42543),
            .I(N__42537));
    LocalMux I__9402 (
            .O(N__42540),
            .I(N__42534));
    LocalMux I__9401 (
            .O(N__42537),
            .I(N__42531));
    Span4Mux_v I__9400 (
            .O(N__42534),
            .I(N__42527));
    Span4Mux_v I__9399 (
            .O(N__42531),
            .I(N__42524));
    InMux I__9398 (
            .O(N__42530),
            .I(N__42521));
    Span4Mux_h I__9397 (
            .O(N__42527),
            .I(N__42518));
    Span4Mux_h I__9396 (
            .O(N__42524),
            .I(N__42515));
    LocalMux I__9395 (
            .O(N__42521),
            .I(buf_dds1_7));
    Odrv4 I__9394 (
            .O(N__42518),
            .I(buf_dds1_7));
    Odrv4 I__9393 (
            .O(N__42515),
            .I(buf_dds1_7));
    InMux I__9392 (
            .O(N__42508),
            .I(N__42503));
    InMux I__9391 (
            .O(N__42507),
            .I(N__42500));
    InMux I__9390 (
            .O(N__42506),
            .I(N__42497));
    LocalMux I__9389 (
            .O(N__42503),
            .I(data_index_4));
    LocalMux I__9388 (
            .O(N__42500),
            .I(data_index_4));
    LocalMux I__9387 (
            .O(N__42497),
            .I(data_index_4));
    InMux I__9386 (
            .O(N__42490),
            .I(N__42484));
    InMux I__9385 (
            .O(N__42489),
            .I(N__42484));
    LocalMux I__9384 (
            .O(N__42484),
            .I(n7_adj_1540));
    InMux I__9383 (
            .O(N__42481),
            .I(n19329));
    InMux I__9382 (
            .O(N__42478),
            .I(n19330));
    InMux I__9381 (
            .O(N__42475),
            .I(n19331));
    InMux I__9380 (
            .O(N__42472),
            .I(N__42468));
    InMux I__9379 (
            .O(N__42471),
            .I(N__42465));
    LocalMux I__9378 (
            .O(N__42468),
            .I(N__42460));
    LocalMux I__9377 (
            .O(N__42465),
            .I(N__42460));
    Span4Mux_h I__9376 (
            .O(N__42460),
            .I(N__42456));
    InMux I__9375 (
            .O(N__42459),
            .I(N__42453));
    Span4Mux_h I__9374 (
            .O(N__42456),
            .I(N__42450));
    LocalMux I__9373 (
            .O(N__42453),
            .I(N__42447));
    Span4Mux_h I__9372 (
            .O(N__42450),
            .I(N__42444));
    Odrv12 I__9371 (
            .O(N__42447),
            .I(data_index_7));
    Odrv4 I__9370 (
            .O(N__42444),
            .I(data_index_7));
    InMux I__9369 (
            .O(N__42439),
            .I(N__42436));
    LocalMux I__9368 (
            .O(N__42436),
            .I(N__42432));
    InMux I__9367 (
            .O(N__42435),
            .I(N__42429));
    Span4Mux_h I__9366 (
            .O(N__42432),
            .I(N__42426));
    LocalMux I__9365 (
            .O(N__42429),
            .I(N__42423));
    Span4Mux_h I__9364 (
            .O(N__42426),
            .I(N__42420));
    Span12Mux_s11_v I__9363 (
            .O(N__42423),
            .I(N__42417));
    Odrv4 I__9362 (
            .O(N__42420),
            .I(n7_adj_1535));
    Odrv12 I__9361 (
            .O(N__42417),
            .I(n7_adj_1535));
    InMux I__9360 (
            .O(N__42412),
            .I(n19332));
    InMux I__9359 (
            .O(N__42409),
            .I(N__42405));
    InMux I__9358 (
            .O(N__42408),
            .I(N__42402));
    LocalMux I__9357 (
            .O(N__42405),
            .I(N__42397));
    LocalMux I__9356 (
            .O(N__42402),
            .I(N__42397));
    Span4Mux_v I__9355 (
            .O(N__42397),
            .I(N__42393));
    InMux I__9354 (
            .O(N__42396),
            .I(N__42390));
    Span4Mux_h I__9353 (
            .O(N__42393),
            .I(N__42387));
    LocalMux I__9352 (
            .O(N__42390),
            .I(data_index_8));
    Odrv4 I__9351 (
            .O(N__42387),
            .I(data_index_8));
    InMux I__9350 (
            .O(N__42382),
            .I(N__42376));
    InMux I__9349 (
            .O(N__42381),
            .I(N__42376));
    LocalMux I__9348 (
            .O(N__42376),
            .I(N__42373));
    Span4Mux_v I__9347 (
            .O(N__42373),
            .I(N__42370));
    Span4Mux_h I__9346 (
            .O(N__42370),
            .I(N__42367));
    Span4Mux_h I__9345 (
            .O(N__42367),
            .I(N__42364));
    Odrv4 I__9344 (
            .O(N__42364),
            .I(n7_adj_1533));
    InMux I__9343 (
            .O(N__42361),
            .I(bfn_16_16_0_));
    CascadeMux I__9342 (
            .O(N__42358),
            .I(N__42354));
    CascadeMux I__9341 (
            .O(N__42357),
            .I(N__42350));
    InMux I__9340 (
            .O(N__42354),
            .I(N__42347));
    CascadeMux I__9339 (
            .O(N__42353),
            .I(N__42336));
    InMux I__9338 (
            .O(N__42350),
            .I(N__42333));
    LocalMux I__9337 (
            .O(N__42347),
            .I(N__42330));
    CascadeMux I__9336 (
            .O(N__42346),
            .I(N__42327));
    CascadeMux I__9335 (
            .O(N__42345),
            .I(N__42324));
    CascadeMux I__9334 (
            .O(N__42344),
            .I(N__42321));
    CascadeMux I__9333 (
            .O(N__42343),
            .I(N__42318));
    CascadeMux I__9332 (
            .O(N__42342),
            .I(N__42315));
    CascadeMux I__9331 (
            .O(N__42341),
            .I(N__42312));
    CascadeMux I__9330 (
            .O(N__42340),
            .I(N__42309));
    CascadeMux I__9329 (
            .O(N__42339),
            .I(N__42306));
    InMux I__9328 (
            .O(N__42336),
            .I(N__42303));
    LocalMux I__9327 (
            .O(N__42333),
            .I(N__42300));
    Span4Mux_v I__9326 (
            .O(N__42330),
            .I(N__42297));
    InMux I__9325 (
            .O(N__42327),
            .I(N__42288));
    InMux I__9324 (
            .O(N__42324),
            .I(N__42288));
    InMux I__9323 (
            .O(N__42321),
            .I(N__42288));
    InMux I__9322 (
            .O(N__42318),
            .I(N__42288));
    InMux I__9321 (
            .O(N__42315),
            .I(N__42279));
    InMux I__9320 (
            .O(N__42312),
            .I(N__42279));
    InMux I__9319 (
            .O(N__42309),
            .I(N__42279));
    InMux I__9318 (
            .O(N__42306),
            .I(N__42279));
    LocalMux I__9317 (
            .O(N__42303),
            .I(n10579));
    Odrv4 I__9316 (
            .O(N__42300),
            .I(n10579));
    Odrv4 I__9315 (
            .O(N__42297),
            .I(n10579));
    LocalMux I__9314 (
            .O(N__42288),
            .I(n10579));
    LocalMux I__9313 (
            .O(N__42279),
            .I(n10579));
    InMux I__9312 (
            .O(N__42268),
            .I(n19334));
    CascadeMux I__9311 (
            .O(N__42265),
            .I(n17338_cascade_));
    CascadeMux I__9310 (
            .O(N__42262),
            .I(N__42259));
    CascadeBuf I__9309 (
            .O(N__42259),
            .I(N__42256));
    CascadeMux I__9308 (
            .O(N__42256),
            .I(N__42253));
    CascadeBuf I__9307 (
            .O(N__42253),
            .I(N__42250));
    CascadeMux I__9306 (
            .O(N__42250),
            .I(N__42247));
    CascadeBuf I__9305 (
            .O(N__42247),
            .I(N__42244));
    CascadeMux I__9304 (
            .O(N__42244),
            .I(N__42241));
    CascadeBuf I__9303 (
            .O(N__42241),
            .I(N__42238));
    CascadeMux I__9302 (
            .O(N__42238),
            .I(N__42235));
    CascadeBuf I__9301 (
            .O(N__42235),
            .I(N__42232));
    CascadeMux I__9300 (
            .O(N__42232),
            .I(N__42229));
    CascadeBuf I__9299 (
            .O(N__42229),
            .I(N__42226));
    CascadeMux I__9298 (
            .O(N__42226),
            .I(N__42223));
    CascadeBuf I__9297 (
            .O(N__42223),
            .I(N__42220));
    CascadeMux I__9296 (
            .O(N__42220),
            .I(N__42217));
    CascadeBuf I__9295 (
            .O(N__42217),
            .I(N__42213));
    CascadeMux I__9294 (
            .O(N__42216),
            .I(N__42210));
    CascadeMux I__9293 (
            .O(N__42213),
            .I(N__42207));
    CascadeBuf I__9292 (
            .O(N__42210),
            .I(N__42204));
    CascadeBuf I__9291 (
            .O(N__42207),
            .I(N__42201));
    CascadeMux I__9290 (
            .O(N__42204),
            .I(N__42198));
    CascadeMux I__9289 (
            .O(N__42201),
            .I(N__42195));
    InMux I__9288 (
            .O(N__42198),
            .I(N__42192));
    InMux I__9287 (
            .O(N__42195),
            .I(N__42189));
    LocalMux I__9286 (
            .O(N__42192),
            .I(N__42186));
    LocalMux I__9285 (
            .O(N__42189),
            .I(N__42183));
    Span4Mux_v I__9284 (
            .O(N__42186),
            .I(N__42180));
    Span12Mux_s10_v I__9283 (
            .O(N__42183),
            .I(N__42177));
    Sp12to4 I__9282 (
            .O(N__42180),
            .I(N__42172));
    Span12Mux_h I__9281 (
            .O(N__42177),
            .I(N__42172));
    Odrv12 I__9280 (
            .O(N__42172),
            .I(data_index_9_N_212_5));
    InMux I__9279 (
            .O(N__42169),
            .I(N__42166));
    LocalMux I__9278 (
            .O(N__42166),
            .I(N__42163));
    Odrv4 I__9277 (
            .O(N__42163),
            .I(n22_adj_1492));
    CascadeMux I__9276 (
            .O(N__42160),
            .I(n21_adj_1494_cascade_));
    InMux I__9275 (
            .O(N__42157),
            .I(N__42154));
    LocalMux I__9274 (
            .O(N__42154),
            .I(n24_adj_1530));
    InMux I__9273 (
            .O(N__42151),
            .I(N__42148));
    LocalMux I__9272 (
            .O(N__42148),
            .I(n30_adj_1597));
    CascadeMux I__9271 (
            .O(N__42145),
            .I(N__42140));
    InMux I__9270 (
            .O(N__42144),
            .I(N__42136));
    InMux I__9269 (
            .O(N__42143),
            .I(N__42132));
    InMux I__9268 (
            .O(N__42140),
            .I(N__42127));
    InMux I__9267 (
            .O(N__42139),
            .I(N__42127));
    LocalMux I__9266 (
            .O(N__42136),
            .I(N__42123));
    InMux I__9265 (
            .O(N__42135),
            .I(N__42120));
    LocalMux I__9264 (
            .O(N__42132),
            .I(N__42116));
    LocalMux I__9263 (
            .O(N__42127),
            .I(N__42113));
    InMux I__9262 (
            .O(N__42126),
            .I(N__42110));
    Span4Mux_h I__9261 (
            .O(N__42123),
            .I(N__42105));
    LocalMux I__9260 (
            .O(N__42120),
            .I(N__42105));
    InMux I__9259 (
            .O(N__42119),
            .I(N__42102));
    Span4Mux_v I__9258 (
            .O(N__42116),
            .I(N__42095));
    Span4Mux_v I__9257 (
            .O(N__42113),
            .I(N__42095));
    LocalMux I__9256 (
            .O(N__42110),
            .I(N__42095));
    Span4Mux_h I__9255 (
            .O(N__42105),
            .I(N__42090));
    LocalMux I__9254 (
            .O(N__42102),
            .I(N__42090));
    Span4Mux_h I__9253 (
            .O(N__42095),
            .I(N__42087));
    Span4Mux_v I__9252 (
            .O(N__42090),
            .I(N__42084));
    Span4Mux_v I__9251 (
            .O(N__42087),
            .I(N__42081));
    Odrv4 I__9250 (
            .O(N__42084),
            .I(n14_adj_1549));
    Odrv4 I__9249 (
            .O(N__42081),
            .I(n14_adj_1549));
    CascadeMux I__9248 (
            .O(N__42076),
            .I(N__42071));
    CascadeMux I__9247 (
            .O(N__42075),
            .I(N__42068));
    CascadeMux I__9246 (
            .O(N__42074),
            .I(N__42065));
    InMux I__9245 (
            .O(N__42071),
            .I(N__42062));
    InMux I__9244 (
            .O(N__42068),
            .I(N__42057));
    InMux I__9243 (
            .O(N__42065),
            .I(N__42057));
    LocalMux I__9242 (
            .O(N__42062),
            .I(N__42054));
    LocalMux I__9241 (
            .O(N__42057),
            .I(N__42051));
    Span4Mux_v I__9240 (
            .O(N__42054),
            .I(N__42046));
    Span4Mux_h I__9239 (
            .O(N__42051),
            .I(N__42046));
    Span4Mux_v I__9238 (
            .O(N__42046),
            .I(N__42041));
    InMux I__9237 (
            .O(N__42045),
            .I(N__42038));
    InMux I__9236 (
            .O(N__42044),
            .I(N__42035));
    Sp12to4 I__9235 (
            .O(N__42041),
            .I(N__42030));
    LocalMux I__9234 (
            .O(N__42038),
            .I(N__42030));
    LocalMux I__9233 (
            .O(N__42035),
            .I(buf_cfgRTD_4));
    Odrv12 I__9232 (
            .O(N__42030),
            .I(buf_cfgRTD_4));
    CascadeMux I__9231 (
            .O(N__42025),
            .I(N__42021));
    InMux I__9230 (
            .O(N__42024),
            .I(N__42016));
    InMux I__9229 (
            .O(N__42021),
            .I(N__42009));
    InMux I__9228 (
            .O(N__42020),
            .I(N__42009));
    InMux I__9227 (
            .O(N__42019),
            .I(N__42009));
    LocalMux I__9226 (
            .O(N__42016),
            .I(N__42001));
    LocalMux I__9225 (
            .O(N__42009),
            .I(N__41998));
    InMux I__9224 (
            .O(N__42008),
            .I(N__41993));
    InMux I__9223 (
            .O(N__42007),
            .I(N__41993));
    InMux I__9222 (
            .O(N__42006),
            .I(N__41980));
    InMux I__9221 (
            .O(N__42005),
            .I(N__41980));
    InMux I__9220 (
            .O(N__42004),
            .I(N__41980));
    Span4Mux_v I__9219 (
            .O(N__42001),
            .I(N__41973));
    Span4Mux_h I__9218 (
            .O(N__41998),
            .I(N__41973));
    LocalMux I__9217 (
            .O(N__41993),
            .I(N__41973));
    InMux I__9216 (
            .O(N__41992),
            .I(N__41968));
    InMux I__9215 (
            .O(N__41991),
            .I(N__41968));
    InMux I__9214 (
            .O(N__41990),
            .I(N__41959));
    InMux I__9213 (
            .O(N__41989),
            .I(N__41959));
    InMux I__9212 (
            .O(N__41988),
            .I(N__41959));
    InMux I__9211 (
            .O(N__41987),
            .I(N__41959));
    LocalMux I__9210 (
            .O(N__41980),
            .I(n12415));
    Odrv4 I__9209 (
            .O(N__41973),
            .I(n12415));
    LocalMux I__9208 (
            .O(N__41968),
            .I(n12415));
    LocalMux I__9207 (
            .O(N__41959),
            .I(n12415));
    InMux I__9206 (
            .O(N__41950),
            .I(N__41947));
    LocalMux I__9205 (
            .O(N__41947),
            .I(N__41944));
    Span4Mux_v I__9204 (
            .O(N__41944),
            .I(N__41940));
    InMux I__9203 (
            .O(N__41943),
            .I(N__41937));
    Span4Mux_h I__9202 (
            .O(N__41940),
            .I(N__41932));
    LocalMux I__9201 (
            .O(N__41937),
            .I(N__41932));
    Span4Mux_h I__9200 (
            .O(N__41932),
            .I(N__41929));
    Odrv4 I__9199 (
            .O(N__41929),
            .I(n14_adj_1551));
    CascadeMux I__9198 (
            .O(N__41926),
            .I(N__41923));
    InMux I__9197 (
            .O(N__41923),
            .I(N__41920));
    LocalMux I__9196 (
            .O(N__41920),
            .I(N__41917));
    Span4Mux_v I__9195 (
            .O(N__41917),
            .I(N__41914));
    Span4Mux_h I__9194 (
            .O(N__41914),
            .I(N__41909));
    InMux I__9193 (
            .O(N__41913),
            .I(N__41904));
    InMux I__9192 (
            .O(N__41912),
            .I(N__41904));
    Odrv4 I__9191 (
            .O(N__41909),
            .I(req_data_cnt_10));
    LocalMux I__9190 (
            .O(N__41904),
            .I(req_data_cnt_10));
    InMux I__9189 (
            .O(N__41899),
            .I(N__41896));
    LocalMux I__9188 (
            .O(N__41896),
            .I(N__41892));
    InMux I__9187 (
            .O(N__41895),
            .I(N__41888));
    Span12Mux_h I__9186 (
            .O(N__41892),
            .I(N__41885));
    InMux I__9185 (
            .O(N__41891),
            .I(N__41882));
    LocalMux I__9184 (
            .O(N__41888),
            .I(req_data_cnt_8));
    Odrv12 I__9183 (
            .O(N__41885),
            .I(req_data_cnt_8));
    LocalMux I__9182 (
            .O(N__41882),
            .I(req_data_cnt_8));
    InMux I__9181 (
            .O(N__41875),
            .I(N__41872));
    LocalMux I__9180 (
            .O(N__41872),
            .I(n19_adj_1499));
    InMux I__9179 (
            .O(N__41869),
            .I(bfn_16_15_0_));
    InMux I__9178 (
            .O(N__41866),
            .I(n19326));
    InMux I__9177 (
            .O(N__41863),
            .I(N__41858));
    InMux I__9176 (
            .O(N__41862),
            .I(N__41855));
    InMux I__9175 (
            .O(N__41861),
            .I(N__41852));
    LocalMux I__9174 (
            .O(N__41858),
            .I(N__41847));
    LocalMux I__9173 (
            .O(N__41855),
            .I(N__41847));
    LocalMux I__9172 (
            .O(N__41852),
            .I(data_index_2));
    Odrv12 I__9171 (
            .O(N__41847),
            .I(data_index_2));
    InMux I__9170 (
            .O(N__41842),
            .I(N__41836));
    InMux I__9169 (
            .O(N__41841),
            .I(N__41836));
    LocalMux I__9168 (
            .O(N__41836),
            .I(N__41833));
    Odrv4 I__9167 (
            .O(N__41833),
            .I(n7_adj_1544));
    InMux I__9166 (
            .O(N__41830),
            .I(n19327));
    InMux I__9165 (
            .O(N__41827),
            .I(N__41822));
    InMux I__9164 (
            .O(N__41826),
            .I(N__41819));
    InMux I__9163 (
            .O(N__41825),
            .I(N__41816));
    LocalMux I__9162 (
            .O(N__41822),
            .I(N__41813));
    LocalMux I__9161 (
            .O(N__41819),
            .I(N__41808));
    LocalMux I__9160 (
            .O(N__41816),
            .I(N__41808));
    Span4Mux_v I__9159 (
            .O(N__41813),
            .I(N__41805));
    Span4Mux_h I__9158 (
            .O(N__41808),
            .I(N__41802));
    Odrv4 I__9157 (
            .O(N__41805),
            .I(data_index_3));
    Odrv4 I__9156 (
            .O(N__41802),
            .I(data_index_3));
    InMux I__9155 (
            .O(N__41797),
            .I(N__41791));
    InMux I__9154 (
            .O(N__41796),
            .I(N__41791));
    LocalMux I__9153 (
            .O(N__41791),
            .I(N__41788));
    Odrv12 I__9152 (
            .O(N__41788),
            .I(n7_adj_1542));
    InMux I__9151 (
            .O(N__41785),
            .I(n19328));
    InMux I__9150 (
            .O(N__41782),
            .I(N__41778));
    InMux I__9149 (
            .O(N__41781),
            .I(N__41775));
    LocalMux I__9148 (
            .O(N__41778),
            .I(N__41772));
    LocalMux I__9147 (
            .O(N__41775),
            .I(N__41769));
    Span4Mux_v I__9146 (
            .O(N__41772),
            .I(N__41766));
    Span4Mux_v I__9145 (
            .O(N__41769),
            .I(N__41763));
    Span4Mux_h I__9144 (
            .O(N__41766),
            .I(N__41760));
    Span4Mux_v I__9143 (
            .O(N__41763),
            .I(N__41757));
    Odrv4 I__9142 (
            .O(N__41760),
            .I(n14_adj_1524));
    Odrv4 I__9141 (
            .O(N__41757),
            .I(n14_adj_1524));
    InMux I__9140 (
            .O(N__41752),
            .I(N__41748));
    CascadeMux I__9139 (
            .O(N__41751),
            .I(N__41745));
    LocalMux I__9138 (
            .O(N__41748),
            .I(N__41741));
    InMux I__9137 (
            .O(N__41745),
            .I(N__41738));
    InMux I__9136 (
            .O(N__41744),
            .I(N__41735));
    Span4Mux_v I__9135 (
            .O(N__41741),
            .I(N__41732));
    LocalMux I__9134 (
            .O(N__41738),
            .I(N__41729));
    LocalMux I__9133 (
            .O(N__41735),
            .I(req_data_cnt_0));
    Odrv4 I__9132 (
            .O(N__41732),
            .I(req_data_cnt_0));
    Odrv4 I__9131 (
            .O(N__41729),
            .I(req_data_cnt_0));
    InMux I__9130 (
            .O(N__41722),
            .I(N__41719));
    LocalMux I__9129 (
            .O(N__41719),
            .I(N__41715));
    InMux I__9128 (
            .O(N__41718),
            .I(N__41711));
    Span12Mux_v I__9127 (
            .O(N__41715),
            .I(N__41708));
    InMux I__9126 (
            .O(N__41714),
            .I(N__41705));
    LocalMux I__9125 (
            .O(N__41711),
            .I(req_data_cnt_6));
    Odrv12 I__9124 (
            .O(N__41708),
            .I(req_data_cnt_6));
    LocalMux I__9123 (
            .O(N__41705),
            .I(req_data_cnt_6));
    InMux I__9122 (
            .O(N__41698),
            .I(N__41695));
    LocalMux I__9121 (
            .O(N__41695),
            .I(n17_adj_1554));
    InMux I__9120 (
            .O(N__41692),
            .I(N__41688));
    CascadeMux I__9119 (
            .O(N__41691),
            .I(N__41685));
    LocalMux I__9118 (
            .O(N__41688),
            .I(N__41681));
    InMux I__9117 (
            .O(N__41685),
            .I(N__41678));
    InMux I__9116 (
            .O(N__41684),
            .I(N__41675));
    Span4Mux_h I__9115 (
            .O(N__41681),
            .I(N__41672));
    LocalMux I__9114 (
            .O(N__41678),
            .I(N__41669));
    LocalMux I__9113 (
            .O(N__41675),
            .I(N__41664));
    Span4Mux_v I__9112 (
            .O(N__41672),
            .I(N__41664));
    Span4Mux_v I__9111 (
            .O(N__41669),
            .I(N__41661));
    Odrv4 I__9110 (
            .O(N__41664),
            .I(req_data_cnt_15));
    Odrv4 I__9109 (
            .O(N__41661),
            .I(req_data_cnt_15));
    CascadeMux I__9108 (
            .O(N__41656),
            .I(N__41653));
    InMux I__9107 (
            .O(N__41653),
            .I(N__41650));
    LocalMux I__9106 (
            .O(N__41650),
            .I(N__41647));
    Span4Mux_h I__9105 (
            .O(N__41647),
            .I(N__41643));
    InMux I__9104 (
            .O(N__41646),
            .I(N__41639));
    Span4Mux_h I__9103 (
            .O(N__41643),
            .I(N__41636));
    InMux I__9102 (
            .O(N__41642),
            .I(N__41633));
    LocalMux I__9101 (
            .O(N__41639),
            .I(req_data_cnt_9));
    Odrv4 I__9100 (
            .O(N__41636),
            .I(req_data_cnt_9));
    LocalMux I__9099 (
            .O(N__41633),
            .I(req_data_cnt_9));
    InMux I__9098 (
            .O(N__41626),
            .I(N__41623));
    LocalMux I__9097 (
            .O(N__41623),
            .I(N__41619));
    InMux I__9096 (
            .O(N__41622),
            .I(N__41616));
    Span4Mux_v I__9095 (
            .O(N__41619),
            .I(N__41609));
    LocalMux I__9094 (
            .O(N__41616),
            .I(N__41609));
    InMux I__9093 (
            .O(N__41615),
            .I(N__41606));
    InMux I__9092 (
            .O(N__41614),
            .I(N__41603));
    Odrv4 I__9091 (
            .O(N__41609),
            .I(n20613));
    LocalMux I__9090 (
            .O(N__41606),
            .I(n20613));
    LocalMux I__9089 (
            .O(N__41603),
            .I(n20613));
    InMux I__9088 (
            .O(N__41596),
            .I(N__41593));
    LocalMux I__9087 (
            .O(N__41593),
            .I(N__41588));
    CascadeMux I__9086 (
            .O(N__41592),
            .I(N__41585));
    InMux I__9085 (
            .O(N__41591),
            .I(N__41582));
    Span4Mux_v I__9084 (
            .O(N__41588),
            .I(N__41579));
    InMux I__9083 (
            .O(N__41585),
            .I(N__41576));
    LocalMux I__9082 (
            .O(N__41582),
            .I(req_data_cnt_2));
    Odrv4 I__9081 (
            .O(N__41579),
            .I(req_data_cnt_2));
    LocalMux I__9080 (
            .O(N__41576),
            .I(req_data_cnt_2));
    InMux I__9079 (
            .O(N__41569),
            .I(N__41566));
    LocalMux I__9078 (
            .O(N__41566),
            .I(N__41562));
    InMux I__9077 (
            .O(N__41565),
            .I(N__41558));
    Span12Mux_v I__9076 (
            .O(N__41562),
            .I(N__41555));
    InMux I__9075 (
            .O(N__41561),
            .I(N__41552));
    LocalMux I__9074 (
            .O(N__41558),
            .I(req_data_cnt_7));
    Odrv12 I__9073 (
            .O(N__41555),
            .I(req_data_cnt_7));
    LocalMux I__9072 (
            .O(N__41552),
            .I(req_data_cnt_7));
    CascadeMux I__9071 (
            .O(N__41545),
            .I(N__41541));
    InMux I__9070 (
            .O(N__41544),
            .I(N__41536));
    InMux I__9069 (
            .O(N__41541),
            .I(N__41536));
    LocalMux I__9068 (
            .O(N__41536),
            .I(N__41532));
    CascadeMux I__9067 (
            .O(N__41535),
            .I(N__41529));
    Span4Mux_v I__9066 (
            .O(N__41532),
            .I(N__41523));
    InMux I__9065 (
            .O(N__41529),
            .I(N__41518));
    InMux I__9064 (
            .O(N__41528),
            .I(N__41518));
    InMux I__9063 (
            .O(N__41527),
            .I(N__41515));
    InMux I__9062 (
            .O(N__41526),
            .I(N__41512));
    Span4Mux_h I__9061 (
            .O(N__41523),
            .I(N__41507));
    LocalMux I__9060 (
            .O(N__41518),
            .I(N__41507));
    LocalMux I__9059 (
            .O(N__41515),
            .I(N__41503));
    LocalMux I__9058 (
            .O(N__41512),
            .I(N__41500));
    Span4Mux_v I__9057 (
            .O(N__41507),
            .I(N__41497));
    InMux I__9056 (
            .O(N__41506),
            .I(N__41494));
    Span4Mux_v I__9055 (
            .O(N__41503),
            .I(N__41491));
    Span4Mux_h I__9054 (
            .O(N__41500),
            .I(N__41488));
    Span4Mux_v I__9053 (
            .O(N__41497),
            .I(N__41485));
    LocalMux I__9052 (
            .O(N__41494),
            .I(N__41482));
    Span4Mux_h I__9051 (
            .O(N__41491),
            .I(N__41477));
    Span4Mux_v I__9050 (
            .O(N__41488),
            .I(N__41477));
    Odrv4 I__9049 (
            .O(N__41485),
            .I(n14_adj_1548));
    Odrv12 I__9048 (
            .O(N__41482),
            .I(n14_adj_1548));
    Odrv4 I__9047 (
            .O(N__41477),
            .I(n14_adj_1548));
    CascadeMux I__9046 (
            .O(N__41470),
            .I(N__41466));
    InMux I__9045 (
            .O(N__41469),
            .I(N__41463));
    InMux I__9044 (
            .O(N__41466),
            .I(N__41460));
    LocalMux I__9043 (
            .O(N__41463),
            .I(N__41457));
    LocalMux I__9042 (
            .O(N__41460),
            .I(N__41452));
    Span4Mux_h I__9041 (
            .O(N__41457),
            .I(N__41452));
    Odrv4 I__9040 (
            .O(N__41452),
            .I(data_idxvec_8));
    InMux I__9039 (
            .O(N__41449),
            .I(N__41446));
    LocalMux I__9038 (
            .O(N__41446),
            .I(N__41443));
    Odrv12 I__9037 (
            .O(N__41443),
            .I(n20779));
    CascadeMux I__9036 (
            .O(N__41440),
            .I(n12415_cascade_));
    CascadeMux I__9035 (
            .O(N__41437),
            .I(N__41433));
    CascadeMux I__9034 (
            .O(N__41436),
            .I(N__41430));
    InMux I__9033 (
            .O(N__41433),
            .I(N__41427));
    InMux I__9032 (
            .O(N__41430),
            .I(N__41422));
    LocalMux I__9031 (
            .O(N__41427),
            .I(N__41419));
    InMux I__9030 (
            .O(N__41426),
            .I(N__41416));
    InMux I__9029 (
            .O(N__41425),
            .I(N__41413));
    LocalMux I__9028 (
            .O(N__41422),
            .I(N__41410));
    Span4Mux_v I__9027 (
            .O(N__41419),
            .I(N__41405));
    LocalMux I__9026 (
            .O(N__41416),
            .I(N__41405));
    LocalMux I__9025 (
            .O(N__41413),
            .I(N__41402));
    Span4Mux_v I__9024 (
            .O(N__41410),
            .I(N__41399));
    Span4Mux_v I__9023 (
            .O(N__41405),
            .I(N__41396));
    Span4Mux_h I__9022 (
            .O(N__41402),
            .I(N__41393));
    Span4Mux_h I__9021 (
            .O(N__41399),
            .I(N__41390));
    Span4Mux_h I__9020 (
            .O(N__41396),
            .I(N__41387));
    Span4Mux_h I__9019 (
            .O(N__41393),
            .I(N__41383));
    Sp12to4 I__9018 (
            .O(N__41390),
            .I(N__41378));
    Sp12to4 I__9017 (
            .O(N__41387),
            .I(N__41378));
    InMux I__9016 (
            .O(N__41386),
            .I(N__41375));
    Span4Mux_h I__9015 (
            .O(N__41383),
            .I(N__41372));
    Odrv12 I__9014 (
            .O(N__41378),
            .I(buf_cfgRTD_5));
    LocalMux I__9013 (
            .O(N__41375),
            .I(buf_cfgRTD_5));
    Odrv4 I__9012 (
            .O(N__41372),
            .I(buf_cfgRTD_5));
    InMux I__9011 (
            .O(N__41365),
            .I(N__41360));
    CascadeMux I__9010 (
            .O(N__41364),
            .I(N__41357));
    CascadeMux I__9009 (
            .O(N__41363),
            .I(N__41351));
    LocalMux I__9008 (
            .O(N__41360),
            .I(N__41348));
    InMux I__9007 (
            .O(N__41357),
            .I(N__41342));
    InMux I__9006 (
            .O(N__41356),
            .I(N__41342));
    InMux I__9005 (
            .O(N__41355),
            .I(N__41339));
    InMux I__9004 (
            .O(N__41354),
            .I(N__41336));
    InMux I__9003 (
            .O(N__41351),
            .I(N__41333));
    Span4Mux_h I__9002 (
            .O(N__41348),
            .I(N__41330));
    InMux I__9001 (
            .O(N__41347),
            .I(N__41327));
    LocalMux I__9000 (
            .O(N__41342),
            .I(N__41324));
    LocalMux I__8999 (
            .O(N__41339),
            .I(N__41321));
    LocalMux I__8998 (
            .O(N__41336),
            .I(N__41318));
    LocalMux I__8997 (
            .O(N__41333),
            .I(N__41315));
    Span4Mux_v I__8996 (
            .O(N__41330),
            .I(N__41312));
    LocalMux I__8995 (
            .O(N__41327),
            .I(N__41309));
    Span4Mux_h I__8994 (
            .O(N__41324),
            .I(N__41306));
    Span12Mux_v I__8993 (
            .O(N__41321),
            .I(N__41303));
    Span4Mux_v I__8992 (
            .O(N__41318),
            .I(N__41300));
    Span4Mux_v I__8991 (
            .O(N__41315),
            .I(N__41293));
    Span4Mux_h I__8990 (
            .O(N__41312),
            .I(N__41293));
    Span4Mux_v I__8989 (
            .O(N__41309),
            .I(N__41293));
    Odrv4 I__8988 (
            .O(N__41306),
            .I(comm_buf_1_0));
    Odrv12 I__8987 (
            .O(N__41303),
            .I(comm_buf_1_0));
    Odrv4 I__8986 (
            .O(N__41300),
            .I(comm_buf_1_0));
    Odrv4 I__8985 (
            .O(N__41293),
            .I(comm_buf_1_0));
    InMux I__8984 (
            .O(N__41284),
            .I(N__41280));
    InMux I__8983 (
            .O(N__41283),
            .I(N__41277));
    LocalMux I__8982 (
            .O(N__41280),
            .I(N__41274));
    LocalMux I__8981 (
            .O(N__41277),
            .I(N__41269));
    Span4Mux_h I__8980 (
            .O(N__41274),
            .I(N__41269));
    Span4Mux_h I__8979 (
            .O(N__41269),
            .I(N__41266));
    Odrv4 I__8978 (
            .O(N__41266),
            .I(n14_adj_1528));
    InMux I__8977 (
            .O(N__41263),
            .I(N__41260));
    LocalMux I__8976 (
            .O(N__41260),
            .I(N__41256));
    InMux I__8975 (
            .O(N__41259),
            .I(N__41253));
    Span4Mux_h I__8974 (
            .O(N__41256),
            .I(N__41248));
    LocalMux I__8973 (
            .O(N__41253),
            .I(N__41248));
    Span4Mux_h I__8972 (
            .O(N__41248),
            .I(N__41245));
    Odrv4 I__8971 (
            .O(N__41245),
            .I(n14_adj_1525));
    InMux I__8970 (
            .O(N__41242),
            .I(N__41239));
    LocalMux I__8969 (
            .O(N__41239),
            .I(N__41236));
    Span12Mux_v I__8968 (
            .O(N__41236),
            .I(N__41233));
    Odrv12 I__8967 (
            .O(N__41233),
            .I(n20850));
    InMux I__8966 (
            .O(N__41230),
            .I(N__41227));
    LocalMux I__8965 (
            .O(N__41227),
            .I(N__41224));
    Span4Mux_h I__8964 (
            .O(N__41224),
            .I(N__41221));
    Span4Mux_h I__8963 (
            .O(N__41221),
            .I(N__41218));
    Odrv4 I__8962 (
            .O(N__41218),
            .I(n30_adj_1520));
    InMux I__8961 (
            .O(N__41215),
            .I(N__41212));
    LocalMux I__8960 (
            .O(N__41212),
            .I(N__41209));
    Span4Mux_v I__8959 (
            .O(N__41209),
            .I(N__41206));
    Odrv4 I__8958 (
            .O(N__41206),
            .I(n22_adj_1594));
    InMux I__8957 (
            .O(N__41203),
            .I(N__41200));
    LocalMux I__8956 (
            .O(N__41200),
            .I(n10_adj_1582));
    CascadeMux I__8955 (
            .O(N__41197),
            .I(N__41193));
    InMux I__8954 (
            .O(N__41196),
            .I(N__41190));
    InMux I__8953 (
            .O(N__41193),
            .I(N__41186));
    LocalMux I__8952 (
            .O(N__41190),
            .I(N__41183));
    InMux I__8951 (
            .O(N__41189),
            .I(N__41180));
    LocalMux I__8950 (
            .O(N__41186),
            .I(N__41177));
    Odrv12 I__8949 (
            .O(N__41183),
            .I(clk_cnt_1));
    LocalMux I__8948 (
            .O(N__41180),
            .I(clk_cnt_1));
    Odrv4 I__8947 (
            .O(N__41177),
            .I(clk_cnt_1));
    InMux I__8946 (
            .O(N__41170),
            .I(N__41166));
    InMux I__8945 (
            .O(N__41169),
            .I(N__41161));
    LocalMux I__8944 (
            .O(N__41166),
            .I(N__41158));
    InMux I__8943 (
            .O(N__41165),
            .I(N__41153));
    InMux I__8942 (
            .O(N__41164),
            .I(N__41153));
    LocalMux I__8941 (
            .O(N__41161),
            .I(N__41150));
    Odrv12 I__8940 (
            .O(N__41158),
            .I(clk_cnt_0));
    LocalMux I__8939 (
            .O(N__41153),
            .I(clk_cnt_0));
    Odrv4 I__8938 (
            .O(N__41150),
            .I(clk_cnt_0));
    ClkMux I__8937 (
            .O(N__41143),
            .I(N__41138));
    ClkMux I__8936 (
            .O(N__41142),
            .I(N__41135));
    ClkMux I__8935 (
            .O(N__41141),
            .I(N__41126));
    LocalMux I__8934 (
            .O(N__41138),
            .I(N__41123));
    LocalMux I__8933 (
            .O(N__41135),
            .I(N__41120));
    ClkMux I__8932 (
            .O(N__41134),
            .I(N__41117));
    ClkMux I__8931 (
            .O(N__41133),
            .I(N__41112));
    ClkMux I__8930 (
            .O(N__41132),
            .I(N__41109));
    ClkMux I__8929 (
            .O(N__41131),
            .I(N__41106));
    ClkMux I__8928 (
            .O(N__41130),
            .I(N__41103));
    ClkMux I__8927 (
            .O(N__41129),
            .I(N__41100));
    LocalMux I__8926 (
            .O(N__41126),
            .I(N__41094));
    Span4Mux_h I__8925 (
            .O(N__41123),
            .I(N__41087));
    Span4Mux_v I__8924 (
            .O(N__41120),
            .I(N__41087));
    LocalMux I__8923 (
            .O(N__41117),
            .I(N__41087));
    ClkMux I__8922 (
            .O(N__41116),
            .I(N__41084));
    ClkMux I__8921 (
            .O(N__41115),
            .I(N__41076));
    LocalMux I__8920 (
            .O(N__41112),
            .I(N__41073));
    LocalMux I__8919 (
            .O(N__41109),
            .I(N__41070));
    LocalMux I__8918 (
            .O(N__41106),
            .I(N__41067));
    LocalMux I__8917 (
            .O(N__41103),
            .I(N__41062));
    LocalMux I__8916 (
            .O(N__41100),
            .I(N__41062));
    ClkMux I__8915 (
            .O(N__41099),
            .I(N__41059));
    ClkMux I__8914 (
            .O(N__41098),
            .I(N__41056));
    ClkMux I__8913 (
            .O(N__41097),
            .I(N__41053));
    Span4Mux_h I__8912 (
            .O(N__41094),
            .I(N__41046));
    Span4Mux_h I__8911 (
            .O(N__41087),
            .I(N__41046));
    LocalMux I__8910 (
            .O(N__41084),
            .I(N__41046));
    ClkMux I__8909 (
            .O(N__41083),
            .I(N__41043));
    ClkMux I__8908 (
            .O(N__41082),
            .I(N__41040));
    ClkMux I__8907 (
            .O(N__41081),
            .I(N__41037));
    ClkMux I__8906 (
            .O(N__41080),
            .I(N__41034));
    ClkMux I__8905 (
            .O(N__41079),
            .I(N__41031));
    LocalMux I__8904 (
            .O(N__41076),
            .I(N__41026));
    Span4Mux_v I__8903 (
            .O(N__41073),
            .I(N__41026));
    Span4Mux_v I__8902 (
            .O(N__41070),
            .I(N__41017));
    Span4Mux_h I__8901 (
            .O(N__41067),
            .I(N__41017));
    Span4Mux_v I__8900 (
            .O(N__41062),
            .I(N__41017));
    LocalMux I__8899 (
            .O(N__41059),
            .I(N__41017));
    LocalMux I__8898 (
            .O(N__41056),
            .I(N__41012));
    LocalMux I__8897 (
            .O(N__41053),
            .I(N__41012));
    Span4Mux_v I__8896 (
            .O(N__41046),
            .I(N__41009));
    LocalMux I__8895 (
            .O(N__41043),
            .I(N__41006));
    LocalMux I__8894 (
            .O(N__41040),
            .I(N__41003));
    LocalMux I__8893 (
            .O(N__41037),
            .I(N__41000));
    LocalMux I__8892 (
            .O(N__41034),
            .I(N__40997));
    LocalMux I__8891 (
            .O(N__41031),
            .I(N__40994));
    Span4Mux_h I__8890 (
            .O(N__41026),
            .I(N__40987));
    Span4Mux_h I__8889 (
            .O(N__41017),
            .I(N__40987));
    Span4Mux_v I__8888 (
            .O(N__41012),
            .I(N__40987));
    Span4Mux_h I__8887 (
            .O(N__41009),
            .I(N__40984));
    Span4Mux_v I__8886 (
            .O(N__41006),
            .I(N__40979));
    Span4Mux_v I__8885 (
            .O(N__41003),
            .I(N__40979));
    Span4Mux_v I__8884 (
            .O(N__41000),
            .I(N__40970));
    Span4Mux_v I__8883 (
            .O(N__40997),
            .I(N__40970));
    Span4Mux_v I__8882 (
            .O(N__40994),
            .I(N__40970));
    Span4Mux_h I__8881 (
            .O(N__40987),
            .I(N__40970));
    Span4Mux_h I__8880 (
            .O(N__40984),
            .I(N__40967));
    Sp12to4 I__8879 (
            .O(N__40979),
            .I(N__40962));
    Sp12to4 I__8878 (
            .O(N__40970),
            .I(N__40962));
    Span4Mux_h I__8877 (
            .O(N__40967),
            .I(N__40958));
    Span12Mux_h I__8876 (
            .O(N__40962),
            .I(N__40955));
    InMux I__8875 (
            .O(N__40961),
            .I(N__40952));
    Odrv4 I__8874 (
            .O(N__40958),
            .I(clk_RTD));
    Odrv12 I__8873 (
            .O(N__40955),
            .I(clk_RTD));
    LocalMux I__8872 (
            .O(N__40952),
            .I(clk_RTD));
    IoInMux I__8871 (
            .O(N__40945),
            .I(N__40942));
    LocalMux I__8870 (
            .O(N__40942),
            .I(N__40939));
    IoSpan4Mux I__8869 (
            .O(N__40939),
            .I(N__40935));
    ClkMux I__8868 (
            .O(N__40938),
            .I(N__40932));
    Span4Mux_s1_v I__8867 (
            .O(N__40935),
            .I(N__40929));
    LocalMux I__8866 (
            .O(N__40932),
            .I(N__40925));
    Sp12to4 I__8865 (
            .O(N__40929),
            .I(N__40922));
    ClkMux I__8864 (
            .O(N__40928),
            .I(N__40919));
    Span4Mux_h I__8863 (
            .O(N__40925),
            .I(N__40916));
    Span12Mux_h I__8862 (
            .O(N__40922),
            .I(N__40913));
    LocalMux I__8861 (
            .O(N__40919),
            .I(N__40910));
    Span4Mux_v I__8860 (
            .O(N__40916),
            .I(N__40907));
    Span12Mux_v I__8859 (
            .O(N__40913),
            .I(N__40901));
    Span12Mux_h I__8858 (
            .O(N__40910),
            .I(N__40901));
    Span4Mux_h I__8857 (
            .O(N__40907),
            .I(N__40898));
    InMux I__8856 (
            .O(N__40906),
            .I(N__40895));
    Odrv12 I__8855 (
            .O(N__40901),
            .I(TEST_LED));
    Odrv4 I__8854 (
            .O(N__40898),
            .I(TEST_LED));
    LocalMux I__8853 (
            .O(N__40895),
            .I(TEST_LED));
    InMux I__8852 (
            .O(N__40888),
            .I(N__40885));
    LocalMux I__8851 (
            .O(N__40885),
            .I(N__40882));
    Span4Mux_h I__8850 (
            .O(N__40882),
            .I(N__40878));
    CascadeMux I__8849 (
            .O(N__40881),
            .I(N__40875));
    Span4Mux_v I__8848 (
            .O(N__40878),
            .I(N__40872));
    InMux I__8847 (
            .O(N__40875),
            .I(N__40869));
    Odrv4 I__8846 (
            .O(N__40872),
            .I(buf_adcdata_vdc_6));
    LocalMux I__8845 (
            .O(N__40869),
            .I(buf_adcdata_vdc_6));
    InMux I__8844 (
            .O(N__40864),
            .I(N__40861));
    LocalMux I__8843 (
            .O(N__40861),
            .I(N__40857));
    InMux I__8842 (
            .O(N__40860),
            .I(N__40854));
    Span4Mux_v I__8841 (
            .O(N__40857),
            .I(N__40850));
    LocalMux I__8840 (
            .O(N__40854),
            .I(N__40847));
    InMux I__8839 (
            .O(N__40853),
            .I(N__40844));
    Sp12to4 I__8838 (
            .O(N__40850),
            .I(N__40841));
    Span4Mux_v I__8837 (
            .O(N__40847),
            .I(N__40838));
    LocalMux I__8836 (
            .O(N__40844),
            .I(buf_adcdata_vac_6));
    Odrv12 I__8835 (
            .O(N__40841),
            .I(buf_adcdata_vac_6));
    Odrv4 I__8834 (
            .O(N__40838),
            .I(buf_adcdata_vac_6));
    InMux I__8833 (
            .O(N__40831),
            .I(N__40828));
    LocalMux I__8832 (
            .O(N__40828),
            .I(n19_adj_1593));
    CascadeMux I__8831 (
            .O(N__40825),
            .I(N__40822));
    InMux I__8830 (
            .O(N__40822),
            .I(N__40819));
    LocalMux I__8829 (
            .O(N__40819),
            .I(N__40816));
    Odrv12 I__8828 (
            .O(N__40816),
            .I(n21071));
    InMux I__8827 (
            .O(N__40813),
            .I(N__40810));
    LocalMux I__8826 (
            .O(N__40810),
            .I(N__40807));
    Odrv4 I__8825 (
            .O(N__40807),
            .I(n20_adj_1607));
    InMux I__8824 (
            .O(N__40804),
            .I(N__40801));
    LocalMux I__8823 (
            .O(N__40801),
            .I(N__40798));
    Odrv12 I__8822 (
            .O(N__40798),
            .I(comm_buf_5_4));
    InMux I__8821 (
            .O(N__40795),
            .I(N__40792));
    LocalMux I__8820 (
            .O(N__40792),
            .I(N__40789));
    Odrv12 I__8819 (
            .O(N__40789),
            .I(comm_buf_4_4));
    InMux I__8818 (
            .O(N__40786),
            .I(N__40781));
    InMux I__8817 (
            .O(N__40785),
            .I(N__40778));
    InMux I__8816 (
            .O(N__40784),
            .I(N__40775));
    LocalMux I__8815 (
            .O(N__40781),
            .I(N__40772));
    LocalMux I__8814 (
            .O(N__40778),
            .I(N__40769));
    LocalMux I__8813 (
            .O(N__40775),
            .I(N__40766));
    Span4Mux_v I__8812 (
            .O(N__40772),
            .I(N__40763));
    Span4Mux_v I__8811 (
            .O(N__40769),
            .I(N__40760));
    Sp12to4 I__8810 (
            .O(N__40766),
            .I(N__40757));
    Sp12to4 I__8809 (
            .O(N__40763),
            .I(N__40750));
    Sp12to4 I__8808 (
            .O(N__40760),
            .I(N__40750));
    Span12Mux_v I__8807 (
            .O(N__40757),
            .I(N__40750));
    Odrv12 I__8806 (
            .O(N__40750),
            .I(comm_buf_0_6));
    InMux I__8805 (
            .O(N__40747),
            .I(N__40744));
    LocalMux I__8804 (
            .O(N__40744),
            .I(n28));
    InMux I__8803 (
            .O(N__40741),
            .I(N__40738));
    LocalMux I__8802 (
            .O(N__40738),
            .I(n27));
    CascadeMux I__8801 (
            .O(N__40735),
            .I(n26_adj_1625_cascade_));
    InMux I__8800 (
            .O(N__40732),
            .I(N__40729));
    LocalMux I__8799 (
            .O(N__40729),
            .I(n25_adj_1616));
    CascadeMux I__8798 (
            .O(N__40726),
            .I(n19553_cascade_));
    SRMux I__8797 (
            .O(N__40723),
            .I(N__40720));
    LocalMux I__8796 (
            .O(N__40720),
            .I(N__40717));
    Span4Mux_v I__8795 (
            .O(N__40717),
            .I(N__40714));
    Odrv4 I__8794 (
            .O(N__40714),
            .I(n17393));
    CascadeMux I__8793 (
            .O(N__40711),
            .I(N__40708));
    InMux I__8792 (
            .O(N__40708),
            .I(N__40705));
    LocalMux I__8791 (
            .O(N__40705),
            .I(N__40702));
    Span4Mux_h I__8790 (
            .O(N__40702),
            .I(N__40699));
    Span4Mux_v I__8789 (
            .O(N__40699),
            .I(N__40696));
    Span4Mux_h I__8788 (
            .O(N__40696),
            .I(N__40693));
    Odrv4 I__8787 (
            .O(N__40693),
            .I(n30));
    CascadeMux I__8786 (
            .O(N__40690),
            .I(comm_state_3_N_412_3_cascade_));
    CascadeMux I__8785 (
            .O(N__40687),
            .I(n20700_cascade_));
    SRMux I__8784 (
            .O(N__40684),
            .I(N__40680));
    SRMux I__8783 (
            .O(N__40683),
            .I(N__40677));
    LocalMux I__8782 (
            .O(N__40680),
            .I(N__40674));
    LocalMux I__8781 (
            .O(N__40677),
            .I(N__40671));
    Span4Mux_v I__8780 (
            .O(N__40674),
            .I(N__40668));
    Span4Mux_h I__8779 (
            .O(N__40671),
            .I(N__40665));
    Odrv4 I__8778 (
            .O(N__40668),
            .I(flagcntwd));
    Odrv4 I__8777 (
            .O(N__40665),
            .I(flagcntwd));
    CEMux I__8776 (
            .O(N__40660),
            .I(N__40657));
    LocalMux I__8775 (
            .O(N__40657),
            .I(N__40654));
    Span4Mux_h I__8774 (
            .O(N__40654),
            .I(N__40651));
    Odrv4 I__8773 (
            .O(N__40651),
            .I(n11411));
    SRMux I__8772 (
            .O(N__40648),
            .I(N__40645));
    LocalMux I__8771 (
            .O(N__40645),
            .I(N__40642));
    Span4Mux_v I__8770 (
            .O(N__40642),
            .I(N__40638));
    SRMux I__8769 (
            .O(N__40641),
            .I(N__40635));
    Span4Mux_v I__8768 (
            .O(N__40638),
            .I(N__40632));
    LocalMux I__8767 (
            .O(N__40635),
            .I(N__40629));
    Span4Mux_h I__8766 (
            .O(N__40632),
            .I(N__40626));
    Odrv4 I__8765 (
            .O(N__40629),
            .I(n20081));
    Odrv4 I__8764 (
            .O(N__40626),
            .I(n20081));
    CascadeMux I__8763 (
            .O(N__40621),
            .I(N__40618));
    InMux I__8762 (
            .O(N__40618),
            .I(N__40615));
    LocalMux I__8761 (
            .O(N__40615),
            .I(N__40612));
    Span4Mux_h I__8760 (
            .O(N__40612),
            .I(N__40609));
    Span4Mux_h I__8759 (
            .O(N__40609),
            .I(N__40606));
    Odrv4 I__8758 (
            .O(N__40606),
            .I(n11333));
    CascadeMux I__8757 (
            .O(N__40603),
            .I(N__40600));
    CascadeBuf I__8756 (
            .O(N__40600),
            .I(N__40597));
    CascadeMux I__8755 (
            .O(N__40597),
            .I(N__40594));
    CascadeBuf I__8754 (
            .O(N__40594),
            .I(N__40591));
    CascadeMux I__8753 (
            .O(N__40591),
            .I(N__40588));
    CascadeBuf I__8752 (
            .O(N__40588),
            .I(N__40585));
    CascadeMux I__8751 (
            .O(N__40585),
            .I(N__40582));
    CascadeBuf I__8750 (
            .O(N__40582),
            .I(N__40579));
    CascadeMux I__8749 (
            .O(N__40579),
            .I(N__40576));
    CascadeBuf I__8748 (
            .O(N__40576),
            .I(N__40573));
    CascadeMux I__8747 (
            .O(N__40573),
            .I(N__40570));
    CascadeBuf I__8746 (
            .O(N__40570),
            .I(N__40567));
    CascadeMux I__8745 (
            .O(N__40567),
            .I(N__40564));
    CascadeBuf I__8744 (
            .O(N__40564),
            .I(N__40561));
    CascadeMux I__8743 (
            .O(N__40561),
            .I(N__40558));
    CascadeBuf I__8742 (
            .O(N__40558),
            .I(N__40555));
    CascadeMux I__8741 (
            .O(N__40555),
            .I(N__40552));
    CascadeBuf I__8740 (
            .O(N__40552),
            .I(N__40548));
    CascadeMux I__8739 (
            .O(N__40551),
            .I(N__40545));
    CascadeMux I__8738 (
            .O(N__40548),
            .I(N__40542));
    CascadeBuf I__8737 (
            .O(N__40545),
            .I(N__40539));
    InMux I__8736 (
            .O(N__40542),
            .I(N__40536));
    CascadeMux I__8735 (
            .O(N__40539),
            .I(N__40533));
    LocalMux I__8734 (
            .O(N__40536),
            .I(N__40530));
    InMux I__8733 (
            .O(N__40533),
            .I(N__40527));
    Span4Mux_h I__8732 (
            .O(N__40530),
            .I(N__40524));
    LocalMux I__8731 (
            .O(N__40527),
            .I(N__40520));
    Span4Mux_h I__8730 (
            .O(N__40524),
            .I(N__40517));
    InMux I__8729 (
            .O(N__40523),
            .I(N__40514));
    Span12Mux_h I__8728 (
            .O(N__40520),
            .I(N__40511));
    Span4Mux_h I__8727 (
            .O(N__40517),
            .I(N__40508));
    LocalMux I__8726 (
            .O(N__40514),
            .I(data_count_8));
    Odrv12 I__8725 (
            .O(N__40511),
            .I(data_count_8));
    Odrv4 I__8724 (
            .O(N__40508),
            .I(data_count_8));
    InMux I__8723 (
            .O(N__40501),
            .I(bfn_15_18_0_));
    InMux I__8722 (
            .O(N__40498),
            .I(n19295));
    CascadeMux I__8721 (
            .O(N__40495),
            .I(N__40492));
    CascadeBuf I__8720 (
            .O(N__40492),
            .I(N__40489));
    CascadeMux I__8719 (
            .O(N__40489),
            .I(N__40486));
    CascadeBuf I__8718 (
            .O(N__40486),
            .I(N__40483));
    CascadeMux I__8717 (
            .O(N__40483),
            .I(N__40480));
    CascadeBuf I__8716 (
            .O(N__40480),
            .I(N__40477));
    CascadeMux I__8715 (
            .O(N__40477),
            .I(N__40474));
    CascadeBuf I__8714 (
            .O(N__40474),
            .I(N__40471));
    CascadeMux I__8713 (
            .O(N__40471),
            .I(N__40468));
    CascadeBuf I__8712 (
            .O(N__40468),
            .I(N__40465));
    CascadeMux I__8711 (
            .O(N__40465),
            .I(N__40462));
    CascadeBuf I__8710 (
            .O(N__40462),
            .I(N__40459));
    CascadeMux I__8709 (
            .O(N__40459),
            .I(N__40456));
    CascadeBuf I__8708 (
            .O(N__40456),
            .I(N__40453));
    CascadeMux I__8707 (
            .O(N__40453),
            .I(N__40450));
    CascadeBuf I__8706 (
            .O(N__40450),
            .I(N__40447));
    CascadeMux I__8705 (
            .O(N__40447),
            .I(N__40443));
    CascadeMux I__8704 (
            .O(N__40446),
            .I(N__40440));
    CascadeBuf I__8703 (
            .O(N__40443),
            .I(N__40437));
    CascadeBuf I__8702 (
            .O(N__40440),
            .I(N__40434));
    CascadeMux I__8701 (
            .O(N__40437),
            .I(N__40431));
    CascadeMux I__8700 (
            .O(N__40434),
            .I(N__40428));
    InMux I__8699 (
            .O(N__40431),
            .I(N__40425));
    InMux I__8698 (
            .O(N__40428),
            .I(N__40422));
    LocalMux I__8697 (
            .O(N__40425),
            .I(N__40419));
    LocalMux I__8696 (
            .O(N__40422),
            .I(N__40416));
    Span4Mux_h I__8695 (
            .O(N__40419),
            .I(N__40413));
    Span4Mux_h I__8694 (
            .O(N__40416),
            .I(N__40409));
    Span4Mux_h I__8693 (
            .O(N__40413),
            .I(N__40406));
    InMux I__8692 (
            .O(N__40412),
            .I(N__40403));
    Span4Mux_v I__8691 (
            .O(N__40409),
            .I(N__40400));
    Span4Mux_h I__8690 (
            .O(N__40406),
            .I(N__40397));
    LocalMux I__8689 (
            .O(N__40403),
            .I(data_count_9));
    Odrv4 I__8688 (
            .O(N__40400),
            .I(data_count_9));
    Odrv4 I__8687 (
            .O(N__40397),
            .I(data_count_9));
    CascadeMux I__8686 (
            .O(N__40390),
            .I(N__40387));
    InMux I__8685 (
            .O(N__40387),
            .I(N__40384));
    LocalMux I__8684 (
            .O(N__40384),
            .I(N__40381));
    Span4Mux_h I__8683 (
            .O(N__40381),
            .I(N__40378));
    Odrv4 I__8682 (
            .O(N__40378),
            .I(\SIG_DDS.tmp_buf_14 ));
    InMux I__8681 (
            .O(N__40375),
            .I(N__40370));
    InMux I__8680 (
            .O(N__40374),
            .I(N__40367));
    CascadeMux I__8679 (
            .O(N__40373),
            .I(N__40364));
    LocalMux I__8678 (
            .O(N__40370),
            .I(N__40361));
    LocalMux I__8677 (
            .O(N__40367),
            .I(N__40358));
    InMux I__8676 (
            .O(N__40364),
            .I(N__40355));
    Span4Mux_h I__8675 (
            .O(N__40361),
            .I(N__40352));
    Span4Mux_h I__8674 (
            .O(N__40358),
            .I(N__40349));
    LocalMux I__8673 (
            .O(N__40355),
            .I(buf_dds0_0));
    Odrv4 I__8672 (
            .O(N__40352),
            .I(buf_dds0_0));
    Odrv4 I__8671 (
            .O(N__40349),
            .I(buf_dds0_0));
    CascadeMux I__8670 (
            .O(N__40342),
            .I(N__40339));
    InMux I__8669 (
            .O(N__40339),
            .I(N__40336));
    LocalMux I__8668 (
            .O(N__40336),
            .I(N__40333));
    Odrv4 I__8667 (
            .O(N__40333),
            .I(\SIG_DDS.tmp_buf_0 ));
    CEMux I__8666 (
            .O(N__40330),
            .I(N__40326));
    CEMux I__8665 (
            .O(N__40329),
            .I(N__40323));
    LocalMux I__8664 (
            .O(N__40326),
            .I(N__40320));
    LocalMux I__8663 (
            .O(N__40323),
            .I(N__40317));
    Span4Mux_h I__8662 (
            .O(N__40320),
            .I(N__40311));
    Span4Mux_h I__8661 (
            .O(N__40317),
            .I(N__40308));
    CEMux I__8660 (
            .O(N__40316),
            .I(N__40305));
    CEMux I__8659 (
            .O(N__40315),
            .I(N__40302));
    CEMux I__8658 (
            .O(N__40314),
            .I(N__40299));
    Odrv4 I__8657 (
            .O(N__40311),
            .I(\SIG_DDS.n12700 ));
    Odrv4 I__8656 (
            .O(N__40308),
            .I(\SIG_DDS.n12700 ));
    LocalMux I__8655 (
            .O(N__40305),
            .I(\SIG_DDS.n12700 ));
    LocalMux I__8654 (
            .O(N__40302),
            .I(\SIG_DDS.n12700 ));
    LocalMux I__8653 (
            .O(N__40299),
            .I(\SIG_DDS.n12700 ));
    InMux I__8652 (
            .O(N__40288),
            .I(N__40285));
    LocalMux I__8651 (
            .O(N__40285),
            .I(N__40282));
    Span4Mux_v I__8650 (
            .O(N__40282),
            .I(N__40279));
    Span4Mux_v I__8649 (
            .O(N__40279),
            .I(N__40276));
    Span4Mux_h I__8648 (
            .O(N__40276),
            .I(N__40271));
    InMux I__8647 (
            .O(N__40275),
            .I(N__40266));
    InMux I__8646 (
            .O(N__40274),
            .I(N__40266));
    Odrv4 I__8645 (
            .O(N__40271),
            .I(comm_tx_buf_6));
    LocalMux I__8644 (
            .O(N__40266),
            .I(comm_tx_buf_6));
    SRMux I__8643 (
            .O(N__40261),
            .I(N__40257));
    SRMux I__8642 (
            .O(N__40260),
            .I(N__40253));
    LocalMux I__8641 (
            .O(N__40257),
            .I(N__40250));
    SRMux I__8640 (
            .O(N__40256),
            .I(N__40247));
    LocalMux I__8639 (
            .O(N__40253),
            .I(N__40242));
    Span4Mux_h I__8638 (
            .O(N__40250),
            .I(N__40242));
    LocalMux I__8637 (
            .O(N__40247),
            .I(N__40239));
    Odrv4 I__8636 (
            .O(N__40242),
            .I(\comm_spi.data_tx_7__N_758 ));
    Odrv4 I__8635 (
            .O(N__40239),
            .I(\comm_spi.data_tx_7__N_758 ));
    InMux I__8634 (
            .O(N__40234),
            .I(N__40231));
    LocalMux I__8633 (
            .O(N__40231),
            .I(N__40226));
    InMux I__8632 (
            .O(N__40230),
            .I(N__40223));
    InMux I__8631 (
            .O(N__40229),
            .I(N__40220));
    Odrv4 I__8630 (
            .O(N__40226),
            .I(\comm_spi.n22623 ));
    LocalMux I__8629 (
            .O(N__40223),
            .I(\comm_spi.n22623 ));
    LocalMux I__8628 (
            .O(N__40220),
            .I(\comm_spi.n22623 ));
    InMux I__8627 (
            .O(N__40213),
            .I(N__40210));
    LocalMux I__8626 (
            .O(N__40210),
            .I(N__40206));
    InMux I__8625 (
            .O(N__40209),
            .I(N__40203));
    Span4Mux_v I__8624 (
            .O(N__40206),
            .I(N__40200));
    LocalMux I__8623 (
            .O(N__40203),
            .I(N__40197));
    Odrv4 I__8622 (
            .O(N__40200),
            .I(\comm_spi.n14592 ));
    Odrv4 I__8621 (
            .O(N__40197),
            .I(\comm_spi.n14592 ));
    InMux I__8620 (
            .O(N__40192),
            .I(N__40189));
    LocalMux I__8619 (
            .O(N__40189),
            .I(N__40186));
    Span4Mux_v I__8618 (
            .O(N__40186),
            .I(N__40182));
    InMux I__8617 (
            .O(N__40185),
            .I(N__40179));
    Odrv4 I__8616 (
            .O(N__40182),
            .I(\comm_spi.n14593 ));
    LocalMux I__8615 (
            .O(N__40179),
            .I(\comm_spi.n14593 ));
    CascadeMux I__8614 (
            .O(N__40174),
            .I(N__40171));
    CascadeBuf I__8613 (
            .O(N__40171),
            .I(N__40168));
    CascadeMux I__8612 (
            .O(N__40168),
            .I(N__40165));
    CascadeBuf I__8611 (
            .O(N__40165),
            .I(N__40162));
    CascadeMux I__8610 (
            .O(N__40162),
            .I(N__40159));
    CascadeBuf I__8609 (
            .O(N__40159),
            .I(N__40156));
    CascadeMux I__8608 (
            .O(N__40156),
            .I(N__40153));
    CascadeBuf I__8607 (
            .O(N__40153),
            .I(N__40150));
    CascadeMux I__8606 (
            .O(N__40150),
            .I(N__40147));
    CascadeBuf I__8605 (
            .O(N__40147),
            .I(N__40144));
    CascadeMux I__8604 (
            .O(N__40144),
            .I(N__40141));
    CascadeBuf I__8603 (
            .O(N__40141),
            .I(N__40138));
    CascadeMux I__8602 (
            .O(N__40138),
            .I(N__40135));
    CascadeBuf I__8601 (
            .O(N__40135),
            .I(N__40132));
    CascadeMux I__8600 (
            .O(N__40132),
            .I(N__40129));
    CascadeBuf I__8599 (
            .O(N__40129),
            .I(N__40126));
    CascadeMux I__8598 (
            .O(N__40126),
            .I(N__40122));
    CascadeMux I__8597 (
            .O(N__40125),
            .I(N__40119));
    CascadeBuf I__8596 (
            .O(N__40122),
            .I(N__40116));
    CascadeBuf I__8595 (
            .O(N__40119),
            .I(N__40113));
    CascadeMux I__8594 (
            .O(N__40116),
            .I(N__40110));
    CascadeMux I__8593 (
            .O(N__40113),
            .I(N__40107));
    InMux I__8592 (
            .O(N__40110),
            .I(N__40104));
    InMux I__8591 (
            .O(N__40107),
            .I(N__40101));
    LocalMux I__8590 (
            .O(N__40104),
            .I(N__40098));
    LocalMux I__8589 (
            .O(N__40101),
            .I(N__40094));
    Span4Mux_v I__8588 (
            .O(N__40098),
            .I(N__40091));
    CascadeMux I__8587 (
            .O(N__40097),
            .I(N__40088));
    Span4Mux_v I__8586 (
            .O(N__40094),
            .I(N__40085));
    Span4Mux_h I__8585 (
            .O(N__40091),
            .I(N__40082));
    InMux I__8584 (
            .O(N__40088),
            .I(N__40079));
    Span4Mux_h I__8583 (
            .O(N__40085),
            .I(N__40074));
    Span4Mux_h I__8582 (
            .O(N__40082),
            .I(N__40074));
    LocalMux I__8581 (
            .O(N__40079),
            .I(data_count_0));
    Odrv4 I__8580 (
            .O(N__40074),
            .I(data_count_0));
    CascadeMux I__8579 (
            .O(N__40069),
            .I(N__40066));
    CascadeBuf I__8578 (
            .O(N__40066),
            .I(N__40063));
    CascadeMux I__8577 (
            .O(N__40063),
            .I(N__40060));
    CascadeBuf I__8576 (
            .O(N__40060),
            .I(N__40057));
    CascadeMux I__8575 (
            .O(N__40057),
            .I(N__40054));
    CascadeBuf I__8574 (
            .O(N__40054),
            .I(N__40051));
    CascadeMux I__8573 (
            .O(N__40051),
            .I(N__40048));
    CascadeBuf I__8572 (
            .O(N__40048),
            .I(N__40045));
    CascadeMux I__8571 (
            .O(N__40045),
            .I(N__40042));
    CascadeBuf I__8570 (
            .O(N__40042),
            .I(N__40039));
    CascadeMux I__8569 (
            .O(N__40039),
            .I(N__40036));
    CascadeBuf I__8568 (
            .O(N__40036),
            .I(N__40033));
    CascadeMux I__8567 (
            .O(N__40033),
            .I(N__40030));
    CascadeBuf I__8566 (
            .O(N__40030),
            .I(N__40027));
    CascadeMux I__8565 (
            .O(N__40027),
            .I(N__40024));
    CascadeBuf I__8564 (
            .O(N__40024),
            .I(N__40021));
    CascadeMux I__8563 (
            .O(N__40021),
            .I(N__40017));
    CascadeMux I__8562 (
            .O(N__40020),
            .I(N__40014));
    CascadeBuf I__8561 (
            .O(N__40017),
            .I(N__40011));
    CascadeBuf I__8560 (
            .O(N__40014),
            .I(N__40008));
    CascadeMux I__8559 (
            .O(N__40011),
            .I(N__40005));
    CascadeMux I__8558 (
            .O(N__40008),
            .I(N__40002));
    InMux I__8557 (
            .O(N__40005),
            .I(N__39999));
    InMux I__8556 (
            .O(N__40002),
            .I(N__39996));
    LocalMux I__8555 (
            .O(N__39999),
            .I(N__39993));
    LocalMux I__8554 (
            .O(N__39996),
            .I(N__39990));
    Span4Mux_v I__8553 (
            .O(N__39993),
            .I(N__39987));
    Span4Mux_v I__8552 (
            .O(N__39990),
            .I(N__39983));
    Span4Mux_h I__8551 (
            .O(N__39987),
            .I(N__39980));
    InMux I__8550 (
            .O(N__39986),
            .I(N__39977));
    Span4Mux_h I__8549 (
            .O(N__39983),
            .I(N__39972));
    Span4Mux_h I__8548 (
            .O(N__39980),
            .I(N__39972));
    LocalMux I__8547 (
            .O(N__39977),
            .I(data_count_1));
    Odrv4 I__8546 (
            .O(N__39972),
            .I(data_count_1));
    InMux I__8545 (
            .O(N__39967),
            .I(n19287));
    CascadeMux I__8544 (
            .O(N__39964),
            .I(N__39961));
    CascadeBuf I__8543 (
            .O(N__39961),
            .I(N__39958));
    CascadeMux I__8542 (
            .O(N__39958),
            .I(N__39955));
    CascadeBuf I__8541 (
            .O(N__39955),
            .I(N__39952));
    CascadeMux I__8540 (
            .O(N__39952),
            .I(N__39949));
    CascadeBuf I__8539 (
            .O(N__39949),
            .I(N__39946));
    CascadeMux I__8538 (
            .O(N__39946),
            .I(N__39943));
    CascadeBuf I__8537 (
            .O(N__39943),
            .I(N__39940));
    CascadeMux I__8536 (
            .O(N__39940),
            .I(N__39937));
    CascadeBuf I__8535 (
            .O(N__39937),
            .I(N__39934));
    CascadeMux I__8534 (
            .O(N__39934),
            .I(N__39931));
    CascadeBuf I__8533 (
            .O(N__39931),
            .I(N__39928));
    CascadeMux I__8532 (
            .O(N__39928),
            .I(N__39925));
    CascadeBuf I__8531 (
            .O(N__39925),
            .I(N__39922));
    CascadeMux I__8530 (
            .O(N__39922),
            .I(N__39919));
    CascadeBuf I__8529 (
            .O(N__39919),
            .I(N__39916));
    CascadeMux I__8528 (
            .O(N__39916),
            .I(N__39912));
    CascadeMux I__8527 (
            .O(N__39915),
            .I(N__39909));
    CascadeBuf I__8526 (
            .O(N__39912),
            .I(N__39906));
    CascadeBuf I__8525 (
            .O(N__39909),
            .I(N__39903));
    CascadeMux I__8524 (
            .O(N__39906),
            .I(N__39900));
    CascadeMux I__8523 (
            .O(N__39903),
            .I(N__39897));
    InMux I__8522 (
            .O(N__39900),
            .I(N__39894));
    InMux I__8521 (
            .O(N__39897),
            .I(N__39891));
    LocalMux I__8520 (
            .O(N__39894),
            .I(N__39888));
    LocalMux I__8519 (
            .O(N__39891),
            .I(N__39885));
    Span4Mux_h I__8518 (
            .O(N__39888),
            .I(N__39882));
    Span4Mux_h I__8517 (
            .O(N__39885),
            .I(N__39878));
    Span4Mux_h I__8516 (
            .O(N__39882),
            .I(N__39875));
    InMux I__8515 (
            .O(N__39881),
            .I(N__39872));
    Span4Mux_h I__8514 (
            .O(N__39878),
            .I(N__39869));
    Span4Mux_h I__8513 (
            .O(N__39875),
            .I(N__39866));
    LocalMux I__8512 (
            .O(N__39872),
            .I(data_count_2));
    Odrv4 I__8511 (
            .O(N__39869),
            .I(data_count_2));
    Odrv4 I__8510 (
            .O(N__39866),
            .I(data_count_2));
    InMux I__8509 (
            .O(N__39859),
            .I(n19288));
    CascadeMux I__8508 (
            .O(N__39856),
            .I(N__39853));
    CascadeBuf I__8507 (
            .O(N__39853),
            .I(N__39850));
    CascadeMux I__8506 (
            .O(N__39850),
            .I(N__39847));
    CascadeBuf I__8505 (
            .O(N__39847),
            .I(N__39844));
    CascadeMux I__8504 (
            .O(N__39844),
            .I(N__39841));
    CascadeBuf I__8503 (
            .O(N__39841),
            .I(N__39838));
    CascadeMux I__8502 (
            .O(N__39838),
            .I(N__39835));
    CascadeBuf I__8501 (
            .O(N__39835),
            .I(N__39832));
    CascadeMux I__8500 (
            .O(N__39832),
            .I(N__39829));
    CascadeBuf I__8499 (
            .O(N__39829),
            .I(N__39826));
    CascadeMux I__8498 (
            .O(N__39826),
            .I(N__39823));
    CascadeBuf I__8497 (
            .O(N__39823),
            .I(N__39820));
    CascadeMux I__8496 (
            .O(N__39820),
            .I(N__39817));
    CascadeBuf I__8495 (
            .O(N__39817),
            .I(N__39814));
    CascadeMux I__8494 (
            .O(N__39814),
            .I(N__39810));
    CascadeMux I__8493 (
            .O(N__39813),
            .I(N__39807));
    CascadeBuf I__8492 (
            .O(N__39810),
            .I(N__39804));
    CascadeBuf I__8491 (
            .O(N__39807),
            .I(N__39801));
    CascadeMux I__8490 (
            .O(N__39804),
            .I(N__39798));
    CascadeMux I__8489 (
            .O(N__39801),
            .I(N__39795));
    CascadeBuf I__8488 (
            .O(N__39798),
            .I(N__39792));
    InMux I__8487 (
            .O(N__39795),
            .I(N__39789));
    CascadeMux I__8486 (
            .O(N__39792),
            .I(N__39786));
    LocalMux I__8485 (
            .O(N__39789),
            .I(N__39783));
    InMux I__8484 (
            .O(N__39786),
            .I(N__39780));
    Span4Mux_h I__8483 (
            .O(N__39783),
            .I(N__39776));
    LocalMux I__8482 (
            .O(N__39780),
            .I(N__39773));
    InMux I__8481 (
            .O(N__39779),
            .I(N__39770));
    Span4Mux_h I__8480 (
            .O(N__39776),
            .I(N__39767));
    Span12Mux_h I__8479 (
            .O(N__39773),
            .I(N__39764));
    LocalMux I__8478 (
            .O(N__39770),
            .I(data_count_3));
    Odrv4 I__8477 (
            .O(N__39767),
            .I(data_count_3));
    Odrv12 I__8476 (
            .O(N__39764),
            .I(data_count_3));
    InMux I__8475 (
            .O(N__39757),
            .I(n19289));
    CascadeMux I__8474 (
            .O(N__39754),
            .I(N__39751));
    CascadeBuf I__8473 (
            .O(N__39751),
            .I(N__39748));
    CascadeMux I__8472 (
            .O(N__39748),
            .I(N__39745));
    CascadeBuf I__8471 (
            .O(N__39745),
            .I(N__39742));
    CascadeMux I__8470 (
            .O(N__39742),
            .I(N__39739));
    CascadeBuf I__8469 (
            .O(N__39739),
            .I(N__39736));
    CascadeMux I__8468 (
            .O(N__39736),
            .I(N__39733));
    CascadeBuf I__8467 (
            .O(N__39733),
            .I(N__39730));
    CascadeMux I__8466 (
            .O(N__39730),
            .I(N__39727));
    CascadeBuf I__8465 (
            .O(N__39727),
            .I(N__39724));
    CascadeMux I__8464 (
            .O(N__39724),
            .I(N__39721));
    CascadeBuf I__8463 (
            .O(N__39721),
            .I(N__39718));
    CascadeMux I__8462 (
            .O(N__39718),
            .I(N__39715));
    CascadeBuf I__8461 (
            .O(N__39715),
            .I(N__39712));
    CascadeMux I__8460 (
            .O(N__39712),
            .I(N__39709));
    CascadeBuf I__8459 (
            .O(N__39709),
            .I(N__39706));
    CascadeMux I__8458 (
            .O(N__39706),
            .I(N__39702));
    CascadeMux I__8457 (
            .O(N__39705),
            .I(N__39699));
    CascadeBuf I__8456 (
            .O(N__39702),
            .I(N__39696));
    CascadeBuf I__8455 (
            .O(N__39699),
            .I(N__39693));
    CascadeMux I__8454 (
            .O(N__39696),
            .I(N__39690));
    CascadeMux I__8453 (
            .O(N__39693),
            .I(N__39687));
    InMux I__8452 (
            .O(N__39690),
            .I(N__39684));
    InMux I__8451 (
            .O(N__39687),
            .I(N__39681));
    LocalMux I__8450 (
            .O(N__39684),
            .I(N__39678));
    LocalMux I__8449 (
            .O(N__39681),
            .I(N__39675));
    Span4Mux_h I__8448 (
            .O(N__39678),
            .I(N__39672));
    Span4Mux_v I__8447 (
            .O(N__39675),
            .I(N__39668));
    Span4Mux_h I__8446 (
            .O(N__39672),
            .I(N__39665));
    InMux I__8445 (
            .O(N__39671),
            .I(N__39662));
    Span4Mux_h I__8444 (
            .O(N__39668),
            .I(N__39659));
    Span4Mux_h I__8443 (
            .O(N__39665),
            .I(N__39656));
    LocalMux I__8442 (
            .O(N__39662),
            .I(data_count_4));
    Odrv4 I__8441 (
            .O(N__39659),
            .I(data_count_4));
    Odrv4 I__8440 (
            .O(N__39656),
            .I(data_count_4));
    InMux I__8439 (
            .O(N__39649),
            .I(n19290));
    CascadeMux I__8438 (
            .O(N__39646),
            .I(N__39643));
    CascadeBuf I__8437 (
            .O(N__39643),
            .I(N__39640));
    CascadeMux I__8436 (
            .O(N__39640),
            .I(N__39637));
    CascadeBuf I__8435 (
            .O(N__39637),
            .I(N__39634));
    CascadeMux I__8434 (
            .O(N__39634),
            .I(N__39631));
    CascadeBuf I__8433 (
            .O(N__39631),
            .I(N__39628));
    CascadeMux I__8432 (
            .O(N__39628),
            .I(N__39625));
    CascadeBuf I__8431 (
            .O(N__39625),
            .I(N__39622));
    CascadeMux I__8430 (
            .O(N__39622),
            .I(N__39619));
    CascadeBuf I__8429 (
            .O(N__39619),
            .I(N__39616));
    CascadeMux I__8428 (
            .O(N__39616),
            .I(N__39613));
    CascadeBuf I__8427 (
            .O(N__39613),
            .I(N__39610));
    CascadeMux I__8426 (
            .O(N__39610),
            .I(N__39607));
    CascadeBuf I__8425 (
            .O(N__39607),
            .I(N__39604));
    CascadeMux I__8424 (
            .O(N__39604),
            .I(N__39601));
    CascadeBuf I__8423 (
            .O(N__39601),
            .I(N__39598));
    CascadeMux I__8422 (
            .O(N__39598),
            .I(N__39594));
    CascadeMux I__8421 (
            .O(N__39597),
            .I(N__39591));
    CascadeBuf I__8420 (
            .O(N__39594),
            .I(N__39588));
    CascadeBuf I__8419 (
            .O(N__39591),
            .I(N__39585));
    CascadeMux I__8418 (
            .O(N__39588),
            .I(N__39582));
    CascadeMux I__8417 (
            .O(N__39585),
            .I(N__39579));
    InMux I__8416 (
            .O(N__39582),
            .I(N__39576));
    InMux I__8415 (
            .O(N__39579),
            .I(N__39573));
    LocalMux I__8414 (
            .O(N__39576),
            .I(N__39570));
    LocalMux I__8413 (
            .O(N__39573),
            .I(N__39567));
    Span4Mux_h I__8412 (
            .O(N__39570),
            .I(N__39564));
    Span4Mux_v I__8411 (
            .O(N__39567),
            .I(N__39560));
    Span4Mux_h I__8410 (
            .O(N__39564),
            .I(N__39557));
    InMux I__8409 (
            .O(N__39563),
            .I(N__39554));
    Span4Mux_h I__8408 (
            .O(N__39560),
            .I(N__39551));
    Span4Mux_h I__8407 (
            .O(N__39557),
            .I(N__39548));
    LocalMux I__8406 (
            .O(N__39554),
            .I(data_count_5));
    Odrv4 I__8405 (
            .O(N__39551),
            .I(data_count_5));
    Odrv4 I__8404 (
            .O(N__39548),
            .I(data_count_5));
    InMux I__8403 (
            .O(N__39541),
            .I(n19291));
    CascadeMux I__8402 (
            .O(N__39538),
            .I(N__39535));
    CascadeBuf I__8401 (
            .O(N__39535),
            .I(N__39532));
    CascadeMux I__8400 (
            .O(N__39532),
            .I(N__39529));
    CascadeBuf I__8399 (
            .O(N__39529),
            .I(N__39526));
    CascadeMux I__8398 (
            .O(N__39526),
            .I(N__39523));
    CascadeBuf I__8397 (
            .O(N__39523),
            .I(N__39520));
    CascadeMux I__8396 (
            .O(N__39520),
            .I(N__39517));
    CascadeBuf I__8395 (
            .O(N__39517),
            .I(N__39514));
    CascadeMux I__8394 (
            .O(N__39514),
            .I(N__39511));
    CascadeBuf I__8393 (
            .O(N__39511),
            .I(N__39508));
    CascadeMux I__8392 (
            .O(N__39508),
            .I(N__39505));
    CascadeBuf I__8391 (
            .O(N__39505),
            .I(N__39502));
    CascadeMux I__8390 (
            .O(N__39502),
            .I(N__39499));
    CascadeBuf I__8389 (
            .O(N__39499),
            .I(N__39496));
    CascadeMux I__8388 (
            .O(N__39496),
            .I(N__39493));
    CascadeBuf I__8387 (
            .O(N__39493),
            .I(N__39489));
    CascadeMux I__8386 (
            .O(N__39492),
            .I(N__39486));
    CascadeMux I__8385 (
            .O(N__39489),
            .I(N__39483));
    CascadeBuf I__8384 (
            .O(N__39486),
            .I(N__39480));
    CascadeBuf I__8383 (
            .O(N__39483),
            .I(N__39477));
    CascadeMux I__8382 (
            .O(N__39480),
            .I(N__39474));
    CascadeMux I__8381 (
            .O(N__39477),
            .I(N__39471));
    InMux I__8380 (
            .O(N__39474),
            .I(N__39468));
    InMux I__8379 (
            .O(N__39471),
            .I(N__39465));
    LocalMux I__8378 (
            .O(N__39468),
            .I(N__39462));
    LocalMux I__8377 (
            .O(N__39465),
            .I(N__39459));
    Span4Mux_h I__8376 (
            .O(N__39462),
            .I(N__39455));
    Span4Mux_v I__8375 (
            .O(N__39459),
            .I(N__39452));
    InMux I__8374 (
            .O(N__39458),
            .I(N__39449));
    Span4Mux_h I__8373 (
            .O(N__39455),
            .I(N__39446));
    Sp12to4 I__8372 (
            .O(N__39452),
            .I(N__39443));
    LocalMux I__8371 (
            .O(N__39449),
            .I(data_count_6));
    Odrv4 I__8370 (
            .O(N__39446),
            .I(data_count_6));
    Odrv12 I__8369 (
            .O(N__39443),
            .I(data_count_6));
    InMux I__8368 (
            .O(N__39436),
            .I(n19292));
    CascadeMux I__8367 (
            .O(N__39433),
            .I(N__39430));
    CascadeBuf I__8366 (
            .O(N__39430),
            .I(N__39427));
    CascadeMux I__8365 (
            .O(N__39427),
            .I(N__39424));
    CascadeBuf I__8364 (
            .O(N__39424),
            .I(N__39421));
    CascadeMux I__8363 (
            .O(N__39421),
            .I(N__39418));
    CascadeBuf I__8362 (
            .O(N__39418),
            .I(N__39415));
    CascadeMux I__8361 (
            .O(N__39415),
            .I(N__39412));
    CascadeBuf I__8360 (
            .O(N__39412),
            .I(N__39409));
    CascadeMux I__8359 (
            .O(N__39409),
            .I(N__39406));
    CascadeBuf I__8358 (
            .O(N__39406),
            .I(N__39403));
    CascadeMux I__8357 (
            .O(N__39403),
            .I(N__39400));
    CascadeBuf I__8356 (
            .O(N__39400),
            .I(N__39397));
    CascadeMux I__8355 (
            .O(N__39397),
            .I(N__39394));
    CascadeBuf I__8354 (
            .O(N__39394),
            .I(N__39391));
    CascadeMux I__8353 (
            .O(N__39391),
            .I(N__39387));
    CascadeMux I__8352 (
            .O(N__39390),
            .I(N__39384));
    CascadeBuf I__8351 (
            .O(N__39387),
            .I(N__39381));
    CascadeBuf I__8350 (
            .O(N__39384),
            .I(N__39378));
    CascadeMux I__8349 (
            .O(N__39381),
            .I(N__39375));
    CascadeMux I__8348 (
            .O(N__39378),
            .I(N__39372));
    CascadeBuf I__8347 (
            .O(N__39375),
            .I(N__39369));
    InMux I__8346 (
            .O(N__39372),
            .I(N__39366));
    CascadeMux I__8345 (
            .O(N__39369),
            .I(N__39363));
    LocalMux I__8344 (
            .O(N__39366),
            .I(N__39360));
    InMux I__8343 (
            .O(N__39363),
            .I(N__39357));
    Span4Mux_v I__8342 (
            .O(N__39360),
            .I(N__39353));
    LocalMux I__8341 (
            .O(N__39357),
            .I(N__39350));
    InMux I__8340 (
            .O(N__39356),
            .I(N__39347));
    Span4Mux_h I__8339 (
            .O(N__39353),
            .I(N__39344));
    Span12Mux_s9_v I__8338 (
            .O(N__39350),
            .I(N__39341));
    LocalMux I__8337 (
            .O(N__39347),
            .I(data_count_7));
    Odrv4 I__8336 (
            .O(N__39344),
            .I(data_count_7));
    Odrv12 I__8335 (
            .O(N__39341),
            .I(data_count_7));
    InMux I__8334 (
            .O(N__39334),
            .I(n19293));
    CascadeMux I__8333 (
            .O(N__39331),
            .I(N__39324));
    InMux I__8332 (
            .O(N__39330),
            .I(N__39318));
    InMux I__8331 (
            .O(N__39329),
            .I(N__39318));
    InMux I__8330 (
            .O(N__39328),
            .I(N__39308));
    InMux I__8329 (
            .O(N__39327),
            .I(N__39308));
    InMux I__8328 (
            .O(N__39324),
            .I(N__39303));
    InMux I__8327 (
            .O(N__39323),
            .I(N__39303));
    LocalMux I__8326 (
            .O(N__39318),
            .I(N__39300));
    InMux I__8325 (
            .O(N__39317),
            .I(N__39293));
    InMux I__8324 (
            .O(N__39316),
            .I(N__39293));
    InMux I__8323 (
            .O(N__39315),
            .I(N__39293));
    InMux I__8322 (
            .O(N__39314),
            .I(N__39288));
    InMux I__8321 (
            .O(N__39313),
            .I(N__39288));
    LocalMux I__8320 (
            .O(N__39308),
            .I(N__39280));
    LocalMux I__8319 (
            .O(N__39303),
            .I(N__39280));
    Span4Mux_v I__8318 (
            .O(N__39300),
            .I(N__39277));
    LocalMux I__8317 (
            .O(N__39293),
            .I(N__39274));
    LocalMux I__8316 (
            .O(N__39288),
            .I(N__39269));
    InMux I__8315 (
            .O(N__39287),
            .I(N__39262));
    InMux I__8314 (
            .O(N__39286),
            .I(N__39262));
    InMux I__8313 (
            .O(N__39285),
            .I(N__39262));
    Span4Mux_h I__8312 (
            .O(N__39280),
            .I(N__39255));
    Span4Mux_h I__8311 (
            .O(N__39277),
            .I(N__39255));
    Span4Mux_h I__8310 (
            .O(N__39274),
            .I(N__39255));
    InMux I__8309 (
            .O(N__39273),
            .I(N__39250));
    InMux I__8308 (
            .O(N__39272),
            .I(N__39250));
    Odrv4 I__8307 (
            .O(N__39269),
            .I(n12391));
    LocalMux I__8306 (
            .O(N__39262),
            .I(n12391));
    Odrv4 I__8305 (
            .O(N__39255),
            .I(n12391));
    LocalMux I__8304 (
            .O(N__39250),
            .I(n12391));
    InMux I__8303 (
            .O(N__39241),
            .I(N__39233));
    InMux I__8302 (
            .O(N__39240),
            .I(N__39226));
    InMux I__8301 (
            .O(N__39239),
            .I(N__39226));
    InMux I__8300 (
            .O(N__39238),
            .I(N__39226));
    InMux I__8299 (
            .O(N__39237),
            .I(N__39223));
    InMux I__8298 (
            .O(N__39236),
            .I(N__39220));
    LocalMux I__8297 (
            .O(N__39233),
            .I(N__39212));
    LocalMux I__8296 (
            .O(N__39226),
            .I(N__39212));
    LocalMux I__8295 (
            .O(N__39223),
            .I(N__39212));
    LocalMux I__8294 (
            .O(N__39220),
            .I(N__39209));
    InMux I__8293 (
            .O(N__39219),
            .I(N__39206));
    Span4Mux_v I__8292 (
            .O(N__39212),
            .I(N__39198));
    Span4Mux_h I__8291 (
            .O(N__39209),
            .I(N__39198));
    LocalMux I__8290 (
            .O(N__39206),
            .I(N__39198));
    InMux I__8289 (
            .O(N__39205),
            .I(N__39195));
    Sp12to4 I__8288 (
            .O(N__39198),
            .I(N__39190));
    LocalMux I__8287 (
            .O(N__39195),
            .I(N__39190));
    Odrv12 I__8286 (
            .O(N__39190),
            .I(n12367));
    InMux I__8285 (
            .O(N__39187),
            .I(N__39184));
    LocalMux I__8284 (
            .O(N__39184),
            .I(N__39180));
    CascadeMux I__8283 (
            .O(N__39183),
            .I(N__39177));
    Span4Mux_v I__8282 (
            .O(N__39180),
            .I(N__39174));
    InMux I__8281 (
            .O(N__39177),
            .I(N__39171));
    Span4Mux_h I__8280 (
            .O(N__39174),
            .I(N__39168));
    LocalMux I__8279 (
            .O(N__39171),
            .I(N__39165));
    Odrv4 I__8278 (
            .O(N__39168),
            .I(n11324));
    Odrv12 I__8277 (
            .O(N__39165),
            .I(n11324));
    CascadeMux I__8276 (
            .O(N__39160),
            .I(n8780_cascade_));
    CascadeMux I__8275 (
            .O(N__39157),
            .I(N__39153));
    InMux I__8274 (
            .O(N__39156),
            .I(N__39143));
    InMux I__8273 (
            .O(N__39153),
            .I(N__39143));
    InMux I__8272 (
            .O(N__39152),
            .I(N__39143));
    CascadeMux I__8271 (
            .O(N__39151),
            .I(N__39138));
    InMux I__8270 (
            .O(N__39150),
            .I(N__39134));
    LocalMux I__8269 (
            .O(N__39143),
            .I(N__39131));
    InMux I__8268 (
            .O(N__39142),
            .I(N__39128));
    InMux I__8267 (
            .O(N__39141),
            .I(N__39123));
    InMux I__8266 (
            .O(N__39138),
            .I(N__39123));
    InMux I__8265 (
            .O(N__39137),
            .I(N__39119));
    LocalMux I__8264 (
            .O(N__39134),
            .I(N__39116));
    Span4Mux_v I__8263 (
            .O(N__39131),
            .I(N__39109));
    LocalMux I__8262 (
            .O(N__39128),
            .I(N__39109));
    LocalMux I__8261 (
            .O(N__39123),
            .I(N__39109));
    CascadeMux I__8260 (
            .O(N__39122),
            .I(N__39102));
    LocalMux I__8259 (
            .O(N__39119),
            .I(N__39099));
    Span4Mux_v I__8258 (
            .O(N__39116),
            .I(N__39094));
    Span4Mux_v I__8257 (
            .O(N__39109),
            .I(N__39094));
    InMux I__8256 (
            .O(N__39108),
            .I(N__39089));
    InMux I__8255 (
            .O(N__39107),
            .I(N__39089));
    InMux I__8254 (
            .O(N__39106),
            .I(N__39086));
    InMux I__8253 (
            .O(N__39105),
            .I(N__39081));
    InMux I__8252 (
            .O(N__39102),
            .I(N__39081));
    Span4Mux_v I__8251 (
            .O(N__39099),
            .I(N__39076));
    Span4Mux_h I__8250 (
            .O(N__39094),
            .I(N__39076));
    LocalMux I__8249 (
            .O(N__39089),
            .I(N__39073));
    LocalMux I__8248 (
            .O(N__39086),
            .I(eis_state_1));
    LocalMux I__8247 (
            .O(N__39081),
            .I(eis_state_1));
    Odrv4 I__8246 (
            .O(N__39076),
            .I(eis_state_1));
    Odrv12 I__8245 (
            .O(N__39073),
            .I(eis_state_1));
    InMux I__8244 (
            .O(N__39064),
            .I(N__39058));
    InMux I__8243 (
            .O(N__39063),
            .I(N__39058));
    LocalMux I__8242 (
            .O(N__39058),
            .I(N__39054));
    InMux I__8241 (
            .O(N__39057),
            .I(N__39051));
    Span4Mux_h I__8240 (
            .O(N__39054),
            .I(N__39048));
    LocalMux I__8239 (
            .O(N__39051),
            .I(buf_dds0_7));
    Odrv4 I__8238 (
            .O(N__39048),
            .I(buf_dds0_7));
    InMux I__8237 (
            .O(N__39043),
            .I(N__39040));
    LocalMux I__8236 (
            .O(N__39040),
            .I(n8_adj_1541));
    CascadeMux I__8235 (
            .O(N__39037),
            .I(n8_adj_1541_cascade_));
    CascadeMux I__8234 (
            .O(N__39034),
            .I(N__39031));
    CascadeBuf I__8233 (
            .O(N__39031),
            .I(N__39028));
    CascadeMux I__8232 (
            .O(N__39028),
            .I(N__39025));
    CascadeBuf I__8231 (
            .O(N__39025),
            .I(N__39022));
    CascadeMux I__8230 (
            .O(N__39022),
            .I(N__39019));
    CascadeBuf I__8229 (
            .O(N__39019),
            .I(N__39016));
    CascadeMux I__8228 (
            .O(N__39016),
            .I(N__39013));
    CascadeBuf I__8227 (
            .O(N__39013),
            .I(N__39010));
    CascadeMux I__8226 (
            .O(N__39010),
            .I(N__39007));
    CascadeBuf I__8225 (
            .O(N__39007),
            .I(N__39004));
    CascadeMux I__8224 (
            .O(N__39004),
            .I(N__39001));
    CascadeBuf I__8223 (
            .O(N__39001),
            .I(N__38998));
    CascadeMux I__8222 (
            .O(N__38998),
            .I(N__38995));
    CascadeBuf I__8221 (
            .O(N__38995),
            .I(N__38992));
    CascadeMux I__8220 (
            .O(N__38992),
            .I(N__38988));
    CascadeMux I__8219 (
            .O(N__38991),
            .I(N__38985));
    CascadeBuf I__8218 (
            .O(N__38988),
            .I(N__38982));
    CascadeBuf I__8217 (
            .O(N__38985),
            .I(N__38979));
    CascadeMux I__8216 (
            .O(N__38982),
            .I(N__38976));
    CascadeMux I__8215 (
            .O(N__38979),
            .I(N__38973));
    CascadeBuf I__8214 (
            .O(N__38976),
            .I(N__38970));
    InMux I__8213 (
            .O(N__38973),
            .I(N__38967));
    CascadeMux I__8212 (
            .O(N__38970),
            .I(N__38964));
    LocalMux I__8211 (
            .O(N__38967),
            .I(N__38961));
    InMux I__8210 (
            .O(N__38964),
            .I(N__38958));
    Span4Mux_h I__8209 (
            .O(N__38961),
            .I(N__38955));
    LocalMux I__8208 (
            .O(N__38958),
            .I(N__38952));
    Span4Mux_h I__8207 (
            .O(N__38955),
            .I(N__38949));
    Span12Mux_s10_v I__8206 (
            .O(N__38952),
            .I(N__38946));
    Odrv4 I__8205 (
            .O(N__38949),
            .I(data_index_9_N_212_4));
    Odrv12 I__8204 (
            .O(N__38946),
            .I(data_index_9_N_212_4));
    InMux I__8203 (
            .O(N__38941),
            .I(N__38938));
    LocalMux I__8202 (
            .O(N__38938),
            .I(N__38932));
    InMux I__8201 (
            .O(N__38937),
            .I(N__38929));
    InMux I__8200 (
            .O(N__38936),
            .I(N__38926));
    InMux I__8199 (
            .O(N__38935),
            .I(N__38923));
    Span4Mux_h I__8198 (
            .O(N__38932),
            .I(N__38920));
    LocalMux I__8197 (
            .O(N__38929),
            .I(N__38917));
    LocalMux I__8196 (
            .O(N__38926),
            .I(N__38914));
    LocalMux I__8195 (
            .O(N__38923),
            .I(N__38907));
    Span4Mux_v I__8194 (
            .O(N__38920),
            .I(N__38907));
    Span4Mux_h I__8193 (
            .O(N__38917),
            .I(N__38907));
    Odrv4 I__8192 (
            .O(N__38914),
            .I(eis_stop));
    Odrv4 I__8191 (
            .O(N__38907),
            .I(eis_stop));
    CascadeMux I__8190 (
            .O(N__38902),
            .I(n29_cascade_));
    InMux I__8189 (
            .O(N__38899),
            .I(N__38894));
    InMux I__8188 (
            .O(N__38898),
            .I(N__38891));
    InMux I__8187 (
            .O(N__38897),
            .I(N__38888));
    LocalMux I__8186 (
            .O(N__38894),
            .I(N__38885));
    LocalMux I__8185 (
            .O(N__38891),
            .I(N__38882));
    LocalMux I__8184 (
            .O(N__38888),
            .I(N__38879));
    Span4Mux_h I__8183 (
            .O(N__38885),
            .I(N__38874));
    Span4Mux_h I__8182 (
            .O(N__38882),
            .I(N__38874));
    Odrv12 I__8181 (
            .O(N__38879),
            .I(n16_adj_1609));
    Odrv4 I__8180 (
            .O(N__38874),
            .I(n16_adj_1609));
    CascadeMux I__8179 (
            .O(N__38869),
            .I(N__38866));
    InMux I__8178 (
            .O(N__38866),
            .I(N__38862));
    InMux I__8177 (
            .O(N__38865),
            .I(N__38859));
    LocalMux I__8176 (
            .O(N__38862),
            .I(N__38856));
    LocalMux I__8175 (
            .O(N__38859),
            .I(N__38852));
    Span4Mux_h I__8174 (
            .O(N__38856),
            .I(N__38849));
    InMux I__8173 (
            .O(N__38855),
            .I(N__38846));
    Span4Mux_v I__8172 (
            .O(N__38852),
            .I(N__38843));
    Span4Mux_v I__8171 (
            .O(N__38849),
            .I(N__38838));
    LocalMux I__8170 (
            .O(N__38846),
            .I(N__38838));
    Odrv4 I__8169 (
            .O(N__38843),
            .I(n14_adj_1558));
    Odrv4 I__8168 (
            .O(N__38838),
            .I(n14_adj_1558));
    InMux I__8167 (
            .O(N__38833),
            .I(N__38830));
    LocalMux I__8166 (
            .O(N__38830),
            .I(N__38827));
    Span4Mux_h I__8165 (
            .O(N__38827),
            .I(N__38822));
    InMux I__8164 (
            .O(N__38826),
            .I(N__38817));
    InMux I__8163 (
            .O(N__38825),
            .I(N__38817));
    Odrv4 I__8162 (
            .O(N__38822),
            .I(req_data_cnt_3));
    LocalMux I__8161 (
            .O(N__38817),
            .I(req_data_cnt_3));
    InMux I__8160 (
            .O(N__38812),
            .I(N__38809));
    LocalMux I__8159 (
            .O(N__38809),
            .I(N__38805));
    InMux I__8158 (
            .O(N__38808),
            .I(N__38802));
    Span4Mux_h I__8157 (
            .O(N__38805),
            .I(N__38799));
    LocalMux I__8156 (
            .O(N__38802),
            .I(acadc_skipcnt_12));
    Odrv4 I__8155 (
            .O(N__38799),
            .I(acadc_skipcnt_12));
    InMux I__8154 (
            .O(N__38794),
            .I(N__38791));
    LocalMux I__8153 (
            .O(N__38791),
            .I(N__38787));
    InMux I__8152 (
            .O(N__38790),
            .I(N__38784));
    Span4Mux_h I__8151 (
            .O(N__38787),
            .I(N__38781));
    LocalMux I__8150 (
            .O(N__38784),
            .I(acadc_skipcnt_10));
    Odrv4 I__8149 (
            .O(N__38781),
            .I(acadc_skipcnt_10));
    InMux I__8148 (
            .O(N__38776),
            .I(N__38773));
    LocalMux I__8147 (
            .O(N__38773),
            .I(n21));
    CascadeMux I__8146 (
            .O(N__38770),
            .I(n9_adj_1408_cascade_));
    InMux I__8145 (
            .O(N__38767),
            .I(N__38764));
    LocalMux I__8144 (
            .O(N__38764),
            .I(N__38760));
    CascadeMux I__8143 (
            .O(N__38763),
            .I(N__38756));
    Span4Mux_v I__8142 (
            .O(N__38760),
            .I(N__38753));
    CascadeMux I__8141 (
            .O(N__38759),
            .I(N__38750));
    InMux I__8140 (
            .O(N__38756),
            .I(N__38747));
    Span4Mux_h I__8139 (
            .O(N__38753),
            .I(N__38744));
    InMux I__8138 (
            .O(N__38750),
            .I(N__38741));
    LocalMux I__8137 (
            .O(N__38747),
            .I(cmd_rdadctmp_14_adj_1429));
    Odrv4 I__8136 (
            .O(N__38744),
            .I(cmd_rdadctmp_14_adj_1429));
    LocalMux I__8135 (
            .O(N__38741),
            .I(cmd_rdadctmp_14_adj_1429));
    CascadeMux I__8134 (
            .O(N__38734),
            .I(N__38726));
    CascadeMux I__8133 (
            .O(N__38733),
            .I(N__38723));
    CascadeMux I__8132 (
            .O(N__38732),
            .I(N__38720));
    CascadeMux I__8131 (
            .O(N__38731),
            .I(N__38716));
    CascadeMux I__8130 (
            .O(N__38730),
            .I(N__38713));
    CascadeMux I__8129 (
            .O(N__38729),
            .I(N__38709));
    InMux I__8128 (
            .O(N__38726),
            .I(N__38706));
    InMux I__8127 (
            .O(N__38723),
            .I(N__38703));
    InMux I__8126 (
            .O(N__38720),
            .I(N__38700));
    InMux I__8125 (
            .O(N__38719),
            .I(N__38697));
    InMux I__8124 (
            .O(N__38716),
            .I(N__38694));
    InMux I__8123 (
            .O(N__38713),
            .I(N__38691));
    InMux I__8122 (
            .O(N__38712),
            .I(N__38688));
    InMux I__8121 (
            .O(N__38709),
            .I(N__38685));
    LocalMux I__8120 (
            .O(N__38706),
            .I(N__38682));
    LocalMux I__8119 (
            .O(N__38703),
            .I(N__38679));
    LocalMux I__8118 (
            .O(N__38700),
            .I(N__38676));
    LocalMux I__8117 (
            .O(N__38697),
            .I(N__38673));
    LocalMux I__8116 (
            .O(N__38694),
            .I(N__38668));
    LocalMux I__8115 (
            .O(N__38691),
            .I(N__38668));
    LocalMux I__8114 (
            .O(N__38688),
            .I(N__38665));
    LocalMux I__8113 (
            .O(N__38685),
            .I(N__38662));
    Span4Mux_v I__8112 (
            .O(N__38682),
            .I(N__38659));
    Span4Mux_v I__8111 (
            .O(N__38679),
            .I(N__38654));
    Span4Mux_h I__8110 (
            .O(N__38676),
            .I(N__38654));
    Span4Mux_h I__8109 (
            .O(N__38673),
            .I(N__38651));
    Span4Mux_v I__8108 (
            .O(N__38668),
            .I(N__38645));
    Span4Mux_h I__8107 (
            .O(N__38665),
            .I(N__38645));
    Span12Mux_v I__8106 (
            .O(N__38662),
            .I(N__38640));
    Sp12to4 I__8105 (
            .O(N__38659),
            .I(N__38640));
    Span4Mux_v I__8104 (
            .O(N__38654),
            .I(N__38635));
    Span4Mux_h I__8103 (
            .O(N__38651),
            .I(N__38635));
    InMux I__8102 (
            .O(N__38650),
            .I(N__38632));
    Odrv4 I__8101 (
            .O(N__38645),
            .I(comm_buf_0_2));
    Odrv12 I__8100 (
            .O(N__38640),
            .I(comm_buf_0_2));
    Odrv4 I__8099 (
            .O(N__38635),
            .I(comm_buf_0_2));
    LocalMux I__8098 (
            .O(N__38632),
            .I(comm_buf_0_2));
    InMux I__8097 (
            .O(N__38623),
            .I(N__38620));
    LocalMux I__8096 (
            .O(N__38620),
            .I(N__38617));
    Span4Mux_h I__8095 (
            .O(N__38617),
            .I(N__38614));
    Span4Mux_h I__8094 (
            .O(N__38614),
            .I(N__38609));
    CascadeMux I__8093 (
            .O(N__38613),
            .I(N__38606));
    InMux I__8092 (
            .O(N__38612),
            .I(N__38603));
    Span4Mux_v I__8091 (
            .O(N__38609),
            .I(N__38600));
    InMux I__8090 (
            .O(N__38606),
            .I(N__38597));
    LocalMux I__8089 (
            .O(N__38603),
            .I(acadc_skipCount_10));
    Odrv4 I__8088 (
            .O(N__38600),
            .I(acadc_skipCount_10));
    LocalMux I__8087 (
            .O(N__38597),
            .I(acadc_skipCount_10));
    InMux I__8086 (
            .O(N__38590),
            .I(N__38587));
    LocalMux I__8085 (
            .O(N__38587),
            .I(N__38584));
    Odrv4 I__8084 (
            .O(N__38584),
            .I(n14_adj_1550));
    CEMux I__8083 (
            .O(N__38581),
            .I(N__38577));
    CEMux I__8082 (
            .O(N__38580),
            .I(N__38574));
    LocalMux I__8081 (
            .O(N__38577),
            .I(N__38571));
    LocalMux I__8080 (
            .O(N__38574),
            .I(N__38568));
    Span4Mux_h I__8079 (
            .O(N__38571),
            .I(N__38565));
    Span4Mux_h I__8078 (
            .O(N__38568),
            .I(N__38562));
    Odrv4 I__8077 (
            .O(N__38565),
            .I(n12254));
    Odrv4 I__8076 (
            .O(N__38562),
            .I(n12254));
    CEMux I__8075 (
            .O(N__38557),
            .I(N__38554));
    LocalMux I__8074 (
            .O(N__38554),
            .I(N__38551));
    Span4Mux_v I__8073 (
            .O(N__38551),
            .I(N__38547));
    CEMux I__8072 (
            .O(N__38550),
            .I(N__38541));
    Span4Mux_h I__8071 (
            .O(N__38547),
            .I(N__38537));
    CEMux I__8070 (
            .O(N__38546),
            .I(N__38534));
    CEMux I__8069 (
            .O(N__38545),
            .I(N__38530));
    CEMux I__8068 (
            .O(N__38544),
            .I(N__38527));
    LocalMux I__8067 (
            .O(N__38541),
            .I(N__38524));
    CEMux I__8066 (
            .O(N__38540),
            .I(N__38520));
    Span4Mux_h I__8065 (
            .O(N__38537),
            .I(N__38515));
    LocalMux I__8064 (
            .O(N__38534),
            .I(N__38515));
    CEMux I__8063 (
            .O(N__38533),
            .I(N__38512));
    LocalMux I__8062 (
            .O(N__38530),
            .I(N__38509));
    LocalMux I__8061 (
            .O(N__38527),
            .I(N__38504));
    Span4Mux_v I__8060 (
            .O(N__38524),
            .I(N__38504));
    CEMux I__8059 (
            .O(N__38523),
            .I(N__38501));
    LocalMux I__8058 (
            .O(N__38520),
            .I(N__38498));
    Span4Mux_h I__8057 (
            .O(N__38515),
            .I(N__38494));
    LocalMux I__8056 (
            .O(N__38512),
            .I(N__38487));
    Span4Mux_v I__8055 (
            .O(N__38509),
            .I(N__38487));
    Span4Mux_h I__8054 (
            .O(N__38504),
            .I(N__38487));
    LocalMux I__8053 (
            .O(N__38501),
            .I(N__38482));
    Span4Mux_v I__8052 (
            .O(N__38498),
            .I(N__38482));
    InMux I__8051 (
            .O(N__38497),
            .I(N__38479));
    Odrv4 I__8050 (
            .O(N__38494),
            .I(n12007));
    Odrv4 I__8049 (
            .O(N__38487),
            .I(n12007));
    Odrv4 I__8048 (
            .O(N__38482),
            .I(n12007));
    LocalMux I__8047 (
            .O(N__38479),
            .I(n12007));
    InMux I__8046 (
            .O(N__38470),
            .I(N__38466));
    InMux I__8045 (
            .O(N__38469),
            .I(N__38463));
    LocalMux I__8044 (
            .O(N__38466),
            .I(N__38460));
    LocalMux I__8043 (
            .O(N__38463),
            .I(N__38457));
    Span4Mux_v I__8042 (
            .O(N__38460),
            .I(N__38454));
    Span4Mux_h I__8041 (
            .O(N__38457),
            .I(N__38451));
    Span4Mux_h I__8040 (
            .O(N__38454),
            .I(N__38446));
    Span4Mux_v I__8039 (
            .O(N__38451),
            .I(N__38446));
    Odrv4 I__8038 (
            .O(N__38446),
            .I(n14_adj_1527));
    InMux I__8037 (
            .O(N__38443),
            .I(N__38439));
    InMux I__8036 (
            .O(N__38442),
            .I(N__38436));
    LocalMux I__8035 (
            .O(N__38439),
            .I(N__38433));
    LocalMux I__8034 (
            .O(N__38436),
            .I(N__38430));
    Span4Mux_h I__8033 (
            .O(N__38433),
            .I(N__38427));
    Odrv12 I__8032 (
            .O(N__38430),
            .I(n14_adj_1529));
    Odrv4 I__8031 (
            .O(N__38427),
            .I(n14_adj_1529));
    InMux I__8030 (
            .O(N__38422),
            .I(N__38419));
    LocalMux I__8029 (
            .O(N__38419),
            .I(N__38414));
    CascadeMux I__8028 (
            .O(N__38418),
            .I(N__38411));
    InMux I__8027 (
            .O(N__38417),
            .I(N__38408));
    Span4Mux_h I__8026 (
            .O(N__38414),
            .I(N__38405));
    InMux I__8025 (
            .O(N__38411),
            .I(N__38402));
    LocalMux I__8024 (
            .O(N__38408),
            .I(req_data_cnt_5));
    Odrv4 I__8023 (
            .O(N__38405),
            .I(req_data_cnt_5));
    LocalMux I__8022 (
            .O(N__38402),
            .I(req_data_cnt_5));
    InMux I__8021 (
            .O(N__38395),
            .I(N__38391));
    CascadeMux I__8020 (
            .O(N__38394),
            .I(N__38387));
    LocalMux I__8019 (
            .O(N__38391),
            .I(N__38384));
    InMux I__8018 (
            .O(N__38390),
            .I(N__38379));
    InMux I__8017 (
            .O(N__38387),
            .I(N__38379));
    Odrv4 I__8016 (
            .O(N__38384),
            .I(req_data_cnt_4));
    LocalMux I__8015 (
            .O(N__38379),
            .I(req_data_cnt_4));
    InMux I__8014 (
            .O(N__38374),
            .I(N__38369));
    InMux I__8013 (
            .O(N__38373),
            .I(N__38364));
    InMux I__8012 (
            .O(N__38372),
            .I(N__38364));
    LocalMux I__8011 (
            .O(N__38369),
            .I(req_data_cnt_1));
    LocalMux I__8010 (
            .O(N__38364),
            .I(req_data_cnt_1));
    InMux I__8009 (
            .O(N__38359),
            .I(N__38356));
    LocalMux I__8008 (
            .O(N__38356),
            .I(n20_adj_1496));
    CascadeMux I__8007 (
            .O(N__38353),
            .I(n18_adj_1553_cascade_));
    SRMux I__8006 (
            .O(N__38350),
            .I(N__38347));
    LocalMux I__8005 (
            .O(N__38347),
            .I(N__38343));
    SRMux I__8004 (
            .O(N__38346),
            .I(N__38340));
    Span4Mux_h I__8003 (
            .O(N__38343),
            .I(N__38337));
    LocalMux I__8002 (
            .O(N__38340),
            .I(N__38334));
    Odrv4 I__8001 (
            .O(N__38337),
            .I(n14749));
    Odrv12 I__8000 (
            .O(N__38334),
            .I(n14749));
    InMux I__7999 (
            .O(N__38329),
            .I(N__38326));
    LocalMux I__7998 (
            .O(N__38326),
            .I(N__38323));
    Span4Mux_v I__7997 (
            .O(N__38323),
            .I(N__38320));
    Span4Mux_h I__7996 (
            .O(N__38320),
            .I(N__38316));
    InMux I__7995 (
            .O(N__38319),
            .I(N__38313));
    Odrv4 I__7994 (
            .O(N__38316),
            .I(buf_adcdata_vdc_5));
    LocalMux I__7993 (
            .O(N__38313),
            .I(buf_adcdata_vdc_5));
    InMux I__7992 (
            .O(N__38308),
            .I(N__38305));
    LocalMux I__7991 (
            .O(N__38305),
            .I(N__38300));
    CascadeMux I__7990 (
            .O(N__38304),
            .I(N__38297));
    InMux I__7989 (
            .O(N__38303),
            .I(N__38294));
    Span4Mux_v I__7988 (
            .O(N__38300),
            .I(N__38291));
    InMux I__7987 (
            .O(N__38297),
            .I(N__38288));
    LocalMux I__7986 (
            .O(N__38294),
            .I(N__38285));
    Span4Mux_h I__7985 (
            .O(N__38291),
            .I(N__38282));
    LocalMux I__7984 (
            .O(N__38288),
            .I(buf_adcdata_vac_5));
    Odrv4 I__7983 (
            .O(N__38285),
            .I(buf_adcdata_vac_5));
    Odrv4 I__7982 (
            .O(N__38282),
            .I(buf_adcdata_vac_5));
    InMux I__7981 (
            .O(N__38275),
            .I(N__38272));
    LocalMux I__7980 (
            .O(N__38272),
            .I(n19_adj_1598));
    InMux I__7979 (
            .O(N__38269),
            .I(N__38266));
    LocalMux I__7978 (
            .O(N__38266),
            .I(comm_buf_2_5));
    CascadeMux I__7977 (
            .O(N__38263),
            .I(N__38260));
    InMux I__7976 (
            .O(N__38260),
            .I(N__38256));
    InMux I__7975 (
            .O(N__38259),
            .I(N__38253));
    LocalMux I__7974 (
            .O(N__38256),
            .I(N__38250));
    LocalMux I__7973 (
            .O(N__38253),
            .I(N__38245));
    Span4Mux_h I__7972 (
            .O(N__38250),
            .I(N__38245));
    Odrv4 I__7971 (
            .O(N__38245),
            .I(comm_buf_6_5));
    InMux I__7970 (
            .O(N__38242),
            .I(N__38239));
    LocalMux I__7969 (
            .O(N__38239),
            .I(N__38236));
    Span4Mux_h I__7968 (
            .O(N__38236),
            .I(N__38233));
    Span4Mux_h I__7967 (
            .O(N__38233),
            .I(N__38230));
    Span4Mux_v I__7966 (
            .O(N__38230),
            .I(N__38227));
    Odrv4 I__7965 (
            .O(N__38227),
            .I(comm_buf_4_5));
    CascadeMux I__7964 (
            .O(N__38224),
            .I(n22123_cascade_));
    InMux I__7963 (
            .O(N__38221),
            .I(N__38218));
    LocalMux I__7962 (
            .O(N__38218),
            .I(N__38215));
    Span4Mux_h I__7961 (
            .O(N__38215),
            .I(N__38212));
    Odrv4 I__7960 (
            .O(N__38212),
            .I(n22126));
    InMux I__7959 (
            .O(N__38209),
            .I(N__38203));
    InMux I__7958 (
            .O(N__38208),
            .I(N__38203));
    LocalMux I__7957 (
            .O(N__38203),
            .I(N__38198));
    InMux I__7956 (
            .O(N__38202),
            .I(N__38193));
    InMux I__7955 (
            .O(N__38201),
            .I(N__38193));
    Span4Mux_h I__7954 (
            .O(N__38198),
            .I(N__38190));
    LocalMux I__7953 (
            .O(N__38193),
            .I(n20602));
    Odrv4 I__7952 (
            .O(N__38190),
            .I(n20602));
    IoInMux I__7951 (
            .O(N__38185),
            .I(N__38182));
    LocalMux I__7950 (
            .O(N__38182),
            .I(N__38179));
    IoSpan4Mux I__7949 (
            .O(N__38179),
            .I(N__38176));
    IoSpan4Mux I__7948 (
            .O(N__38176),
            .I(N__38172));
    InMux I__7947 (
            .O(N__38175),
            .I(N__38169));
    Span4Mux_s3_v I__7946 (
            .O(N__38172),
            .I(N__38166));
    LocalMux I__7945 (
            .O(N__38169),
            .I(N__38163));
    Span4Mux_v I__7944 (
            .O(N__38166),
            .I(N__38159));
    Span4Mux_h I__7943 (
            .O(N__38163),
            .I(N__38156));
    InMux I__7942 (
            .O(N__38162),
            .I(N__38153));
    Span4Mux_v I__7941 (
            .O(N__38159),
            .I(N__38148));
    Span4Mux_h I__7940 (
            .O(N__38156),
            .I(N__38148));
    LocalMux I__7939 (
            .O(N__38153),
            .I(SELIRNG0));
    Odrv4 I__7938 (
            .O(N__38148),
            .I(SELIRNG0));
    InMux I__7937 (
            .O(N__38143),
            .I(N__38140));
    LocalMux I__7936 (
            .O(N__38140),
            .I(N__38137));
    Odrv12 I__7935 (
            .O(N__38137),
            .I(n14_adj_1552));
    CascadeMux I__7934 (
            .O(N__38134),
            .I(n14_adj_1552_cascade_));
    InMux I__7933 (
            .O(N__38131),
            .I(N__38128));
    LocalMux I__7932 (
            .O(N__38128),
            .I(n16_adj_1570));
    CascadeMux I__7931 (
            .O(N__38125),
            .I(n12080_cascade_));
    InMux I__7930 (
            .O(N__38122),
            .I(N__38119));
    LocalMux I__7929 (
            .O(N__38119),
            .I(N__38116));
    Odrv4 I__7928 (
            .O(N__38116),
            .I(comm_buf_4_0));
    InMux I__7927 (
            .O(N__38113),
            .I(N__38110));
    LocalMux I__7926 (
            .O(N__38110),
            .I(N__38107));
    Odrv4 I__7925 (
            .O(N__38107),
            .I(n22132));
    CEMux I__7924 (
            .O(N__38104),
            .I(N__38101));
    LocalMux I__7923 (
            .O(N__38101),
            .I(N__38098));
    Odrv4 I__7922 (
            .O(N__38098),
            .I(n12206));
    CascadeMux I__7921 (
            .O(N__38095),
            .I(n12206_cascade_));
    SRMux I__7920 (
            .O(N__38092),
            .I(N__38089));
    LocalMux I__7919 (
            .O(N__38089),
            .I(N__38086));
    Odrv4 I__7918 (
            .O(N__38086),
            .I(n14770));
    InMux I__7917 (
            .O(N__38083),
            .I(N__38080));
    LocalMux I__7916 (
            .O(N__38080),
            .I(N__38077));
    Span4Mux_v I__7915 (
            .O(N__38077),
            .I(N__38073));
    CascadeMux I__7914 (
            .O(N__38076),
            .I(N__38070));
    Span4Mux_h I__7913 (
            .O(N__38073),
            .I(N__38067));
    InMux I__7912 (
            .O(N__38070),
            .I(N__38064));
    Span4Mux_v I__7911 (
            .O(N__38067),
            .I(N__38061));
    LocalMux I__7910 (
            .O(N__38064),
            .I(comm_buf_6_0));
    Odrv4 I__7909 (
            .O(N__38061),
            .I(comm_buf_6_0));
    CascadeMux I__7908 (
            .O(N__38056),
            .I(N__38053));
    InMux I__7907 (
            .O(N__38053),
            .I(N__38050));
    LocalMux I__7906 (
            .O(N__38050),
            .I(comm_buf_2_0));
    InMux I__7905 (
            .O(N__38047),
            .I(N__38044));
    LocalMux I__7904 (
            .O(N__38044),
            .I(n22129));
    InMux I__7903 (
            .O(N__38041),
            .I(N__38038));
    LocalMux I__7902 (
            .O(N__38038),
            .I(N__38035));
    Span12Mux_v I__7901 (
            .O(N__38035),
            .I(N__38032));
    Odrv12 I__7900 (
            .O(N__38032),
            .I(buf_data_iac_5));
    CascadeMux I__7899 (
            .O(N__38029),
            .I(n22_adj_1599_cascade_));
    CascadeMux I__7898 (
            .O(N__38026),
            .I(n30_adj_1600_cascade_));
    CascadeMux I__7897 (
            .O(N__38023),
            .I(N__38019));
    InMux I__7896 (
            .O(N__38022),
            .I(N__38013));
    InMux I__7895 (
            .O(N__38019),
            .I(N__38010));
    InMux I__7894 (
            .O(N__38018),
            .I(N__38007));
    InMux I__7893 (
            .O(N__38017),
            .I(N__38004));
    CascadeMux I__7892 (
            .O(N__38016),
            .I(N__38001));
    LocalMux I__7891 (
            .O(N__38013),
            .I(N__37996));
    LocalMux I__7890 (
            .O(N__38010),
            .I(N__37996));
    LocalMux I__7889 (
            .O(N__38007),
            .I(N__37991));
    LocalMux I__7888 (
            .O(N__38004),
            .I(N__37988));
    InMux I__7887 (
            .O(N__38001),
            .I(N__37985));
    Span4Mux_v I__7886 (
            .O(N__37996),
            .I(N__37982));
    InMux I__7885 (
            .O(N__37995),
            .I(N__37978));
    CascadeMux I__7884 (
            .O(N__37994),
            .I(N__37975));
    Span4Mux_v I__7883 (
            .O(N__37991),
            .I(N__37972));
    Span4Mux_v I__7882 (
            .O(N__37988),
            .I(N__37969));
    LocalMux I__7881 (
            .O(N__37985),
            .I(N__37966));
    Span4Mux_h I__7880 (
            .O(N__37982),
            .I(N__37963));
    InMux I__7879 (
            .O(N__37981),
            .I(N__37960));
    LocalMux I__7878 (
            .O(N__37978),
            .I(N__37957));
    InMux I__7877 (
            .O(N__37975),
            .I(N__37954));
    Span4Mux_v I__7876 (
            .O(N__37972),
            .I(N__37948));
    Span4Mux_v I__7875 (
            .O(N__37969),
            .I(N__37948));
    Span4Mux_h I__7874 (
            .O(N__37966),
            .I(N__37941));
    Span4Mux_h I__7873 (
            .O(N__37963),
            .I(N__37941));
    LocalMux I__7872 (
            .O(N__37960),
            .I(N__37941));
    Span4Mux_h I__7871 (
            .O(N__37957),
            .I(N__37938));
    LocalMux I__7870 (
            .O(N__37954),
            .I(N__37935));
    InMux I__7869 (
            .O(N__37953),
            .I(N__37932));
    Odrv4 I__7868 (
            .O(N__37948),
            .I(comm_rx_buf_5));
    Odrv4 I__7867 (
            .O(N__37941),
            .I(comm_rx_buf_5));
    Odrv4 I__7866 (
            .O(N__37938),
            .I(comm_rx_buf_5));
    Odrv4 I__7865 (
            .O(N__37935),
            .I(comm_rx_buf_5));
    LocalMux I__7864 (
            .O(N__37932),
            .I(comm_rx_buf_5));
    CEMux I__7863 (
            .O(N__37921),
            .I(N__37917));
    CEMux I__7862 (
            .O(N__37920),
            .I(N__37914));
    LocalMux I__7861 (
            .O(N__37917),
            .I(n12080));
    LocalMux I__7860 (
            .O(N__37914),
            .I(n12080));
    CascadeMux I__7859 (
            .O(N__37909),
            .I(n11839_cascade_));
    InMux I__7858 (
            .O(N__37906),
            .I(N__37902));
    InMux I__7857 (
            .O(N__37905),
            .I(N__37899));
    LocalMux I__7856 (
            .O(N__37902),
            .I(n9222));
    LocalMux I__7855 (
            .O(N__37899),
            .I(n9222));
    CascadeMux I__7854 (
            .O(N__37894),
            .I(n9222_cascade_));
    CascadeMux I__7853 (
            .O(N__37891),
            .I(n24_adj_1579_cascade_));
    CascadeMux I__7852 (
            .O(N__37888),
            .I(n21079_cascade_));
    InMux I__7851 (
            .O(N__37885),
            .I(N__37879));
    InMux I__7850 (
            .O(N__37884),
            .I(N__37879));
    LocalMux I__7849 (
            .O(N__37879),
            .I(N__37865));
    InMux I__7848 (
            .O(N__37878),
            .I(N__37860));
    InMux I__7847 (
            .O(N__37877),
            .I(N__37860));
    InMux I__7846 (
            .O(N__37876),
            .I(N__37851));
    InMux I__7845 (
            .O(N__37875),
            .I(N__37851));
    InMux I__7844 (
            .O(N__37874),
            .I(N__37851));
    InMux I__7843 (
            .O(N__37873),
            .I(N__37851));
    InMux I__7842 (
            .O(N__37872),
            .I(N__37848));
    InMux I__7841 (
            .O(N__37871),
            .I(N__37845));
    InMux I__7840 (
            .O(N__37870),
            .I(N__37841));
    InMux I__7839 (
            .O(N__37869),
            .I(N__37827));
    InMux I__7838 (
            .O(N__37868),
            .I(N__37827));
    Span4Mux_v I__7837 (
            .O(N__37865),
            .I(N__37824));
    LocalMux I__7836 (
            .O(N__37860),
            .I(N__37817));
    LocalMux I__7835 (
            .O(N__37851),
            .I(N__37817));
    LocalMux I__7834 (
            .O(N__37848),
            .I(N__37817));
    LocalMux I__7833 (
            .O(N__37845),
            .I(N__37814));
    InMux I__7832 (
            .O(N__37844),
            .I(N__37811));
    LocalMux I__7831 (
            .O(N__37841),
            .I(N__37808));
    InMux I__7830 (
            .O(N__37840),
            .I(N__37801));
    InMux I__7829 (
            .O(N__37839),
            .I(N__37801));
    InMux I__7828 (
            .O(N__37838),
            .I(N__37801));
    InMux I__7827 (
            .O(N__37837),
            .I(N__37788));
    InMux I__7826 (
            .O(N__37836),
            .I(N__37788));
    InMux I__7825 (
            .O(N__37835),
            .I(N__37788));
    InMux I__7824 (
            .O(N__37834),
            .I(N__37788));
    InMux I__7823 (
            .O(N__37833),
            .I(N__37788));
    InMux I__7822 (
            .O(N__37832),
            .I(N__37788));
    LocalMux I__7821 (
            .O(N__37827),
            .I(N__37776));
    Span4Mux_h I__7820 (
            .O(N__37824),
            .I(N__37771));
    Span4Mux_v I__7819 (
            .O(N__37817),
            .I(N__37771));
    Span12Mux_h I__7818 (
            .O(N__37814),
            .I(N__37766));
    LocalMux I__7817 (
            .O(N__37811),
            .I(N__37766));
    Span4Mux_v I__7816 (
            .O(N__37808),
            .I(N__37759));
    LocalMux I__7815 (
            .O(N__37801),
            .I(N__37759));
    LocalMux I__7814 (
            .O(N__37788),
            .I(N__37759));
    InMux I__7813 (
            .O(N__37787),
            .I(N__37752));
    InMux I__7812 (
            .O(N__37786),
            .I(N__37752));
    InMux I__7811 (
            .O(N__37785),
            .I(N__37752));
    InMux I__7810 (
            .O(N__37784),
            .I(N__37739));
    InMux I__7809 (
            .O(N__37783),
            .I(N__37739));
    InMux I__7808 (
            .O(N__37782),
            .I(N__37739));
    InMux I__7807 (
            .O(N__37781),
            .I(N__37739));
    InMux I__7806 (
            .O(N__37780),
            .I(N__37739));
    InMux I__7805 (
            .O(N__37779),
            .I(N__37739));
    Odrv4 I__7804 (
            .O(N__37776),
            .I(n12643));
    Odrv4 I__7803 (
            .O(N__37771),
            .I(n12643));
    Odrv12 I__7802 (
            .O(N__37766),
            .I(n12643));
    Odrv4 I__7801 (
            .O(N__37759),
            .I(n12643));
    LocalMux I__7800 (
            .O(N__37752),
            .I(n12643));
    LocalMux I__7799 (
            .O(N__37739),
            .I(n12643));
    InMux I__7798 (
            .O(N__37726),
            .I(N__37723));
    LocalMux I__7797 (
            .O(N__37723),
            .I(N__37720));
    Span4Mux_v I__7796 (
            .O(N__37720),
            .I(N__37715));
    InMux I__7795 (
            .O(N__37719),
            .I(N__37712));
    InMux I__7794 (
            .O(N__37718),
            .I(N__37709));
    Odrv4 I__7793 (
            .O(N__37715),
            .I(\comm_spi.n22644 ));
    LocalMux I__7792 (
            .O(N__37712),
            .I(\comm_spi.n22644 ));
    LocalMux I__7791 (
            .O(N__37709),
            .I(\comm_spi.n22644 ));
    SRMux I__7790 (
            .O(N__37702),
            .I(N__37699));
    LocalMux I__7789 (
            .O(N__37699),
            .I(N__37696));
    Odrv4 I__7788 (
            .O(N__37696),
            .I(\comm_spi.data_tx_7__N_778 ));
    InMux I__7787 (
            .O(N__37693),
            .I(N__37690));
    LocalMux I__7786 (
            .O(N__37690),
            .I(N__37686));
    InMux I__7785 (
            .O(N__37689),
            .I(N__37683));
    Odrv4 I__7784 (
            .O(N__37686),
            .I(\comm_spi.n14608 ));
    LocalMux I__7783 (
            .O(N__37683),
            .I(\comm_spi.n14608 ));
    SRMux I__7782 (
            .O(N__37678),
            .I(N__37675));
    LocalMux I__7781 (
            .O(N__37675),
            .I(N__37672));
    Span4Mux_h I__7780 (
            .O(N__37672),
            .I(N__37669));
    Odrv4 I__7779 (
            .O(N__37669),
            .I(\comm_spi.data_tx_7__N_781 ));
    InMux I__7778 (
            .O(N__37666),
            .I(N__37663));
    LocalMux I__7777 (
            .O(N__37663),
            .I(N__37659));
    InMux I__7776 (
            .O(N__37662),
            .I(N__37656));
    Span4Mux_v I__7775 (
            .O(N__37659),
            .I(N__37653));
    LocalMux I__7774 (
            .O(N__37656),
            .I(N__37650));
    Odrv4 I__7773 (
            .O(N__37653),
            .I(\comm_spi.n14607 ));
    Odrv4 I__7772 (
            .O(N__37650),
            .I(\comm_spi.n14607 ));
    SRMux I__7771 (
            .O(N__37645),
            .I(N__37642));
    LocalMux I__7770 (
            .O(N__37642),
            .I(N__37639));
    Sp12to4 I__7769 (
            .O(N__37639),
            .I(N__37636));
    Odrv12 I__7768 (
            .O(N__37636),
            .I(\comm_spi.data_tx_7__N_763 ));
    InMux I__7767 (
            .O(N__37633),
            .I(N__37630));
    LocalMux I__7766 (
            .O(N__37630),
            .I(N__37625));
    InMux I__7765 (
            .O(N__37629),
            .I(N__37620));
    InMux I__7764 (
            .O(N__37628),
            .I(N__37620));
    Span4Mux_h I__7763 (
            .O(N__37625),
            .I(N__37617));
    LocalMux I__7762 (
            .O(N__37620),
            .I(N__37614));
    Span4Mux_h I__7761 (
            .O(N__37617),
            .I(N__37609));
    Span4Mux_v I__7760 (
            .O(N__37614),
            .I(N__37609));
    Odrv4 I__7759 (
            .O(N__37609),
            .I(comm_tx_buf_3));
    InMux I__7758 (
            .O(N__37606),
            .I(N__37599));
    CascadeMux I__7757 (
            .O(N__37605),
            .I(N__37596));
    InMux I__7756 (
            .O(N__37604),
            .I(N__37590));
    InMux I__7755 (
            .O(N__37603),
            .I(N__37587));
    InMux I__7754 (
            .O(N__37602),
            .I(N__37584));
    LocalMux I__7753 (
            .O(N__37599),
            .I(N__37577));
    InMux I__7752 (
            .O(N__37596),
            .I(N__37574));
    InMux I__7751 (
            .O(N__37595),
            .I(N__37569));
    InMux I__7750 (
            .O(N__37594),
            .I(N__37569));
    InMux I__7749 (
            .O(N__37593),
            .I(N__37566));
    LocalMux I__7748 (
            .O(N__37590),
            .I(N__37559));
    LocalMux I__7747 (
            .O(N__37587),
            .I(N__37559));
    LocalMux I__7746 (
            .O(N__37584),
            .I(N__37559));
    InMux I__7745 (
            .O(N__37583),
            .I(N__37550));
    InMux I__7744 (
            .O(N__37582),
            .I(N__37550));
    InMux I__7743 (
            .O(N__37581),
            .I(N__37550));
    InMux I__7742 (
            .O(N__37580),
            .I(N__37550));
    Span4Mux_h I__7741 (
            .O(N__37577),
            .I(N__37547));
    LocalMux I__7740 (
            .O(N__37574),
            .I(N__37540));
    LocalMux I__7739 (
            .O(N__37569),
            .I(N__37540));
    LocalMux I__7738 (
            .O(N__37566),
            .I(N__37540));
    Span4Mux_v I__7737 (
            .O(N__37559),
            .I(N__37537));
    LocalMux I__7736 (
            .O(N__37550),
            .I(eis_state_0));
    Odrv4 I__7735 (
            .O(N__37547),
            .I(eis_state_0));
    Odrv12 I__7734 (
            .O(N__37540),
            .I(eis_state_0));
    Odrv4 I__7733 (
            .O(N__37537),
            .I(eis_state_0));
    InMux I__7732 (
            .O(N__37528),
            .I(N__37525));
    LocalMux I__7731 (
            .O(N__37525),
            .I(N__37522));
    Span4Mux_v I__7730 (
            .O(N__37522),
            .I(N__37519));
    Odrv4 I__7729 (
            .O(N__37519),
            .I(n21067));
    InMux I__7728 (
            .O(N__37516),
            .I(N__37512));
    InMux I__7727 (
            .O(N__37515),
            .I(N__37509));
    LocalMux I__7726 (
            .O(N__37512),
            .I(N__37506));
    LocalMux I__7725 (
            .O(N__37509),
            .I(n10508));
    Odrv12 I__7724 (
            .O(N__37506),
            .I(n10508));
    InMux I__7723 (
            .O(N__37501),
            .I(\ADC_VDC.genclk.n19439 ));
    CascadeMux I__7722 (
            .O(N__37498),
            .I(N__37494));
    InMux I__7721 (
            .O(N__37497),
            .I(N__37491));
    InMux I__7720 (
            .O(N__37494),
            .I(N__37488));
    LocalMux I__7719 (
            .O(N__37491),
            .I(\ADC_VDC.genclk.t0on_15 ));
    LocalMux I__7718 (
            .O(N__37488),
            .I(\ADC_VDC.genclk.t0on_15 ));
    CEMux I__7717 (
            .O(N__37483),
            .I(N__37479));
    CEMux I__7716 (
            .O(N__37482),
            .I(N__37476));
    LocalMux I__7715 (
            .O(N__37479),
            .I(N__37473));
    LocalMux I__7714 (
            .O(N__37476),
            .I(N__37470));
    Span4Mux_v I__7713 (
            .O(N__37473),
            .I(N__37467));
    Span4Mux_v I__7712 (
            .O(N__37470),
            .I(N__37464));
    Span4Mux_h I__7711 (
            .O(N__37467),
            .I(N__37459));
    Span4Mux_h I__7710 (
            .O(N__37464),
            .I(N__37459));
    Odrv4 I__7709 (
            .O(N__37459),
            .I(\ADC_VDC.genclk.div_state_1__N_1266 ));
    SRMux I__7708 (
            .O(N__37456),
            .I(N__37453));
    LocalMux I__7707 (
            .O(N__37453),
            .I(N__37449));
    SRMux I__7706 (
            .O(N__37452),
            .I(N__37446));
    Span4Mux_v I__7705 (
            .O(N__37449),
            .I(N__37439));
    LocalMux I__7704 (
            .O(N__37446),
            .I(N__37439));
    SRMux I__7703 (
            .O(N__37445),
            .I(N__37436));
    SRMux I__7702 (
            .O(N__37444),
            .I(N__37433));
    Odrv4 I__7701 (
            .O(N__37439),
            .I(\ADC_VDC.genclk.n14695 ));
    LocalMux I__7700 (
            .O(N__37436),
            .I(\ADC_VDC.genclk.n14695 ));
    LocalMux I__7699 (
            .O(N__37433),
            .I(\ADC_VDC.genclk.n14695 ));
    InMux I__7698 (
            .O(N__37426),
            .I(N__37421));
    InMux I__7697 (
            .O(N__37425),
            .I(N__37418));
    InMux I__7696 (
            .O(N__37424),
            .I(N__37415));
    LocalMux I__7695 (
            .O(N__37421),
            .I(N__37412));
    LocalMux I__7694 (
            .O(N__37418),
            .I(N__37407));
    LocalMux I__7693 (
            .O(N__37415),
            .I(N__37407));
    Span4Mux_v I__7692 (
            .O(N__37412),
            .I(N__37404));
    Span4Mux_h I__7691 (
            .O(N__37407),
            .I(N__37401));
    Odrv4 I__7690 (
            .O(N__37404),
            .I(\comm_spi.n14585 ));
    Odrv4 I__7689 (
            .O(N__37401),
            .I(\comm_spi.n14585 ));
    CascadeMux I__7688 (
            .O(N__37396),
            .I(N__37392));
    InMux I__7687 (
            .O(N__37395),
            .I(N__37388));
    InMux I__7686 (
            .O(N__37392),
            .I(N__37383));
    InMux I__7685 (
            .O(N__37391),
            .I(N__37383));
    LocalMux I__7684 (
            .O(N__37388),
            .I(comm_tx_buf_7));
    LocalMux I__7683 (
            .O(N__37383),
            .I(comm_tx_buf_7));
    InMux I__7682 (
            .O(N__37378),
            .I(N__37369));
    InMux I__7681 (
            .O(N__37377),
            .I(N__37369));
    InMux I__7680 (
            .O(N__37376),
            .I(N__37369));
    LocalMux I__7679 (
            .O(N__37369),
            .I(N__37366));
    Odrv4 I__7678 (
            .O(N__37366),
            .I(comm_tx_buf_2));
    SRMux I__7677 (
            .O(N__37363),
            .I(N__37360));
    LocalMux I__7676 (
            .O(N__37360),
            .I(\comm_spi.imosi_N_744 ));
    InMux I__7675 (
            .O(N__37357),
            .I(N__37350));
    InMux I__7674 (
            .O(N__37356),
            .I(N__37350));
    InMux I__7673 (
            .O(N__37355),
            .I(N__37347));
    LocalMux I__7672 (
            .O(N__37350),
            .I(N__37343));
    LocalMux I__7671 (
            .O(N__37347),
            .I(N__37339));
    InMux I__7670 (
            .O(N__37346),
            .I(N__37336));
    Span4Mux_v I__7669 (
            .O(N__37343),
            .I(N__37333));
    InMux I__7668 (
            .O(N__37342),
            .I(N__37330));
    Span4Mux_h I__7667 (
            .O(N__37339),
            .I(N__37325));
    LocalMux I__7666 (
            .O(N__37336),
            .I(N__37325));
    Sp12to4 I__7665 (
            .O(N__37333),
            .I(N__37322));
    LocalMux I__7664 (
            .O(N__37330),
            .I(N__37317));
    Sp12to4 I__7663 (
            .O(N__37325),
            .I(N__37317));
    Span12Mux_h I__7662 (
            .O(N__37322),
            .I(N__37314));
    Span12Mux_v I__7661 (
            .O(N__37317),
            .I(N__37311));
    Span12Mux_v I__7660 (
            .O(N__37314),
            .I(N__37308));
    Span12Mux_h I__7659 (
            .O(N__37311),
            .I(N__37305));
    Odrv12 I__7658 (
            .O(N__37308),
            .I(ICE_SPI_MOSI));
    Odrv12 I__7657 (
            .O(N__37305),
            .I(ICE_SPI_MOSI));
    SRMux I__7656 (
            .O(N__37300),
            .I(N__37297));
    LocalMux I__7655 (
            .O(N__37297),
            .I(N__37294));
    Span4Mux_h I__7654 (
            .O(N__37294),
            .I(N__37291));
    Odrv4 I__7653 (
            .O(N__37291),
            .I(\comm_spi.imosi_N_745 ));
    CascadeMux I__7652 (
            .O(N__37288),
            .I(N__37284));
    InMux I__7651 (
            .O(N__37287),
            .I(N__37281));
    InMux I__7650 (
            .O(N__37284),
            .I(N__37278));
    LocalMux I__7649 (
            .O(N__37281),
            .I(\ADC_VDC.genclk.t0on_7 ));
    LocalMux I__7648 (
            .O(N__37278),
            .I(\ADC_VDC.genclk.t0on_7 ));
    InMux I__7647 (
            .O(N__37273),
            .I(\ADC_VDC.genclk.n19431 ));
    InMux I__7646 (
            .O(N__37270),
            .I(N__37266));
    InMux I__7645 (
            .O(N__37269),
            .I(N__37263));
    LocalMux I__7644 (
            .O(N__37266),
            .I(\ADC_VDC.genclk.t0on_8 ));
    LocalMux I__7643 (
            .O(N__37263),
            .I(\ADC_VDC.genclk.t0on_8 ));
    InMux I__7642 (
            .O(N__37258),
            .I(bfn_15_4_0_));
    CascadeMux I__7641 (
            .O(N__37255),
            .I(N__37252));
    InMux I__7640 (
            .O(N__37252),
            .I(N__37248));
    InMux I__7639 (
            .O(N__37251),
            .I(N__37245));
    LocalMux I__7638 (
            .O(N__37248),
            .I(\ADC_VDC.genclk.t0on_9 ));
    LocalMux I__7637 (
            .O(N__37245),
            .I(\ADC_VDC.genclk.t0on_9 ));
    InMux I__7636 (
            .O(N__37240),
            .I(\ADC_VDC.genclk.n19433 ));
    InMux I__7635 (
            .O(N__37237),
            .I(N__37233));
    InMux I__7634 (
            .O(N__37236),
            .I(N__37230));
    LocalMux I__7633 (
            .O(N__37233),
            .I(\ADC_VDC.genclk.t0on_10 ));
    LocalMux I__7632 (
            .O(N__37230),
            .I(\ADC_VDC.genclk.t0on_10 ));
    InMux I__7631 (
            .O(N__37225),
            .I(\ADC_VDC.genclk.n19434 ));
    CascadeMux I__7630 (
            .O(N__37222),
            .I(N__37219));
    InMux I__7629 (
            .O(N__37219),
            .I(N__37215));
    InMux I__7628 (
            .O(N__37218),
            .I(N__37212));
    LocalMux I__7627 (
            .O(N__37215),
            .I(\ADC_VDC.genclk.t0on_11 ));
    LocalMux I__7626 (
            .O(N__37212),
            .I(\ADC_VDC.genclk.t0on_11 ));
    InMux I__7625 (
            .O(N__37207),
            .I(\ADC_VDC.genclk.n19435 ));
    InMux I__7624 (
            .O(N__37204),
            .I(N__37200));
    InMux I__7623 (
            .O(N__37203),
            .I(N__37197));
    LocalMux I__7622 (
            .O(N__37200),
            .I(\ADC_VDC.genclk.t0on_12 ));
    LocalMux I__7621 (
            .O(N__37197),
            .I(\ADC_VDC.genclk.t0on_12 ));
    InMux I__7620 (
            .O(N__37192),
            .I(\ADC_VDC.genclk.n19436 ));
    CascadeMux I__7619 (
            .O(N__37189),
            .I(N__37186));
    InMux I__7618 (
            .O(N__37186),
            .I(N__37182));
    InMux I__7617 (
            .O(N__37185),
            .I(N__37179));
    LocalMux I__7616 (
            .O(N__37182),
            .I(\ADC_VDC.genclk.t0on_13 ));
    LocalMux I__7615 (
            .O(N__37179),
            .I(\ADC_VDC.genclk.t0on_13 ));
    InMux I__7614 (
            .O(N__37174),
            .I(\ADC_VDC.genclk.n19437 ));
    InMux I__7613 (
            .O(N__37171),
            .I(N__37167));
    InMux I__7612 (
            .O(N__37170),
            .I(N__37164));
    LocalMux I__7611 (
            .O(N__37167),
            .I(\ADC_VDC.genclk.t0on_14 ));
    LocalMux I__7610 (
            .O(N__37164),
            .I(\ADC_VDC.genclk.t0on_14 ));
    InMux I__7609 (
            .O(N__37159),
            .I(\ADC_VDC.genclk.n19438 ));
    CascadeMux I__7608 (
            .O(N__37156),
            .I(N__37153));
    InMux I__7607 (
            .O(N__37153),
            .I(N__37150));
    LocalMux I__7606 (
            .O(N__37150),
            .I(\SIG_DDS.tmp_buf_4 ));
    CascadeMux I__7605 (
            .O(N__37147),
            .I(N__37144));
    InMux I__7604 (
            .O(N__37144),
            .I(N__37141));
    LocalMux I__7603 (
            .O(N__37141),
            .I(\SIG_DDS.tmp_buf_5 ));
    InMux I__7602 (
            .O(N__37138),
            .I(N__37135));
    LocalMux I__7601 (
            .O(N__37135),
            .I(N__37132));
    Span4Mux_h I__7600 (
            .O(N__37132),
            .I(N__37129));
    Odrv4 I__7599 (
            .O(N__37129),
            .I(\SIG_DDS.tmp_buf_6 ));
    InMux I__7598 (
            .O(N__37126),
            .I(N__37122));
    InMux I__7597 (
            .O(N__37125),
            .I(N__37119));
    LocalMux I__7596 (
            .O(N__37122),
            .I(\ADC_VDC.genclk.t0on_0 ));
    LocalMux I__7595 (
            .O(N__37119),
            .I(\ADC_VDC.genclk.t0on_0 ));
    InMux I__7594 (
            .O(N__37114),
            .I(bfn_15_3_0_));
    InMux I__7593 (
            .O(N__37111),
            .I(N__37107));
    InMux I__7592 (
            .O(N__37110),
            .I(N__37104));
    LocalMux I__7591 (
            .O(N__37107),
            .I(\ADC_VDC.genclk.t0on_1 ));
    LocalMux I__7590 (
            .O(N__37104),
            .I(\ADC_VDC.genclk.t0on_1 ));
    InMux I__7589 (
            .O(N__37099),
            .I(\ADC_VDC.genclk.n19425 ));
    CascadeMux I__7588 (
            .O(N__37096),
            .I(N__37093));
    InMux I__7587 (
            .O(N__37093),
            .I(N__37089));
    InMux I__7586 (
            .O(N__37092),
            .I(N__37086));
    LocalMux I__7585 (
            .O(N__37089),
            .I(\ADC_VDC.genclk.t0on_2 ));
    LocalMux I__7584 (
            .O(N__37086),
            .I(\ADC_VDC.genclk.t0on_2 ));
    InMux I__7583 (
            .O(N__37081),
            .I(\ADC_VDC.genclk.n19426 ));
    InMux I__7582 (
            .O(N__37078),
            .I(N__37074));
    InMux I__7581 (
            .O(N__37077),
            .I(N__37071));
    LocalMux I__7580 (
            .O(N__37074),
            .I(\ADC_VDC.genclk.t0on_3 ));
    LocalMux I__7579 (
            .O(N__37071),
            .I(\ADC_VDC.genclk.t0on_3 ));
    InMux I__7578 (
            .O(N__37066),
            .I(\ADC_VDC.genclk.n19427 ));
    CascadeMux I__7577 (
            .O(N__37063),
            .I(N__37059));
    CascadeMux I__7576 (
            .O(N__37062),
            .I(N__37056));
    InMux I__7575 (
            .O(N__37059),
            .I(N__37053));
    InMux I__7574 (
            .O(N__37056),
            .I(N__37050));
    LocalMux I__7573 (
            .O(N__37053),
            .I(N__37047));
    LocalMux I__7572 (
            .O(N__37050),
            .I(\ADC_VDC.genclk.t0on_4 ));
    Odrv4 I__7571 (
            .O(N__37047),
            .I(\ADC_VDC.genclk.t0on_4 ));
    InMux I__7570 (
            .O(N__37042),
            .I(\ADC_VDC.genclk.n19428 ));
    CascadeMux I__7569 (
            .O(N__37039),
            .I(N__37035));
    InMux I__7568 (
            .O(N__37038),
            .I(N__37032));
    InMux I__7567 (
            .O(N__37035),
            .I(N__37029));
    LocalMux I__7566 (
            .O(N__37032),
            .I(\ADC_VDC.genclk.t0on_5 ));
    LocalMux I__7565 (
            .O(N__37029),
            .I(\ADC_VDC.genclk.t0on_5 ));
    InMux I__7564 (
            .O(N__37024),
            .I(\ADC_VDC.genclk.n19429 ));
    CascadeMux I__7563 (
            .O(N__37021),
            .I(N__37018));
    InMux I__7562 (
            .O(N__37018),
            .I(N__37014));
    InMux I__7561 (
            .O(N__37017),
            .I(N__37011));
    LocalMux I__7560 (
            .O(N__37014),
            .I(\ADC_VDC.genclk.t0on_6 ));
    LocalMux I__7559 (
            .O(N__37011),
            .I(\ADC_VDC.genclk.t0on_6 ));
    InMux I__7558 (
            .O(N__37006),
            .I(\ADC_VDC.genclk.n19430 ));
    CascadeMux I__7557 (
            .O(N__37003),
            .I(N__37000));
    InMux I__7556 (
            .O(N__37000),
            .I(N__36997));
    LocalMux I__7555 (
            .O(N__36997),
            .I(N__36994));
    Odrv4 I__7554 (
            .O(N__36994),
            .I(n20949));
    InMux I__7553 (
            .O(N__36991),
            .I(N__36988));
    LocalMux I__7552 (
            .O(N__36988),
            .I(n26_adj_1623));
    CascadeMux I__7551 (
            .O(N__36985),
            .I(n21949_cascade_));
    InMux I__7550 (
            .O(N__36982),
            .I(N__36979));
    LocalMux I__7549 (
            .O(N__36979),
            .I(N__36974));
    InMux I__7548 (
            .O(N__36978),
            .I(N__36969));
    InMux I__7547 (
            .O(N__36977),
            .I(N__36969));
    Odrv4 I__7546 (
            .O(N__36974),
            .I(acadc_skipCount_7));
    LocalMux I__7545 (
            .O(N__36969),
            .I(acadc_skipCount_7));
    InMux I__7544 (
            .O(N__36964),
            .I(N__36961));
    LocalMux I__7543 (
            .O(N__36961),
            .I(N__36958));
    Span4Mux_h I__7542 (
            .O(N__36958),
            .I(N__36955));
    Odrv4 I__7541 (
            .O(N__36955),
            .I(n21964));
    CascadeMux I__7540 (
            .O(N__36952),
            .I(n21952_cascade_));
    InMux I__7539 (
            .O(N__36949),
            .I(N__36944));
    InMux I__7538 (
            .O(N__36948),
            .I(N__36941));
    InMux I__7537 (
            .O(N__36947),
            .I(N__36938));
    LocalMux I__7536 (
            .O(N__36944),
            .I(N__36935));
    LocalMux I__7535 (
            .O(N__36941),
            .I(N__36932));
    LocalMux I__7534 (
            .O(N__36938),
            .I(acadc_skipCount_4));
    Odrv4 I__7533 (
            .O(N__36935),
            .I(acadc_skipCount_4));
    Odrv4 I__7532 (
            .O(N__36932),
            .I(acadc_skipCount_4));
    InMux I__7531 (
            .O(N__36925),
            .I(N__36922));
    LocalMux I__7530 (
            .O(N__36922),
            .I(N__36917));
    CascadeMux I__7529 (
            .O(N__36921),
            .I(N__36914));
    InMux I__7528 (
            .O(N__36920),
            .I(N__36911));
    Span12Mux_h I__7527 (
            .O(N__36917),
            .I(N__36908));
    InMux I__7526 (
            .O(N__36914),
            .I(N__36905));
    LocalMux I__7525 (
            .O(N__36911),
            .I(acadc_skipCount_9));
    Odrv12 I__7524 (
            .O(N__36908),
            .I(acadc_skipCount_9));
    LocalMux I__7523 (
            .O(N__36905),
            .I(acadc_skipCount_9));
    InMux I__7522 (
            .O(N__36898),
            .I(N__36891));
    CascadeMux I__7521 (
            .O(N__36897),
            .I(N__36888));
    InMux I__7520 (
            .O(N__36896),
            .I(N__36885));
    InMux I__7519 (
            .O(N__36895),
            .I(N__36882));
    InMux I__7518 (
            .O(N__36894),
            .I(N__36877));
    LocalMux I__7517 (
            .O(N__36891),
            .I(N__36874));
    InMux I__7516 (
            .O(N__36888),
            .I(N__36871));
    LocalMux I__7515 (
            .O(N__36885),
            .I(N__36868));
    LocalMux I__7514 (
            .O(N__36882),
            .I(N__36865));
    InMux I__7513 (
            .O(N__36881),
            .I(N__36862));
    CascadeMux I__7512 (
            .O(N__36880),
            .I(N__36859));
    LocalMux I__7511 (
            .O(N__36877),
            .I(N__36855));
    Span4Mux_v I__7510 (
            .O(N__36874),
            .I(N__36850));
    LocalMux I__7509 (
            .O(N__36871),
            .I(N__36850));
    Span4Mux_h I__7508 (
            .O(N__36868),
            .I(N__36843));
    Span4Mux_v I__7507 (
            .O(N__36865),
            .I(N__36843));
    LocalMux I__7506 (
            .O(N__36862),
            .I(N__36843));
    InMux I__7505 (
            .O(N__36859),
            .I(N__36840));
    CascadeMux I__7504 (
            .O(N__36858),
            .I(N__36837));
    Span12Mux_v I__7503 (
            .O(N__36855),
            .I(N__36834));
    Span4Mux_h I__7502 (
            .O(N__36850),
            .I(N__36831));
    Span4Mux_h I__7501 (
            .O(N__36843),
            .I(N__36826));
    LocalMux I__7500 (
            .O(N__36840),
            .I(N__36826));
    InMux I__7499 (
            .O(N__36837),
            .I(N__36823));
    Odrv12 I__7498 (
            .O(N__36834),
            .I(comm_rx_buf_7));
    Odrv4 I__7497 (
            .O(N__36831),
            .I(comm_rx_buf_7));
    Odrv4 I__7496 (
            .O(N__36826),
            .I(comm_rx_buf_7));
    LocalMux I__7495 (
            .O(N__36823),
            .I(comm_rx_buf_7));
    InMux I__7494 (
            .O(N__36814),
            .I(N__36811));
    LocalMux I__7493 (
            .O(N__36811),
            .I(n30_adj_1624));
    SRMux I__7492 (
            .O(N__36808),
            .I(N__36804));
    SRMux I__7491 (
            .O(N__36807),
            .I(N__36800));
    LocalMux I__7490 (
            .O(N__36804),
            .I(N__36797));
    SRMux I__7489 (
            .O(N__36803),
            .I(N__36792));
    LocalMux I__7488 (
            .O(N__36800),
            .I(N__36787));
    Span4Mux_h I__7487 (
            .O(N__36797),
            .I(N__36784));
    SRMux I__7486 (
            .O(N__36796),
            .I(N__36781));
    SRMux I__7485 (
            .O(N__36795),
            .I(N__36777));
    LocalMux I__7484 (
            .O(N__36792),
            .I(N__36774));
    SRMux I__7483 (
            .O(N__36791),
            .I(N__36771));
    SRMux I__7482 (
            .O(N__36790),
            .I(N__36768));
    Span4Mux_v I__7481 (
            .O(N__36787),
            .I(N__36761));
    Span4Mux_h I__7480 (
            .O(N__36784),
            .I(N__36761));
    LocalMux I__7479 (
            .O(N__36781),
            .I(N__36761));
    SRMux I__7478 (
            .O(N__36780),
            .I(N__36758));
    LocalMux I__7477 (
            .O(N__36777),
            .I(N__36755));
    Span4Mux_v I__7476 (
            .O(N__36774),
            .I(N__36752));
    LocalMux I__7475 (
            .O(N__36771),
            .I(N__36749));
    LocalMux I__7474 (
            .O(N__36768),
            .I(N__36742));
    Span4Mux_v I__7473 (
            .O(N__36761),
            .I(N__36742));
    LocalMux I__7472 (
            .O(N__36758),
            .I(N__36742));
    Span4Mux_h I__7471 (
            .O(N__36755),
            .I(N__36737));
    Span4Mux_h I__7470 (
            .O(N__36752),
            .I(N__36737));
    Span4Mux_h I__7469 (
            .O(N__36749),
            .I(N__36734));
    Sp12to4 I__7468 (
            .O(N__36742),
            .I(N__36731));
    Odrv4 I__7467 (
            .O(N__36737),
            .I(n14742));
    Odrv4 I__7466 (
            .O(N__36734),
            .I(n14742));
    Odrv12 I__7465 (
            .O(N__36731),
            .I(n14742));
    CascadeMux I__7464 (
            .O(N__36724),
            .I(N__36721));
    InMux I__7463 (
            .O(N__36721),
            .I(N__36718));
    LocalMux I__7462 (
            .O(N__36718),
            .I(N__36714));
    InMux I__7461 (
            .O(N__36717),
            .I(N__36710));
    Span4Mux_v I__7460 (
            .O(N__36714),
            .I(N__36707));
    InMux I__7459 (
            .O(N__36713),
            .I(N__36704));
    LocalMux I__7458 (
            .O(N__36710),
            .I(buf_dds0_3));
    Odrv4 I__7457 (
            .O(N__36707),
            .I(buf_dds0_3));
    LocalMux I__7456 (
            .O(N__36704),
            .I(buf_dds0_3));
    InMux I__7455 (
            .O(N__36697),
            .I(N__36694));
    LocalMux I__7454 (
            .O(N__36694),
            .I(\SIG_DDS.tmp_buf_2 ));
    CascadeMux I__7453 (
            .O(N__36691),
            .I(N__36688));
    InMux I__7452 (
            .O(N__36688),
            .I(N__36685));
    LocalMux I__7451 (
            .O(N__36685),
            .I(\SIG_DDS.tmp_buf_3 ));
    InMux I__7450 (
            .O(N__36682),
            .I(N__36679));
    LocalMux I__7449 (
            .O(N__36679),
            .I(N__36675));
    InMux I__7448 (
            .O(N__36678),
            .I(N__36672));
    Span4Mux_v I__7447 (
            .O(N__36675),
            .I(N__36669));
    LocalMux I__7446 (
            .O(N__36672),
            .I(data_idxvec_7));
    Odrv4 I__7445 (
            .O(N__36669),
            .I(data_idxvec_7));
    InMux I__7444 (
            .O(N__36664),
            .I(N__36661));
    LocalMux I__7443 (
            .O(N__36661),
            .I(N__36658));
    Span4Mux_v I__7442 (
            .O(N__36658),
            .I(N__36654));
    InMux I__7441 (
            .O(N__36657),
            .I(N__36650));
    Span4Mux_h I__7440 (
            .O(N__36654),
            .I(N__36647));
    InMux I__7439 (
            .O(N__36653),
            .I(N__36644));
    LocalMux I__7438 (
            .O(N__36650),
            .I(acadc_skipCount_14));
    Odrv4 I__7437 (
            .O(N__36647),
            .I(acadc_skipCount_14));
    LocalMux I__7436 (
            .O(N__36644),
            .I(acadc_skipCount_14));
    InMux I__7435 (
            .O(N__36637),
            .I(N__36631));
    InMux I__7434 (
            .O(N__36636),
            .I(N__36631));
    LocalMux I__7433 (
            .O(N__36631),
            .I(n8_adj_1545));
    InMux I__7432 (
            .O(N__36628),
            .I(N__36624));
    InMux I__7431 (
            .O(N__36627),
            .I(N__36621));
    LocalMux I__7430 (
            .O(N__36624),
            .I(N__36618));
    LocalMux I__7429 (
            .O(N__36621),
            .I(acadc_skipcnt_9));
    Odrv4 I__7428 (
            .O(N__36618),
            .I(acadc_skipcnt_9));
    InMux I__7427 (
            .O(N__36613),
            .I(N__36609));
    InMux I__7426 (
            .O(N__36612),
            .I(N__36606));
    LocalMux I__7425 (
            .O(N__36609),
            .I(N__36603));
    LocalMux I__7424 (
            .O(N__36606),
            .I(acadc_skipcnt_15));
    Odrv4 I__7423 (
            .O(N__36603),
            .I(acadc_skipcnt_15));
    InMux I__7422 (
            .O(N__36598),
            .I(N__36595));
    LocalMux I__7421 (
            .O(N__36595),
            .I(N__36592));
    Span4Mux_h I__7420 (
            .O(N__36592),
            .I(N__36589));
    Span4Mux_v I__7419 (
            .O(N__36589),
            .I(N__36584));
    InMux I__7418 (
            .O(N__36588),
            .I(N__36579));
    InMux I__7417 (
            .O(N__36587),
            .I(N__36579));
    Odrv4 I__7416 (
            .O(N__36584),
            .I(acadc_skipCount_15));
    LocalMux I__7415 (
            .O(N__36579),
            .I(acadc_skipCount_15));
    InMux I__7414 (
            .O(N__36574),
            .I(N__36571));
    LocalMux I__7413 (
            .O(N__36571),
            .I(n24));
    CascadeMux I__7412 (
            .O(N__36568),
            .I(N__36565));
    InMux I__7411 (
            .O(N__36565),
            .I(N__36560));
    InMux I__7410 (
            .O(N__36564),
            .I(N__36557));
    InMux I__7409 (
            .O(N__36563),
            .I(N__36554));
    LocalMux I__7408 (
            .O(N__36560),
            .I(N__36551));
    LocalMux I__7407 (
            .O(N__36557),
            .I(N__36548));
    LocalMux I__7406 (
            .O(N__36554),
            .I(N__36545));
    Odrv4 I__7405 (
            .O(N__36551),
            .I(acadc_skipCount_1));
    Odrv4 I__7404 (
            .O(N__36548),
            .I(acadc_skipCount_1));
    Odrv12 I__7403 (
            .O(N__36545),
            .I(acadc_skipCount_1));
    InMux I__7402 (
            .O(N__36538),
            .I(N__36535));
    LocalMux I__7401 (
            .O(N__36535),
            .I(N__36532));
    Span4Mux_h I__7400 (
            .O(N__36532),
            .I(N__36529));
    Odrv4 I__7399 (
            .O(N__36529),
            .I(n9_adj_1407));
    CascadeMux I__7398 (
            .O(N__36526),
            .I(N__36523));
    CascadeBuf I__7397 (
            .O(N__36523),
            .I(N__36520));
    CascadeMux I__7396 (
            .O(N__36520),
            .I(N__36517));
    CascadeBuf I__7395 (
            .O(N__36517),
            .I(N__36514));
    CascadeMux I__7394 (
            .O(N__36514),
            .I(N__36511));
    CascadeBuf I__7393 (
            .O(N__36511),
            .I(N__36508));
    CascadeMux I__7392 (
            .O(N__36508),
            .I(N__36505));
    CascadeBuf I__7391 (
            .O(N__36505),
            .I(N__36502));
    CascadeMux I__7390 (
            .O(N__36502),
            .I(N__36499));
    CascadeBuf I__7389 (
            .O(N__36499),
            .I(N__36496));
    CascadeMux I__7388 (
            .O(N__36496),
            .I(N__36493));
    CascadeBuf I__7387 (
            .O(N__36493),
            .I(N__36490));
    CascadeMux I__7386 (
            .O(N__36490),
            .I(N__36487));
    CascadeBuf I__7385 (
            .O(N__36487),
            .I(N__36484));
    CascadeMux I__7384 (
            .O(N__36484),
            .I(N__36481));
    CascadeBuf I__7383 (
            .O(N__36481),
            .I(N__36478));
    CascadeMux I__7382 (
            .O(N__36478),
            .I(N__36474));
    CascadeMux I__7381 (
            .O(N__36477),
            .I(N__36471));
    CascadeBuf I__7380 (
            .O(N__36474),
            .I(N__36468));
    CascadeBuf I__7379 (
            .O(N__36471),
            .I(N__36465));
    CascadeMux I__7378 (
            .O(N__36468),
            .I(N__36462));
    CascadeMux I__7377 (
            .O(N__36465),
            .I(N__36459));
    InMux I__7376 (
            .O(N__36462),
            .I(N__36456));
    InMux I__7375 (
            .O(N__36459),
            .I(N__36453));
    LocalMux I__7374 (
            .O(N__36456),
            .I(N__36450));
    LocalMux I__7373 (
            .O(N__36453),
            .I(N__36447));
    Span4Mux_v I__7372 (
            .O(N__36450),
            .I(N__36444));
    Span4Mux_v I__7371 (
            .O(N__36447),
            .I(N__36441));
    Span4Mux_h I__7370 (
            .O(N__36444),
            .I(N__36438));
    Span4Mux_h I__7369 (
            .O(N__36441),
            .I(N__36433));
    Span4Mux_h I__7368 (
            .O(N__36438),
            .I(N__36433));
    Odrv4 I__7367 (
            .O(N__36433),
            .I(data_index_9_N_212_2));
    InMux I__7366 (
            .O(N__36430),
            .I(N__36427));
    LocalMux I__7365 (
            .O(N__36427),
            .I(N__36423));
    InMux I__7364 (
            .O(N__36426),
            .I(N__36420));
    Span4Mux_v I__7363 (
            .O(N__36423),
            .I(N__36417));
    LocalMux I__7362 (
            .O(N__36420),
            .I(acadc_skipcnt_14));
    Odrv4 I__7361 (
            .O(N__36417),
            .I(acadc_skipcnt_14));
    InMux I__7360 (
            .O(N__36412),
            .I(N__36408));
    InMux I__7359 (
            .O(N__36411),
            .I(N__36405));
    LocalMux I__7358 (
            .O(N__36408),
            .I(N__36402));
    LocalMux I__7357 (
            .O(N__36405),
            .I(acadc_skipcnt_11));
    Odrv4 I__7356 (
            .O(N__36402),
            .I(acadc_skipcnt_11));
    InMux I__7355 (
            .O(N__36397),
            .I(N__36391));
    CascadeMux I__7354 (
            .O(N__36396),
            .I(N__36388));
    InMux I__7353 (
            .O(N__36395),
            .I(N__36385));
    InMux I__7352 (
            .O(N__36394),
            .I(N__36382));
    LocalMux I__7351 (
            .O(N__36391),
            .I(N__36379));
    InMux I__7350 (
            .O(N__36388),
            .I(N__36375));
    LocalMux I__7349 (
            .O(N__36385),
            .I(N__36370));
    LocalMux I__7348 (
            .O(N__36382),
            .I(N__36370));
    Span4Mux_v I__7347 (
            .O(N__36379),
            .I(N__36367));
    InMux I__7346 (
            .O(N__36378),
            .I(N__36364));
    LocalMux I__7345 (
            .O(N__36375),
            .I(N__36361));
    Span12Mux_v I__7344 (
            .O(N__36370),
            .I(N__36358));
    Span4Mux_h I__7343 (
            .O(N__36367),
            .I(N__36353));
    LocalMux I__7342 (
            .O(N__36364),
            .I(N__36353));
    Odrv12 I__7341 (
            .O(N__36361),
            .I(comm_buf_1_3));
    Odrv12 I__7340 (
            .O(N__36358),
            .I(comm_buf_1_3));
    Odrv4 I__7339 (
            .O(N__36353),
            .I(comm_buf_1_3));
    InMux I__7338 (
            .O(N__36346),
            .I(N__36340));
    InMux I__7337 (
            .O(N__36345),
            .I(N__36340));
    LocalMux I__7336 (
            .O(N__36340),
            .I(N__36337));
    Odrv12 I__7335 (
            .O(N__36337),
            .I(n8_adj_1543));
    InMux I__7334 (
            .O(N__36334),
            .I(N__36330));
    InMux I__7333 (
            .O(N__36333),
            .I(N__36327));
    LocalMux I__7332 (
            .O(N__36330),
            .I(N__36324));
    LocalMux I__7331 (
            .O(N__36327),
            .I(acadc_skipcnt_2));
    Odrv4 I__7330 (
            .O(N__36324),
            .I(acadc_skipcnt_2));
    InMux I__7329 (
            .O(N__36319),
            .I(N__36315));
    InMux I__7328 (
            .O(N__36318),
            .I(N__36312));
    LocalMux I__7327 (
            .O(N__36315),
            .I(N__36309));
    LocalMux I__7326 (
            .O(N__36312),
            .I(acadc_skipcnt_7));
    Odrv4 I__7325 (
            .O(N__36309),
            .I(acadc_skipcnt_7));
    InMux I__7324 (
            .O(N__36304),
            .I(N__36299));
    CascadeMux I__7323 (
            .O(N__36303),
            .I(N__36296));
    InMux I__7322 (
            .O(N__36302),
            .I(N__36293));
    LocalMux I__7321 (
            .O(N__36299),
            .I(N__36290));
    InMux I__7320 (
            .O(N__36296),
            .I(N__36287));
    LocalMux I__7319 (
            .O(N__36293),
            .I(acadc_skipCount_2));
    Odrv4 I__7318 (
            .O(N__36290),
            .I(acadc_skipCount_2));
    LocalMux I__7317 (
            .O(N__36287),
            .I(acadc_skipCount_2));
    InMux I__7316 (
            .O(N__36280),
            .I(N__36277));
    LocalMux I__7315 (
            .O(N__36277),
            .I(n23_adj_1586));
    CascadeMux I__7314 (
            .O(N__36274),
            .I(n22_cascade_));
    InMux I__7313 (
            .O(N__36271),
            .I(N__36268));
    LocalMux I__7312 (
            .O(N__36268),
            .I(N__36265));
    Odrv4 I__7311 (
            .O(N__36265),
            .I(n30_adj_1571));
    CascadeMux I__7310 (
            .O(N__36262),
            .I(n30_adj_1478_cascade_));
    InMux I__7309 (
            .O(N__36259),
            .I(N__36256));
    LocalMux I__7308 (
            .O(N__36256),
            .I(N__36249));
    InMux I__7307 (
            .O(N__36255),
            .I(N__36246));
    InMux I__7306 (
            .O(N__36254),
            .I(N__36243));
    InMux I__7305 (
            .O(N__36253),
            .I(N__36238));
    InMux I__7304 (
            .O(N__36252),
            .I(N__36234));
    Span4Mux_v I__7303 (
            .O(N__36249),
            .I(N__36228));
    LocalMux I__7302 (
            .O(N__36246),
            .I(N__36228));
    LocalMux I__7301 (
            .O(N__36243),
            .I(N__36225));
    InMux I__7300 (
            .O(N__36242),
            .I(N__36222));
    InMux I__7299 (
            .O(N__36241),
            .I(N__36219));
    LocalMux I__7298 (
            .O(N__36238),
            .I(N__36216));
    InMux I__7297 (
            .O(N__36237),
            .I(N__36213));
    LocalMux I__7296 (
            .O(N__36234),
            .I(N__36210));
    InMux I__7295 (
            .O(N__36233),
            .I(N__36207));
    Span4Mux_v I__7294 (
            .O(N__36228),
            .I(N__36204));
    Span4Mux_v I__7293 (
            .O(N__36225),
            .I(N__36199));
    LocalMux I__7292 (
            .O(N__36222),
            .I(N__36199));
    LocalMux I__7291 (
            .O(N__36219),
            .I(N__36188));
    Span4Mux_v I__7290 (
            .O(N__36216),
            .I(N__36188));
    LocalMux I__7289 (
            .O(N__36213),
            .I(N__36188));
    Span4Mux_h I__7288 (
            .O(N__36210),
            .I(N__36188));
    LocalMux I__7287 (
            .O(N__36207),
            .I(N__36188));
    Span4Mux_h I__7286 (
            .O(N__36204),
            .I(N__36185));
    Span4Mux_v I__7285 (
            .O(N__36199),
            .I(N__36182));
    Span4Mux_v I__7284 (
            .O(N__36188),
            .I(N__36179));
    Span4Mux_v I__7283 (
            .O(N__36185),
            .I(N__36176));
    Span4Mux_v I__7282 (
            .O(N__36182),
            .I(N__36171));
    Span4Mux_v I__7281 (
            .O(N__36179),
            .I(N__36171));
    Odrv4 I__7280 (
            .O(N__36176),
            .I(comm_rx_buf_0));
    Odrv4 I__7279 (
            .O(N__36171),
            .I(comm_rx_buf_0));
    CascadeMux I__7278 (
            .O(N__36166),
            .I(N__36161));
    InMux I__7277 (
            .O(N__36165),
            .I(N__36154));
    InMux I__7276 (
            .O(N__36164),
            .I(N__36154));
    InMux I__7275 (
            .O(N__36161),
            .I(N__36154));
    LocalMux I__7274 (
            .O(N__36154),
            .I(cmd_rdadctmp_13_adj_1430));
    InMux I__7273 (
            .O(N__36151),
            .I(N__36148));
    LocalMux I__7272 (
            .O(N__36148),
            .I(N__36145));
    Span4Mux_v I__7271 (
            .O(N__36145),
            .I(N__36140));
    InMux I__7270 (
            .O(N__36144),
            .I(N__36137));
    InMux I__7269 (
            .O(N__36143),
            .I(N__36134));
    Span4Mux_h I__7268 (
            .O(N__36140),
            .I(N__36131));
    LocalMux I__7267 (
            .O(N__36137),
            .I(buf_dds1_4));
    LocalMux I__7266 (
            .O(N__36134),
            .I(buf_dds1_4));
    Odrv4 I__7265 (
            .O(N__36131),
            .I(buf_dds1_4));
    InMux I__7264 (
            .O(N__36124),
            .I(N__36121));
    LocalMux I__7263 (
            .O(N__36121),
            .I(N__36118));
    Odrv4 I__7262 (
            .O(N__36118),
            .I(n16));
    InMux I__7261 (
            .O(N__36115),
            .I(N__36112));
    LocalMux I__7260 (
            .O(N__36112),
            .I(N__36109));
    Span4Mux_v I__7259 (
            .O(N__36109),
            .I(N__36105));
    InMux I__7258 (
            .O(N__36108),
            .I(N__36101));
    Span4Mux_h I__7257 (
            .O(N__36105),
            .I(N__36098));
    InMux I__7256 (
            .O(N__36104),
            .I(N__36095));
    LocalMux I__7255 (
            .O(N__36101),
            .I(buf_dds1_6));
    Odrv4 I__7254 (
            .O(N__36098),
            .I(buf_dds1_6));
    LocalMux I__7253 (
            .O(N__36095),
            .I(buf_dds1_6));
    InMux I__7252 (
            .O(N__36088),
            .I(N__36085));
    LocalMux I__7251 (
            .O(N__36085),
            .I(N__36082));
    Odrv4 I__7250 (
            .O(N__36082),
            .I(n16_adj_1488));
    CascadeMux I__7249 (
            .O(N__36079),
            .I(N__36076));
    InMux I__7248 (
            .O(N__36076),
            .I(N__36073));
    LocalMux I__7247 (
            .O(N__36073),
            .I(N__36070));
    Odrv4 I__7246 (
            .O(N__36070),
            .I(n20824));
    InMux I__7245 (
            .O(N__36067),
            .I(N__36064));
    LocalMux I__7244 (
            .O(N__36064),
            .I(N__36061));
    Span4Mux_v I__7243 (
            .O(N__36061),
            .I(N__36058));
    Span4Mux_h I__7242 (
            .O(N__36058),
            .I(N__36055));
    Span4Mux_h I__7241 (
            .O(N__36055),
            .I(N__36052));
    Odrv4 I__7240 (
            .O(N__36052),
            .I(n20836));
    CascadeMux I__7239 (
            .O(N__36049),
            .I(n22069_cascade_));
    InMux I__7238 (
            .O(N__36046),
            .I(N__36043));
    LocalMux I__7237 (
            .O(N__36043),
            .I(n20837));
    InMux I__7236 (
            .O(N__36040),
            .I(N__36036));
    InMux I__7235 (
            .O(N__36039),
            .I(N__36033));
    LocalMux I__7234 (
            .O(N__36036),
            .I(N__36030));
    LocalMux I__7233 (
            .O(N__36033),
            .I(data_idxvec_1));
    Odrv4 I__7232 (
            .O(N__36030),
            .I(data_idxvec_1));
    CascadeMux I__7231 (
            .O(N__36025),
            .I(n26_adj_1509_cascade_));
    InMux I__7230 (
            .O(N__36022),
            .I(N__36019));
    LocalMux I__7229 (
            .O(N__36019),
            .I(N__36016));
    Span4Mux_h I__7228 (
            .O(N__36016),
            .I(N__36013));
    Span4Mux_v I__7227 (
            .O(N__36013),
            .I(N__36010));
    Span4Mux_h I__7226 (
            .O(N__36010),
            .I(N__36007));
    Span4Mux_h I__7225 (
            .O(N__36007),
            .I(N__36004));
    Odrv4 I__7224 (
            .O(N__36004),
            .I(buf_data_iac_9));
    InMux I__7223 (
            .O(N__36001),
            .I(N__35998));
    LocalMux I__7222 (
            .O(N__35998),
            .I(n20825));
    InMux I__7221 (
            .O(N__35995),
            .I(N__35992));
    LocalMux I__7220 (
            .O(N__35992),
            .I(N__35988));
    InMux I__7219 (
            .O(N__35991),
            .I(N__35985));
    Span4Mux_v I__7218 (
            .O(N__35988),
            .I(N__35982));
    LocalMux I__7217 (
            .O(N__35985),
            .I(N__35979));
    Span4Mux_h I__7216 (
            .O(N__35982),
            .I(N__35972));
    Span4Mux_h I__7215 (
            .O(N__35979),
            .I(N__35972));
    CascadeMux I__7214 (
            .O(N__35978),
            .I(N__35968));
    InMux I__7213 (
            .O(N__35977),
            .I(N__35964));
    Span4Mux_h I__7212 (
            .O(N__35972),
            .I(N__35961));
    InMux I__7211 (
            .O(N__35971),
            .I(N__35958));
    InMux I__7210 (
            .O(N__35968),
            .I(N__35955));
    InMux I__7209 (
            .O(N__35967),
            .I(N__35952));
    LocalMux I__7208 (
            .O(N__35964),
            .I(N__35948));
    Span4Mux_h I__7207 (
            .O(N__35961),
            .I(N__35943));
    LocalMux I__7206 (
            .O(N__35958),
            .I(N__35943));
    LocalMux I__7205 (
            .O(N__35955),
            .I(N__35938));
    LocalMux I__7204 (
            .O(N__35952),
            .I(N__35938));
    InMux I__7203 (
            .O(N__35951),
            .I(N__35935));
    Span4Mux_h I__7202 (
            .O(N__35948),
            .I(N__35930));
    Span4Mux_v I__7201 (
            .O(N__35943),
            .I(N__35927));
    Span4Mux_h I__7200 (
            .O(N__35938),
            .I(N__35922));
    LocalMux I__7199 (
            .O(N__35935),
            .I(N__35922));
    InMux I__7198 (
            .O(N__35934),
            .I(N__35919));
    InMux I__7197 (
            .O(N__35933),
            .I(N__35916));
    Odrv4 I__7196 (
            .O(N__35930),
            .I(comm_rx_buf_1));
    Odrv4 I__7195 (
            .O(N__35927),
            .I(comm_rx_buf_1));
    Odrv4 I__7194 (
            .O(N__35922),
            .I(comm_rx_buf_1));
    LocalMux I__7193 (
            .O(N__35919),
            .I(comm_rx_buf_1));
    LocalMux I__7192 (
            .O(N__35916),
            .I(comm_rx_buf_1));
    InMux I__7191 (
            .O(N__35905),
            .I(N__35902));
    LocalMux I__7190 (
            .O(N__35902),
            .I(n22072));
    InMux I__7189 (
            .O(N__35899),
            .I(N__35896));
    LocalMux I__7188 (
            .O(N__35896),
            .I(N__35892));
    InMux I__7187 (
            .O(N__35895),
            .I(N__35889));
    Span4Mux_h I__7186 (
            .O(N__35892),
            .I(N__35886));
    LocalMux I__7185 (
            .O(N__35889),
            .I(data_idxvec_0));
    Odrv4 I__7184 (
            .O(N__35886),
            .I(data_idxvec_0));
    InMux I__7183 (
            .O(N__35881),
            .I(N__35878));
    LocalMux I__7182 (
            .O(N__35878),
            .I(N__35875));
    Span4Mux_h I__7181 (
            .O(N__35875),
            .I(N__35872));
    Span4Mux_h I__7180 (
            .O(N__35872),
            .I(N__35869));
    Span4Mux_h I__7179 (
            .O(N__35869),
            .I(N__35866));
    Odrv4 I__7178 (
            .O(N__35866),
            .I(n21001));
    CascadeMux I__7177 (
            .O(N__35863),
            .I(n26_cascade_));
    InMux I__7176 (
            .O(N__35860),
            .I(N__35857));
    LocalMux I__7175 (
            .O(N__35857),
            .I(N__35852));
    InMux I__7174 (
            .O(N__35856),
            .I(N__35849));
    InMux I__7173 (
            .O(N__35855),
            .I(N__35846));
    Span4Mux_v I__7172 (
            .O(N__35852),
            .I(N__35843));
    LocalMux I__7171 (
            .O(N__35849),
            .I(N__35838));
    LocalMux I__7170 (
            .O(N__35846),
            .I(N__35838));
    Odrv4 I__7169 (
            .O(N__35843),
            .I(acadc_skipCount_0));
    Odrv4 I__7168 (
            .O(N__35838),
            .I(acadc_skipCount_0));
    CascadeMux I__7167 (
            .O(N__35833),
            .I(n22021_cascade_));
    InMux I__7166 (
            .O(N__35830),
            .I(N__35827));
    LocalMux I__7165 (
            .O(N__35827),
            .I(n22024));
    InMux I__7164 (
            .O(N__35824),
            .I(N__35821));
    LocalMux I__7163 (
            .O(N__35821),
            .I(N__35818));
    Span12Mux_v I__7162 (
            .O(N__35818),
            .I(N__35815));
    Odrv12 I__7161 (
            .O(N__35815),
            .I(n21976));
    InMux I__7160 (
            .O(N__35812),
            .I(N__35807));
    CascadeMux I__7159 (
            .O(N__35811),
            .I(N__35803));
    InMux I__7158 (
            .O(N__35810),
            .I(N__35799));
    LocalMux I__7157 (
            .O(N__35807),
            .I(N__35795));
    InMux I__7156 (
            .O(N__35806),
            .I(N__35792));
    InMux I__7155 (
            .O(N__35803),
            .I(N__35789));
    InMux I__7154 (
            .O(N__35802),
            .I(N__35786));
    LocalMux I__7153 (
            .O(N__35799),
            .I(N__35783));
    InMux I__7152 (
            .O(N__35798),
            .I(N__35780));
    Span4Mux_h I__7151 (
            .O(N__35795),
            .I(N__35776));
    LocalMux I__7150 (
            .O(N__35792),
            .I(N__35773));
    LocalMux I__7149 (
            .O(N__35789),
            .I(N__35770));
    LocalMux I__7148 (
            .O(N__35786),
            .I(N__35767));
    Span4Mux_v I__7147 (
            .O(N__35783),
            .I(N__35762));
    LocalMux I__7146 (
            .O(N__35780),
            .I(N__35762));
    InMux I__7145 (
            .O(N__35779),
            .I(N__35759));
    Span4Mux_v I__7144 (
            .O(N__35776),
            .I(N__35754));
    Span4Mux_v I__7143 (
            .O(N__35773),
            .I(N__35751));
    Span4Mux_h I__7142 (
            .O(N__35770),
            .I(N__35748));
    Span4Mux_h I__7141 (
            .O(N__35767),
            .I(N__35745));
    Span4Mux_h I__7140 (
            .O(N__35762),
            .I(N__35742));
    LocalMux I__7139 (
            .O(N__35759),
            .I(N__35739));
    InMux I__7138 (
            .O(N__35758),
            .I(N__35736));
    InMux I__7137 (
            .O(N__35757),
            .I(N__35733));
    Odrv4 I__7136 (
            .O(N__35754),
            .I(comm_rx_buf_6));
    Odrv4 I__7135 (
            .O(N__35751),
            .I(comm_rx_buf_6));
    Odrv4 I__7134 (
            .O(N__35748),
            .I(comm_rx_buf_6));
    Odrv4 I__7133 (
            .O(N__35745),
            .I(comm_rx_buf_6));
    Odrv4 I__7132 (
            .O(N__35742),
            .I(comm_rx_buf_6));
    Odrv12 I__7131 (
            .O(N__35739),
            .I(comm_rx_buf_6));
    LocalMux I__7130 (
            .O(N__35736),
            .I(comm_rx_buf_6));
    LocalMux I__7129 (
            .O(N__35733),
            .I(comm_rx_buf_6));
    InMux I__7128 (
            .O(N__35716),
            .I(N__35713));
    LocalMux I__7127 (
            .O(N__35713),
            .I(N__35710));
    Span4Mux_h I__7126 (
            .O(N__35710),
            .I(N__35707));
    Span4Mux_h I__7125 (
            .O(N__35707),
            .I(N__35704));
    Odrv4 I__7124 (
            .O(N__35704),
            .I(buf_data_vac_6));
    InMux I__7123 (
            .O(N__35701),
            .I(N__35698));
    LocalMux I__7122 (
            .O(N__35698),
            .I(N__35695));
    Span4Mux_v I__7121 (
            .O(N__35695),
            .I(N__35692));
    Odrv4 I__7120 (
            .O(N__35692),
            .I(comm_buf_5_6));
    InMux I__7119 (
            .O(N__35689),
            .I(N__35686));
    LocalMux I__7118 (
            .O(N__35686),
            .I(N__35683));
    Span4Mux_h I__7117 (
            .O(N__35683),
            .I(N__35680));
    Span4Mux_h I__7116 (
            .O(N__35680),
            .I(N__35677));
    Odrv4 I__7115 (
            .O(N__35677),
            .I(buf_data_vac_5));
    InMux I__7114 (
            .O(N__35674),
            .I(N__35671));
    LocalMux I__7113 (
            .O(N__35671),
            .I(comm_buf_5_5));
    InMux I__7112 (
            .O(N__35668),
            .I(N__35665));
    LocalMux I__7111 (
            .O(N__35665),
            .I(N__35658));
    InMux I__7110 (
            .O(N__35664),
            .I(N__35655));
    CascadeMux I__7109 (
            .O(N__35663),
            .I(N__35652));
    InMux I__7108 (
            .O(N__35662),
            .I(N__35649));
    InMux I__7107 (
            .O(N__35661),
            .I(N__35646));
    Span4Mux_h I__7106 (
            .O(N__35658),
            .I(N__35641));
    LocalMux I__7105 (
            .O(N__35655),
            .I(N__35641));
    InMux I__7104 (
            .O(N__35652),
            .I(N__35637));
    LocalMux I__7103 (
            .O(N__35649),
            .I(N__35633));
    LocalMux I__7102 (
            .O(N__35646),
            .I(N__35628));
    Span4Mux_h I__7101 (
            .O(N__35641),
            .I(N__35628));
    InMux I__7100 (
            .O(N__35640),
            .I(N__35625));
    LocalMux I__7099 (
            .O(N__35637),
            .I(N__35622));
    InMux I__7098 (
            .O(N__35636),
            .I(N__35619));
    Span4Mux_h I__7097 (
            .O(N__35633),
            .I(N__35614));
    Sp12to4 I__7096 (
            .O(N__35628),
            .I(N__35611));
    LocalMux I__7095 (
            .O(N__35625),
            .I(N__35608));
    Span4Mux_h I__7094 (
            .O(N__35622),
            .I(N__35603));
    LocalMux I__7093 (
            .O(N__35619),
            .I(N__35603));
    InMux I__7092 (
            .O(N__35618),
            .I(N__35600));
    InMux I__7091 (
            .O(N__35617),
            .I(N__35597));
    Odrv4 I__7090 (
            .O(N__35614),
            .I(comm_rx_buf_4));
    Odrv12 I__7089 (
            .O(N__35611),
            .I(comm_rx_buf_4));
    Odrv12 I__7088 (
            .O(N__35608),
            .I(comm_rx_buf_4));
    Odrv4 I__7087 (
            .O(N__35603),
            .I(comm_rx_buf_4));
    LocalMux I__7086 (
            .O(N__35600),
            .I(comm_rx_buf_4));
    LocalMux I__7085 (
            .O(N__35597),
            .I(comm_rx_buf_4));
    InMux I__7084 (
            .O(N__35584),
            .I(N__35581));
    LocalMux I__7083 (
            .O(N__35581),
            .I(N__35578));
    Span4Mux_h I__7082 (
            .O(N__35578),
            .I(N__35575));
    Span4Mux_h I__7081 (
            .O(N__35575),
            .I(N__35572));
    Odrv4 I__7080 (
            .O(N__35572),
            .I(buf_data_vac_4));
    InMux I__7079 (
            .O(N__35569),
            .I(N__35564));
    CascadeMux I__7078 (
            .O(N__35568),
            .I(N__35560));
    CascadeMux I__7077 (
            .O(N__35567),
            .I(N__35555));
    LocalMux I__7076 (
            .O(N__35564),
            .I(N__35552));
    InMux I__7075 (
            .O(N__35563),
            .I(N__35549));
    InMux I__7074 (
            .O(N__35560),
            .I(N__35546));
    InMux I__7073 (
            .O(N__35559),
            .I(N__35543));
    InMux I__7072 (
            .O(N__35558),
            .I(N__35540));
    InMux I__7071 (
            .O(N__35555),
            .I(N__35537));
    Span4Mux_v I__7070 (
            .O(N__35552),
            .I(N__35534));
    LocalMux I__7069 (
            .O(N__35549),
            .I(N__35531));
    LocalMux I__7068 (
            .O(N__35546),
            .I(N__35525));
    LocalMux I__7067 (
            .O(N__35543),
            .I(N__35525));
    LocalMux I__7066 (
            .O(N__35540),
            .I(N__35522));
    LocalMux I__7065 (
            .O(N__35537),
            .I(N__35519));
    Span4Mux_v I__7064 (
            .O(N__35534),
            .I(N__35514));
    Span4Mux_h I__7063 (
            .O(N__35531),
            .I(N__35514));
    InMux I__7062 (
            .O(N__35530),
            .I(N__35511));
    Span4Mux_v I__7061 (
            .O(N__35525),
            .I(N__35502));
    Span4Mux_h I__7060 (
            .O(N__35522),
            .I(N__35502));
    Span4Mux_v I__7059 (
            .O(N__35519),
            .I(N__35502));
    Span4Mux_h I__7058 (
            .O(N__35514),
            .I(N__35497));
    LocalMux I__7057 (
            .O(N__35511),
            .I(N__35497));
    InMux I__7056 (
            .O(N__35510),
            .I(N__35494));
    InMux I__7055 (
            .O(N__35509),
            .I(N__35491));
    Odrv4 I__7054 (
            .O(N__35502),
            .I(comm_rx_buf_3));
    Odrv4 I__7053 (
            .O(N__35497),
            .I(comm_rx_buf_3));
    LocalMux I__7052 (
            .O(N__35494),
            .I(comm_rx_buf_3));
    LocalMux I__7051 (
            .O(N__35491),
            .I(comm_rx_buf_3));
    InMux I__7050 (
            .O(N__35482),
            .I(N__35479));
    LocalMux I__7049 (
            .O(N__35479),
            .I(N__35476));
    Span4Mux_h I__7048 (
            .O(N__35476),
            .I(N__35473));
    Span4Mux_v I__7047 (
            .O(N__35473),
            .I(N__35470));
    Span4Mux_h I__7046 (
            .O(N__35470),
            .I(N__35467));
    Span4Mux_h I__7045 (
            .O(N__35467),
            .I(N__35464));
    Odrv4 I__7044 (
            .O(N__35464),
            .I(buf_data_vac_3));
    InMux I__7043 (
            .O(N__35461),
            .I(N__35458));
    LocalMux I__7042 (
            .O(N__35458),
            .I(N__35455));
    Odrv4 I__7041 (
            .O(N__35455),
            .I(comm_buf_5_3));
    InMux I__7040 (
            .O(N__35452),
            .I(N__35445));
    InMux I__7039 (
            .O(N__35451),
            .I(N__35442));
    InMux I__7038 (
            .O(N__35450),
            .I(N__35438));
    InMux I__7037 (
            .O(N__35449),
            .I(N__35433));
    InMux I__7036 (
            .O(N__35448),
            .I(N__35433));
    LocalMux I__7035 (
            .O(N__35445),
            .I(N__35428));
    LocalMux I__7034 (
            .O(N__35442),
            .I(N__35428));
    InMux I__7033 (
            .O(N__35441),
            .I(N__35425));
    LocalMux I__7032 (
            .O(N__35438),
            .I(N__35422));
    LocalMux I__7031 (
            .O(N__35433),
            .I(N__35417));
    Span4Mux_v I__7030 (
            .O(N__35428),
            .I(N__35414));
    LocalMux I__7029 (
            .O(N__35425),
            .I(N__35411));
    Span4Mux_v I__7028 (
            .O(N__35422),
            .I(N__35408));
    InMux I__7027 (
            .O(N__35421),
            .I(N__35405));
    CascadeMux I__7026 (
            .O(N__35420),
            .I(N__35402));
    Span4Mux_v I__7025 (
            .O(N__35417),
            .I(N__35398));
    Sp12to4 I__7024 (
            .O(N__35414),
            .I(N__35395));
    Span4Mux_h I__7023 (
            .O(N__35411),
            .I(N__35392));
    Span4Mux_h I__7022 (
            .O(N__35408),
            .I(N__35387));
    LocalMux I__7021 (
            .O(N__35405),
            .I(N__35387));
    InMux I__7020 (
            .O(N__35402),
            .I(N__35384));
    InMux I__7019 (
            .O(N__35401),
            .I(N__35381));
    Odrv4 I__7018 (
            .O(N__35398),
            .I(comm_rx_buf_2));
    Odrv12 I__7017 (
            .O(N__35395),
            .I(comm_rx_buf_2));
    Odrv4 I__7016 (
            .O(N__35392),
            .I(comm_rx_buf_2));
    Odrv4 I__7015 (
            .O(N__35387),
            .I(comm_rx_buf_2));
    LocalMux I__7014 (
            .O(N__35384),
            .I(comm_rx_buf_2));
    LocalMux I__7013 (
            .O(N__35381),
            .I(comm_rx_buf_2));
    InMux I__7012 (
            .O(N__35368),
            .I(N__35365));
    LocalMux I__7011 (
            .O(N__35365),
            .I(N__35362));
    Span12Mux_v I__7010 (
            .O(N__35362),
            .I(N__35359));
    Odrv12 I__7009 (
            .O(N__35359),
            .I(buf_data_vac_2));
    InMux I__7008 (
            .O(N__35356),
            .I(N__35353));
    LocalMux I__7007 (
            .O(N__35353),
            .I(N__35350));
    Odrv12 I__7006 (
            .O(N__35350),
            .I(comm_buf_5_2));
    InMux I__7005 (
            .O(N__35347),
            .I(N__35344));
    LocalMux I__7004 (
            .O(N__35344),
            .I(N__35341));
    Span12Mux_v I__7003 (
            .O(N__35341),
            .I(N__35338));
    Odrv12 I__7002 (
            .O(N__35338),
            .I(buf_data_vac_1));
    InMux I__7001 (
            .O(N__35335),
            .I(N__35332));
    LocalMux I__7000 (
            .O(N__35332),
            .I(N__35329));
    Span4Mux_v I__6999 (
            .O(N__35329),
            .I(N__35326));
    Span4Mux_h I__6998 (
            .O(N__35326),
            .I(N__35322));
    CascadeMux I__6997 (
            .O(N__35325),
            .I(N__35319));
    Span4Mux_h I__6996 (
            .O(N__35322),
            .I(N__35316));
    InMux I__6995 (
            .O(N__35319),
            .I(N__35313));
    Odrv4 I__6994 (
            .O(N__35316),
            .I(buf_readRTD_1));
    LocalMux I__6993 (
            .O(N__35313),
            .I(buf_readRTD_1));
    InMux I__6992 (
            .O(N__35308),
            .I(N__35305));
    LocalMux I__6991 (
            .O(N__35305),
            .I(N__35302));
    Span4Mux_v I__6990 (
            .O(N__35302),
            .I(N__35298));
    CascadeMux I__6989 (
            .O(N__35301),
            .I(N__35295));
    Span4Mux_h I__6988 (
            .O(N__35298),
            .I(N__35292));
    InMux I__6987 (
            .O(N__35295),
            .I(N__35289));
    Odrv4 I__6986 (
            .O(N__35292),
            .I(buf_adcdata_vdc_9));
    LocalMux I__6985 (
            .O(N__35289),
            .I(buf_adcdata_vdc_9));
    InMux I__6984 (
            .O(N__35284),
            .I(N__35280));
    InMux I__6983 (
            .O(N__35283),
            .I(N__35277));
    LocalMux I__6982 (
            .O(N__35280),
            .I(N__35273));
    LocalMux I__6981 (
            .O(N__35277),
            .I(N__35270));
    CascadeMux I__6980 (
            .O(N__35276),
            .I(N__35267));
    Span4Mux_v I__6979 (
            .O(N__35273),
            .I(N__35264));
    Span4Mux_v I__6978 (
            .O(N__35270),
            .I(N__35261));
    InMux I__6977 (
            .O(N__35267),
            .I(N__35258));
    Span4Mux_h I__6976 (
            .O(N__35264),
            .I(N__35255));
    Span4Mux_h I__6975 (
            .O(N__35261),
            .I(N__35252));
    LocalMux I__6974 (
            .O(N__35258),
            .I(buf_adcdata_vac_9));
    Odrv4 I__6973 (
            .O(N__35255),
            .I(buf_adcdata_vac_9));
    Odrv4 I__6972 (
            .O(N__35252),
            .I(buf_adcdata_vac_9));
    InMux I__6971 (
            .O(N__35245),
            .I(N__35242));
    LocalMux I__6970 (
            .O(N__35242),
            .I(n19_adj_1508));
    InMux I__6969 (
            .O(N__35239),
            .I(N__35236));
    LocalMux I__6968 (
            .O(N__35236),
            .I(N__35233));
    Odrv12 I__6967 (
            .O(N__35233),
            .I(n30_adj_1475));
    InMux I__6966 (
            .O(N__35230),
            .I(N__35227));
    LocalMux I__6965 (
            .O(N__35227),
            .I(N__35224));
    Odrv12 I__6964 (
            .O(N__35224),
            .I(comm_buf_2_7));
    InMux I__6963 (
            .O(N__35221),
            .I(N__35218));
    LocalMux I__6962 (
            .O(N__35218),
            .I(N__35215));
    Odrv4 I__6961 (
            .O(N__35215),
            .I(n30_adj_1595));
    InMux I__6960 (
            .O(N__35212),
            .I(N__35209));
    LocalMux I__6959 (
            .O(N__35209),
            .I(N__35206));
    Odrv4 I__6958 (
            .O(N__35206),
            .I(comm_buf_2_6));
    InMux I__6957 (
            .O(N__35203),
            .I(N__35200));
    LocalMux I__6956 (
            .O(N__35200),
            .I(N__35197));
    Span12Mux_h I__6955 (
            .O(N__35197),
            .I(N__35194));
    Odrv12 I__6954 (
            .O(N__35194),
            .I(n30_adj_1612));
    InMux I__6953 (
            .O(N__35191),
            .I(N__35188));
    LocalMux I__6952 (
            .O(N__35188),
            .I(comm_buf_2_3));
    InMux I__6951 (
            .O(N__35185),
            .I(N__35182));
    LocalMux I__6950 (
            .O(N__35182),
            .I(N__35179));
    Span12Mux_h I__6949 (
            .O(N__35179),
            .I(N__35176));
    Odrv12 I__6948 (
            .O(N__35176),
            .I(n30_adj_1615));
    InMux I__6947 (
            .O(N__35173),
            .I(N__35170));
    LocalMux I__6946 (
            .O(N__35170),
            .I(N__35167));
    Odrv4 I__6945 (
            .O(N__35167),
            .I(comm_buf_2_2));
    InMux I__6944 (
            .O(N__35164),
            .I(N__35161));
    LocalMux I__6943 (
            .O(N__35161),
            .I(N__35158));
    Span4Mux_v I__6942 (
            .O(N__35158),
            .I(N__35155));
    Span4Mux_h I__6941 (
            .O(N__35155),
            .I(N__35152));
    Odrv4 I__6940 (
            .O(N__35152),
            .I(n30_adj_1619));
    InMux I__6939 (
            .O(N__35149),
            .I(N__35146));
    LocalMux I__6938 (
            .O(N__35146),
            .I(comm_buf_2_1));
    InMux I__6937 (
            .O(N__35143),
            .I(N__35140));
    LocalMux I__6936 (
            .O(N__35140),
            .I(N__35137));
    Span12Mux_v I__6935 (
            .O(N__35137),
            .I(N__35134));
    Odrv12 I__6934 (
            .O(N__35134),
            .I(buf_data_vac_0));
    InMux I__6933 (
            .O(N__35131),
            .I(N__35128));
    LocalMux I__6932 (
            .O(N__35128),
            .I(N__35125));
    Span4Mux_h I__6931 (
            .O(N__35125),
            .I(N__35122));
    Odrv4 I__6930 (
            .O(N__35122),
            .I(comm_buf_5_0));
    InMux I__6929 (
            .O(N__35119),
            .I(N__35116));
    LocalMux I__6928 (
            .O(N__35116),
            .I(N__35113));
    Odrv12 I__6927 (
            .O(N__35113),
            .I(buf_data_vac_7));
    InMux I__6926 (
            .O(N__35110),
            .I(N__35107));
    LocalMux I__6925 (
            .O(N__35107),
            .I(N__35104));
    Span4Mux_h I__6924 (
            .O(N__35104),
            .I(N__35101));
    Odrv4 I__6923 (
            .O(N__35101),
            .I(comm_buf_5_7));
    InMux I__6922 (
            .O(N__35098),
            .I(N__35095));
    LocalMux I__6921 (
            .O(N__35095),
            .I(N__35092));
    Span4Mux_h I__6920 (
            .O(N__35092),
            .I(N__35089));
    Odrv4 I__6919 (
            .O(N__35089),
            .I(comm_buf_4_2));
    InMux I__6918 (
            .O(N__35086),
            .I(N__35083));
    LocalMux I__6917 (
            .O(N__35083),
            .I(N__35079));
    InMux I__6916 (
            .O(N__35082),
            .I(N__35076));
    Span4Mux_v I__6915 (
            .O(N__35079),
            .I(N__35073));
    LocalMux I__6914 (
            .O(N__35076),
            .I(N__35070));
    Span4Mux_h I__6913 (
            .O(N__35073),
            .I(N__35067));
    Odrv4 I__6912 (
            .O(N__35070),
            .I(comm_buf_6_2));
    Odrv4 I__6911 (
            .O(N__35067),
            .I(comm_buf_6_2));
    CascadeMux I__6910 (
            .O(N__35062),
            .I(n4_adj_1568_cascade_));
    InMux I__6909 (
            .O(N__35059),
            .I(N__35056));
    LocalMux I__6908 (
            .O(N__35056),
            .I(n20786));
    InMux I__6907 (
            .O(N__35053),
            .I(N__35050));
    LocalMux I__6906 (
            .O(N__35050),
            .I(n4_adj_1560));
    CascadeMux I__6905 (
            .O(N__35047),
            .I(n21276_cascade_));
    InMux I__6904 (
            .O(N__35044),
            .I(N__35041));
    LocalMux I__6903 (
            .O(N__35041),
            .I(n22105));
    InMux I__6902 (
            .O(N__35038),
            .I(N__35035));
    LocalMux I__6901 (
            .O(N__35035),
            .I(N__35032));
    Span4Mux_h I__6900 (
            .O(N__35032),
            .I(N__35029));
    Odrv4 I__6899 (
            .O(N__35029),
            .I(comm_buf_3_2));
    CascadeMux I__6898 (
            .O(N__35026),
            .I(n21985_cascade_));
    CascadeMux I__6897 (
            .O(N__35023),
            .I(n21988_cascade_));
    InMux I__6896 (
            .O(N__35020),
            .I(N__35017));
    LocalMux I__6895 (
            .O(N__35017),
            .I(N__35014));
    Span4Mux_v I__6894 (
            .O(N__35014),
            .I(N__35011));
    Odrv4 I__6893 (
            .O(N__35011),
            .I(comm_buf_3_0));
    CascadeMux I__6892 (
            .O(N__35008),
            .I(n17304_cascade_));
    CascadeMux I__6891 (
            .O(N__35005),
            .I(n20906_cascade_));
    InMux I__6890 (
            .O(N__35002),
            .I(N__34999));
    LocalMux I__6889 (
            .O(N__34999),
            .I(\ADC_VDC.genclk.n27_adj_1402 ));
    InMux I__6888 (
            .O(N__34996),
            .I(N__34991));
    InMux I__6887 (
            .O(N__34995),
            .I(N__34988));
    InMux I__6886 (
            .O(N__34994),
            .I(N__34985));
    LocalMux I__6885 (
            .O(N__34991),
            .I(N__34980));
    LocalMux I__6884 (
            .O(N__34988),
            .I(N__34980));
    LocalMux I__6883 (
            .O(N__34985),
            .I(\comm_spi.n14586 ));
    Odrv4 I__6882 (
            .O(N__34980),
            .I(\comm_spi.n14586 ));
    CascadeMux I__6881 (
            .O(N__34975),
            .I(N__34971));
    InMux I__6880 (
            .O(N__34974),
            .I(N__34967));
    InMux I__6879 (
            .O(N__34971),
            .I(N__34964));
    InMux I__6878 (
            .O(N__34970),
            .I(N__34959));
    LocalMux I__6877 (
            .O(N__34967),
            .I(N__34956));
    LocalMux I__6876 (
            .O(N__34964),
            .I(N__34953));
    InMux I__6875 (
            .O(N__34963),
            .I(N__34950));
    InMux I__6874 (
            .O(N__34962),
            .I(N__34947));
    LocalMux I__6873 (
            .O(N__34959),
            .I(\ADC_VDC.genclk.div_state_0 ));
    Odrv4 I__6872 (
            .O(N__34956),
            .I(\ADC_VDC.genclk.div_state_0 ));
    Odrv12 I__6871 (
            .O(N__34953),
            .I(\ADC_VDC.genclk.div_state_0 ));
    LocalMux I__6870 (
            .O(N__34950),
            .I(\ADC_VDC.genclk.div_state_0 ));
    LocalMux I__6869 (
            .O(N__34947),
            .I(\ADC_VDC.genclk.div_state_0 ));
    CascadeMux I__6868 (
            .O(N__34936),
            .I(N__34932));
    InMux I__6867 (
            .O(N__34935),
            .I(N__34927));
    InMux I__6866 (
            .O(N__34932),
            .I(N__34922));
    InMux I__6865 (
            .O(N__34931),
            .I(N__34922));
    InMux I__6864 (
            .O(N__34930),
            .I(N__34919));
    LocalMux I__6863 (
            .O(N__34927),
            .I(N__34915));
    LocalMux I__6862 (
            .O(N__34922),
            .I(N__34908));
    LocalMux I__6861 (
            .O(N__34919),
            .I(N__34908));
    InMux I__6860 (
            .O(N__34918),
            .I(N__34905));
    Span4Mux_h I__6859 (
            .O(N__34915),
            .I(N__34902));
    InMux I__6858 (
            .O(N__34914),
            .I(N__34897));
    InMux I__6857 (
            .O(N__34913),
            .I(N__34897));
    Span4Mux_h I__6856 (
            .O(N__34908),
            .I(N__34894));
    LocalMux I__6855 (
            .O(N__34905),
            .I(\ADC_VDC.genclk.div_state_1 ));
    Odrv4 I__6854 (
            .O(N__34902),
            .I(\ADC_VDC.genclk.div_state_1 ));
    LocalMux I__6853 (
            .O(N__34897),
            .I(\ADC_VDC.genclk.div_state_1 ));
    Odrv4 I__6852 (
            .O(N__34894),
            .I(\ADC_VDC.genclk.div_state_1 ));
    CEMux I__6851 (
            .O(N__34885),
            .I(N__34882));
    LocalMux I__6850 (
            .O(N__34882),
            .I(\ADC_VDC.genclk.n6 ));
    CascadeMux I__6849 (
            .O(N__34879),
            .I(N__34873));
    CascadeMux I__6848 (
            .O(N__34878),
            .I(N__34869));
    CascadeMux I__6847 (
            .O(N__34877),
            .I(N__34866));
    InMux I__6846 (
            .O(N__34876),
            .I(N__34861));
    InMux I__6845 (
            .O(N__34873),
            .I(N__34858));
    InMux I__6844 (
            .O(N__34872),
            .I(N__34855));
    InMux I__6843 (
            .O(N__34869),
            .I(N__34850));
    InMux I__6842 (
            .O(N__34866),
            .I(N__34850));
    InMux I__6841 (
            .O(N__34865),
            .I(N__34847));
    CascadeMux I__6840 (
            .O(N__34864),
            .I(N__34841));
    LocalMux I__6839 (
            .O(N__34861),
            .I(N__34838));
    LocalMux I__6838 (
            .O(N__34858),
            .I(N__34835));
    LocalMux I__6837 (
            .O(N__34855),
            .I(N__34832));
    LocalMux I__6836 (
            .O(N__34850),
            .I(N__34827));
    LocalMux I__6835 (
            .O(N__34847),
            .I(N__34827));
    InMux I__6834 (
            .O(N__34846),
            .I(N__34820));
    InMux I__6833 (
            .O(N__34845),
            .I(N__34820));
    InMux I__6832 (
            .O(N__34844),
            .I(N__34820));
    InMux I__6831 (
            .O(N__34841),
            .I(N__34817));
    Span4Mux_v I__6830 (
            .O(N__34838),
            .I(N__34812));
    Span4Mux_v I__6829 (
            .O(N__34835),
            .I(N__34812));
    Span4Mux_h I__6828 (
            .O(N__34832),
            .I(N__34805));
    Span4Mux_v I__6827 (
            .O(N__34827),
            .I(N__34805));
    LocalMux I__6826 (
            .O(N__34820),
            .I(N__34805));
    LocalMux I__6825 (
            .O(N__34817),
            .I(N__34802));
    Span4Mux_v I__6824 (
            .O(N__34812),
            .I(N__34799));
    Span4Mux_h I__6823 (
            .O(N__34805),
            .I(N__34796));
    Span12Mux_v I__6822 (
            .O(N__34802),
            .I(N__34793));
    Span4Mux_h I__6821 (
            .O(N__34799),
            .I(N__34790));
    Span4Mux_v I__6820 (
            .O(N__34796),
            .I(N__34787));
    Span12Mux_h I__6819 (
            .O(N__34793),
            .I(N__34784));
    Sp12to4 I__6818 (
            .O(N__34790),
            .I(N__34779));
    Sp12to4 I__6817 (
            .O(N__34787),
            .I(N__34779));
    Odrv12 I__6816 (
            .O(N__34784),
            .I(VDC_SDO));
    Odrv12 I__6815 (
            .O(N__34779),
            .I(VDC_SDO));
    InMux I__6814 (
            .O(N__34774),
            .I(N__34765));
    InMux I__6813 (
            .O(N__34773),
            .I(N__34762));
    InMux I__6812 (
            .O(N__34772),
            .I(N__34755));
    InMux I__6811 (
            .O(N__34771),
            .I(N__34755));
    InMux I__6810 (
            .O(N__34770),
            .I(N__34755));
    InMux I__6809 (
            .O(N__34769),
            .I(N__34752));
    CascadeMux I__6808 (
            .O(N__34768),
            .I(N__34748));
    LocalMux I__6807 (
            .O(N__34765),
            .I(N__34736));
    LocalMux I__6806 (
            .O(N__34762),
            .I(N__34731));
    LocalMux I__6805 (
            .O(N__34755),
            .I(N__34731));
    LocalMux I__6804 (
            .O(N__34752),
            .I(N__34728));
    CascadeMux I__6803 (
            .O(N__34751),
            .I(N__34725));
    InMux I__6802 (
            .O(N__34748),
            .I(N__34720));
    InMux I__6801 (
            .O(N__34747),
            .I(N__34717));
    CascadeMux I__6800 (
            .O(N__34746),
            .I(N__34713));
    InMux I__6799 (
            .O(N__34745),
            .I(N__34709));
    InMux I__6798 (
            .O(N__34744),
            .I(N__34704));
    InMux I__6797 (
            .O(N__34743),
            .I(N__34704));
    InMux I__6796 (
            .O(N__34742),
            .I(N__34701));
    InMux I__6795 (
            .O(N__34741),
            .I(N__34698));
    InMux I__6794 (
            .O(N__34740),
            .I(N__34693));
    InMux I__6793 (
            .O(N__34739),
            .I(N__34693));
    Span4Mux_v I__6792 (
            .O(N__34736),
            .I(N__34686));
    Span4Mux_v I__6791 (
            .O(N__34731),
            .I(N__34686));
    Span4Mux_v I__6790 (
            .O(N__34728),
            .I(N__34686));
    InMux I__6789 (
            .O(N__34725),
            .I(N__34679));
    InMux I__6788 (
            .O(N__34724),
            .I(N__34679));
    InMux I__6787 (
            .O(N__34723),
            .I(N__34679));
    LocalMux I__6786 (
            .O(N__34720),
            .I(N__34674));
    LocalMux I__6785 (
            .O(N__34717),
            .I(N__34674));
    InMux I__6784 (
            .O(N__34716),
            .I(N__34667));
    InMux I__6783 (
            .O(N__34713),
            .I(N__34667));
    InMux I__6782 (
            .O(N__34712),
            .I(N__34667));
    LocalMux I__6781 (
            .O(N__34709),
            .I(\ADC_VDC.adc_state_0 ));
    LocalMux I__6780 (
            .O(N__34704),
            .I(\ADC_VDC.adc_state_0 ));
    LocalMux I__6779 (
            .O(N__34701),
            .I(\ADC_VDC.adc_state_0 ));
    LocalMux I__6778 (
            .O(N__34698),
            .I(\ADC_VDC.adc_state_0 ));
    LocalMux I__6777 (
            .O(N__34693),
            .I(\ADC_VDC.adc_state_0 ));
    Odrv4 I__6776 (
            .O(N__34686),
            .I(\ADC_VDC.adc_state_0 ));
    LocalMux I__6775 (
            .O(N__34679),
            .I(\ADC_VDC.adc_state_0 ));
    Odrv4 I__6774 (
            .O(N__34674),
            .I(\ADC_VDC.adc_state_0 ));
    LocalMux I__6773 (
            .O(N__34667),
            .I(\ADC_VDC.adc_state_0 ));
    InMux I__6772 (
            .O(N__34648),
            .I(N__34645));
    LocalMux I__6771 (
            .O(N__34645),
            .I(\ADC_VDC.n62 ));
    CascadeMux I__6770 (
            .O(N__34642),
            .I(N__34621));
    InMux I__6769 (
            .O(N__34641),
            .I(N__34617));
    InMux I__6768 (
            .O(N__34640),
            .I(N__34602));
    InMux I__6767 (
            .O(N__34639),
            .I(N__34602));
    InMux I__6766 (
            .O(N__34638),
            .I(N__34602));
    InMux I__6765 (
            .O(N__34637),
            .I(N__34602));
    InMux I__6764 (
            .O(N__34636),
            .I(N__34602));
    InMux I__6763 (
            .O(N__34635),
            .I(N__34602));
    InMux I__6762 (
            .O(N__34634),
            .I(N__34602));
    InMux I__6761 (
            .O(N__34633),
            .I(N__34595));
    InMux I__6760 (
            .O(N__34632),
            .I(N__34595));
    InMux I__6759 (
            .O(N__34631),
            .I(N__34595));
    CascadeMux I__6758 (
            .O(N__34630),
            .I(N__34590));
    InMux I__6757 (
            .O(N__34629),
            .I(N__34585));
    InMux I__6756 (
            .O(N__34628),
            .I(N__34575));
    InMux I__6755 (
            .O(N__34627),
            .I(N__34575));
    InMux I__6754 (
            .O(N__34626),
            .I(N__34575));
    InMux I__6753 (
            .O(N__34625),
            .I(N__34575));
    InMux I__6752 (
            .O(N__34624),
            .I(N__34556));
    InMux I__6751 (
            .O(N__34621),
            .I(N__34556));
    CascadeMux I__6750 (
            .O(N__34620),
            .I(N__34553));
    LocalMux I__6749 (
            .O(N__34617),
            .I(N__34546));
    LocalMux I__6748 (
            .O(N__34602),
            .I(N__34546));
    LocalMux I__6747 (
            .O(N__34595),
            .I(N__34546));
    InMux I__6746 (
            .O(N__34594),
            .I(N__34541));
    InMux I__6745 (
            .O(N__34593),
            .I(N__34541));
    InMux I__6744 (
            .O(N__34590),
            .I(N__34536));
    InMux I__6743 (
            .O(N__34589),
            .I(N__34536));
    InMux I__6742 (
            .O(N__34588),
            .I(N__34533));
    LocalMux I__6741 (
            .O(N__34585),
            .I(N__34530));
    InMux I__6740 (
            .O(N__34584),
            .I(N__34527));
    LocalMux I__6739 (
            .O(N__34575),
            .I(N__34524));
    InMux I__6738 (
            .O(N__34574),
            .I(N__34507));
    InMux I__6737 (
            .O(N__34573),
            .I(N__34507));
    InMux I__6736 (
            .O(N__34572),
            .I(N__34507));
    InMux I__6735 (
            .O(N__34571),
            .I(N__34507));
    InMux I__6734 (
            .O(N__34570),
            .I(N__34507));
    InMux I__6733 (
            .O(N__34569),
            .I(N__34507));
    InMux I__6732 (
            .O(N__34568),
            .I(N__34507));
    InMux I__6731 (
            .O(N__34567),
            .I(N__34507));
    InMux I__6730 (
            .O(N__34566),
            .I(N__34504));
    CascadeMux I__6729 (
            .O(N__34565),
            .I(N__34500));
    CascadeMux I__6728 (
            .O(N__34564),
            .I(N__34497));
    CascadeMux I__6727 (
            .O(N__34563),
            .I(N__34494));
    CascadeMux I__6726 (
            .O(N__34562),
            .I(N__34491));
    CascadeMux I__6725 (
            .O(N__34561),
            .I(N__34482));
    LocalMux I__6724 (
            .O(N__34556),
            .I(N__34479));
    InMux I__6723 (
            .O(N__34553),
            .I(N__34476));
    Span4Mux_v I__6722 (
            .O(N__34546),
            .I(N__34467));
    LocalMux I__6721 (
            .O(N__34541),
            .I(N__34467));
    LocalMux I__6720 (
            .O(N__34536),
            .I(N__34467));
    LocalMux I__6719 (
            .O(N__34533),
            .I(N__34467));
    Span4Mux_h I__6718 (
            .O(N__34530),
            .I(N__34456));
    LocalMux I__6717 (
            .O(N__34527),
            .I(N__34456));
    Span4Mux_h I__6716 (
            .O(N__34524),
            .I(N__34456));
    LocalMux I__6715 (
            .O(N__34507),
            .I(N__34456));
    LocalMux I__6714 (
            .O(N__34504),
            .I(N__34453));
    InMux I__6713 (
            .O(N__34503),
            .I(N__34446));
    InMux I__6712 (
            .O(N__34500),
            .I(N__34446));
    InMux I__6711 (
            .O(N__34497),
            .I(N__34446));
    InMux I__6710 (
            .O(N__34494),
            .I(N__34443));
    InMux I__6709 (
            .O(N__34491),
            .I(N__34436));
    InMux I__6708 (
            .O(N__34490),
            .I(N__34436));
    InMux I__6707 (
            .O(N__34489),
            .I(N__34436));
    InMux I__6706 (
            .O(N__34488),
            .I(N__34425));
    InMux I__6705 (
            .O(N__34487),
            .I(N__34425));
    InMux I__6704 (
            .O(N__34486),
            .I(N__34425));
    InMux I__6703 (
            .O(N__34485),
            .I(N__34425));
    InMux I__6702 (
            .O(N__34482),
            .I(N__34425));
    Span4Mux_h I__6701 (
            .O(N__34479),
            .I(N__34418));
    LocalMux I__6700 (
            .O(N__34476),
            .I(N__34418));
    Span4Mux_h I__6699 (
            .O(N__34467),
            .I(N__34418));
    InMux I__6698 (
            .O(N__34466),
            .I(N__34413));
    InMux I__6697 (
            .O(N__34465),
            .I(N__34413));
    Span4Mux_v I__6696 (
            .O(N__34456),
            .I(N__34406));
    Span4Mux_v I__6695 (
            .O(N__34453),
            .I(N__34406));
    LocalMux I__6694 (
            .O(N__34446),
            .I(N__34406));
    LocalMux I__6693 (
            .O(N__34443),
            .I(adc_state_2));
    LocalMux I__6692 (
            .O(N__34436),
            .I(adc_state_2));
    LocalMux I__6691 (
            .O(N__34425),
            .I(adc_state_2));
    Odrv4 I__6690 (
            .O(N__34418),
            .I(adc_state_2));
    LocalMux I__6689 (
            .O(N__34413),
            .I(adc_state_2));
    Odrv4 I__6688 (
            .O(N__34406),
            .I(adc_state_2));
    CascadeMux I__6687 (
            .O(N__34393),
            .I(N__34390));
    InMux I__6686 (
            .O(N__34390),
            .I(N__34387));
    LocalMux I__6685 (
            .O(N__34387),
            .I(N__34381));
    InMux I__6684 (
            .O(N__34386),
            .I(N__34376));
    InMux I__6683 (
            .O(N__34385),
            .I(N__34376));
    CascadeMux I__6682 (
            .O(N__34384),
            .I(N__34357));
    Span4Mux_h I__6681 (
            .O(N__34381),
            .I(N__34350));
    LocalMux I__6680 (
            .O(N__34376),
            .I(N__34350));
    InMux I__6679 (
            .O(N__34375),
            .I(N__34347));
    InMux I__6678 (
            .O(N__34374),
            .I(N__34336));
    InMux I__6677 (
            .O(N__34373),
            .I(N__34336));
    InMux I__6676 (
            .O(N__34372),
            .I(N__34336));
    InMux I__6675 (
            .O(N__34371),
            .I(N__34336));
    InMux I__6674 (
            .O(N__34370),
            .I(N__34336));
    InMux I__6673 (
            .O(N__34369),
            .I(N__34333));
    InMux I__6672 (
            .O(N__34368),
            .I(N__34330));
    InMux I__6671 (
            .O(N__34367),
            .I(N__34317));
    InMux I__6670 (
            .O(N__34366),
            .I(N__34317));
    InMux I__6669 (
            .O(N__34365),
            .I(N__34317));
    InMux I__6668 (
            .O(N__34364),
            .I(N__34317));
    InMux I__6667 (
            .O(N__34363),
            .I(N__34317));
    InMux I__6666 (
            .O(N__34362),
            .I(N__34317));
    InMux I__6665 (
            .O(N__34361),
            .I(N__34314));
    InMux I__6664 (
            .O(N__34360),
            .I(N__34311));
    InMux I__6663 (
            .O(N__34357),
            .I(N__34308));
    CascadeMux I__6662 (
            .O(N__34356),
            .I(N__34296));
    InMux I__6661 (
            .O(N__34355),
            .I(N__34286));
    Span4Mux_v I__6660 (
            .O(N__34350),
            .I(N__34281));
    LocalMux I__6659 (
            .O(N__34347),
            .I(N__34281));
    LocalMux I__6658 (
            .O(N__34336),
            .I(N__34276));
    LocalMux I__6657 (
            .O(N__34333),
            .I(N__34276));
    LocalMux I__6656 (
            .O(N__34330),
            .I(N__34273));
    LocalMux I__6655 (
            .O(N__34317),
            .I(N__34268));
    LocalMux I__6654 (
            .O(N__34314),
            .I(N__34268));
    LocalMux I__6653 (
            .O(N__34311),
            .I(N__34263));
    LocalMux I__6652 (
            .O(N__34308),
            .I(N__34263));
    InMux I__6651 (
            .O(N__34307),
            .I(N__34252));
    InMux I__6650 (
            .O(N__34306),
            .I(N__34239));
    InMux I__6649 (
            .O(N__34305),
            .I(N__34239));
    InMux I__6648 (
            .O(N__34304),
            .I(N__34239));
    InMux I__6647 (
            .O(N__34303),
            .I(N__34239));
    InMux I__6646 (
            .O(N__34302),
            .I(N__34239));
    InMux I__6645 (
            .O(N__34301),
            .I(N__34239));
    InMux I__6644 (
            .O(N__34300),
            .I(N__34236));
    InMux I__6643 (
            .O(N__34299),
            .I(N__34233));
    InMux I__6642 (
            .O(N__34296),
            .I(N__34224));
    InMux I__6641 (
            .O(N__34295),
            .I(N__34224));
    InMux I__6640 (
            .O(N__34294),
            .I(N__34224));
    InMux I__6639 (
            .O(N__34293),
            .I(N__34224));
    InMux I__6638 (
            .O(N__34292),
            .I(N__34215));
    InMux I__6637 (
            .O(N__34291),
            .I(N__34215));
    InMux I__6636 (
            .O(N__34290),
            .I(N__34215));
    InMux I__6635 (
            .O(N__34289),
            .I(N__34215));
    LocalMux I__6634 (
            .O(N__34286),
            .I(N__34210));
    Span4Mux_h I__6633 (
            .O(N__34281),
            .I(N__34210));
    Span4Mux_v I__6632 (
            .O(N__34276),
            .I(N__34201));
    Span4Mux_v I__6631 (
            .O(N__34273),
            .I(N__34201));
    Span4Mux_v I__6630 (
            .O(N__34268),
            .I(N__34201));
    Span4Mux_h I__6629 (
            .O(N__34263),
            .I(N__34201));
    InMux I__6628 (
            .O(N__34262),
            .I(N__34184));
    InMux I__6627 (
            .O(N__34261),
            .I(N__34184));
    InMux I__6626 (
            .O(N__34260),
            .I(N__34184));
    InMux I__6625 (
            .O(N__34259),
            .I(N__34184));
    InMux I__6624 (
            .O(N__34258),
            .I(N__34184));
    InMux I__6623 (
            .O(N__34257),
            .I(N__34184));
    InMux I__6622 (
            .O(N__34256),
            .I(N__34184));
    InMux I__6621 (
            .O(N__34255),
            .I(N__34184));
    LocalMux I__6620 (
            .O(N__34252),
            .I(N__34181));
    LocalMux I__6619 (
            .O(N__34239),
            .I(adc_state_3));
    LocalMux I__6618 (
            .O(N__34236),
            .I(adc_state_3));
    LocalMux I__6617 (
            .O(N__34233),
            .I(adc_state_3));
    LocalMux I__6616 (
            .O(N__34224),
            .I(adc_state_3));
    LocalMux I__6615 (
            .O(N__34215),
            .I(adc_state_3));
    Odrv4 I__6614 (
            .O(N__34210),
            .I(adc_state_3));
    Odrv4 I__6613 (
            .O(N__34201),
            .I(adc_state_3));
    LocalMux I__6612 (
            .O(N__34184),
            .I(adc_state_3));
    Odrv4 I__6611 (
            .O(N__34181),
            .I(adc_state_3));
    CascadeMux I__6610 (
            .O(N__34162),
            .I(\ADC_VDC.n62_cascade_ ));
    InMux I__6609 (
            .O(N__34159),
            .I(N__34142));
    InMux I__6608 (
            .O(N__34158),
            .I(N__34142));
    InMux I__6607 (
            .O(N__34157),
            .I(N__34136));
    InMux I__6606 (
            .O(N__34156),
            .I(N__34136));
    InMux I__6605 (
            .O(N__34155),
            .I(N__34133));
    InMux I__6604 (
            .O(N__34154),
            .I(N__34128));
    InMux I__6603 (
            .O(N__34153),
            .I(N__34128));
    InMux I__6602 (
            .O(N__34152),
            .I(N__34123));
    InMux I__6601 (
            .O(N__34151),
            .I(N__34123));
    InMux I__6600 (
            .O(N__34150),
            .I(N__34115));
    InMux I__6599 (
            .O(N__34149),
            .I(N__34115));
    CascadeMux I__6598 (
            .O(N__34148),
            .I(N__34109));
    CascadeMux I__6597 (
            .O(N__34147),
            .I(N__34106));
    LocalMux I__6596 (
            .O(N__34142),
            .I(N__34103));
    InMux I__6595 (
            .O(N__34141),
            .I(N__34100));
    LocalMux I__6594 (
            .O(N__34136),
            .I(N__34097));
    LocalMux I__6593 (
            .O(N__34133),
            .I(N__34089));
    LocalMux I__6592 (
            .O(N__34128),
            .I(N__34089));
    LocalMux I__6591 (
            .O(N__34123),
            .I(N__34086));
    InMux I__6590 (
            .O(N__34122),
            .I(N__34083));
    InMux I__6589 (
            .O(N__34121),
            .I(N__34080));
    InMux I__6588 (
            .O(N__34120),
            .I(N__34077));
    LocalMux I__6587 (
            .O(N__34115),
            .I(N__34074));
    InMux I__6586 (
            .O(N__34114),
            .I(N__34071));
    InMux I__6585 (
            .O(N__34113),
            .I(N__34066));
    InMux I__6584 (
            .O(N__34112),
            .I(N__34066));
    InMux I__6583 (
            .O(N__34109),
            .I(N__34063));
    InMux I__6582 (
            .O(N__34106),
            .I(N__34060));
    Span4Mux_v I__6581 (
            .O(N__34103),
            .I(N__34057));
    LocalMux I__6580 (
            .O(N__34100),
            .I(N__34052));
    Span4Mux_h I__6579 (
            .O(N__34097),
            .I(N__34052));
    InMux I__6578 (
            .O(N__34096),
            .I(N__34045));
    InMux I__6577 (
            .O(N__34095),
            .I(N__34045));
    InMux I__6576 (
            .O(N__34094),
            .I(N__34045));
    Span4Mux_v I__6575 (
            .O(N__34089),
            .I(N__34042));
    Span4Mux_h I__6574 (
            .O(N__34086),
            .I(N__34037));
    LocalMux I__6573 (
            .O(N__34083),
            .I(N__34037));
    LocalMux I__6572 (
            .O(N__34080),
            .I(\ADC_VDC.adc_state_1 ));
    LocalMux I__6571 (
            .O(N__34077),
            .I(\ADC_VDC.adc_state_1 ));
    Odrv12 I__6570 (
            .O(N__34074),
            .I(\ADC_VDC.adc_state_1 ));
    LocalMux I__6569 (
            .O(N__34071),
            .I(\ADC_VDC.adc_state_1 ));
    LocalMux I__6568 (
            .O(N__34066),
            .I(\ADC_VDC.adc_state_1 ));
    LocalMux I__6567 (
            .O(N__34063),
            .I(\ADC_VDC.adc_state_1 ));
    LocalMux I__6566 (
            .O(N__34060),
            .I(\ADC_VDC.adc_state_1 ));
    Odrv4 I__6565 (
            .O(N__34057),
            .I(\ADC_VDC.adc_state_1 ));
    Odrv4 I__6564 (
            .O(N__34052),
            .I(\ADC_VDC.adc_state_1 ));
    LocalMux I__6563 (
            .O(N__34045),
            .I(\ADC_VDC.adc_state_1 ));
    Odrv4 I__6562 (
            .O(N__34042),
            .I(\ADC_VDC.adc_state_1 ));
    Odrv4 I__6561 (
            .O(N__34037),
            .I(\ADC_VDC.adc_state_1 ));
    CEMux I__6560 (
            .O(N__34012),
            .I(N__34009));
    LocalMux I__6559 (
            .O(N__34009),
            .I(N__34006));
    Odrv4 I__6558 (
            .O(N__34006),
            .I(\ADC_VDC.n11736 ));
    InMux I__6557 (
            .O(N__34003),
            .I(N__34000));
    LocalMux I__6556 (
            .O(N__34000),
            .I(N__33997));
    Span4Mux_h I__6555 (
            .O(N__33997),
            .I(N__33994));
    Span4Mux_h I__6554 (
            .O(N__33994),
            .I(N__33991));
    Odrv4 I__6553 (
            .O(N__33991),
            .I(comm_buf_3_7));
    InMux I__6552 (
            .O(N__33988),
            .I(N__33985));
    LocalMux I__6551 (
            .O(N__33985),
            .I(N__33982));
    Odrv4 I__6550 (
            .O(N__33982),
            .I(n1));
    CascadeMux I__6549 (
            .O(N__33979),
            .I(n2_adj_1559_cascade_));
    InMux I__6548 (
            .O(N__33976),
            .I(N__33973));
    LocalMux I__6547 (
            .O(N__33973),
            .I(N__33970));
    Span4Mux_h I__6546 (
            .O(N__33970),
            .I(N__33967));
    Odrv4 I__6545 (
            .O(N__33967),
            .I(comm_buf_4_7));
    InMux I__6544 (
            .O(N__33964),
            .I(N__33961));
    LocalMux I__6543 (
            .O(N__33961),
            .I(N__33957));
    CascadeMux I__6542 (
            .O(N__33960),
            .I(N__33954));
    Span4Mux_h I__6541 (
            .O(N__33957),
            .I(N__33951));
    InMux I__6540 (
            .O(N__33954),
            .I(N__33948));
    Span4Mux_v I__6539 (
            .O(N__33951),
            .I(N__33945));
    LocalMux I__6538 (
            .O(N__33948),
            .I(comm_buf_6_7));
    Odrv4 I__6537 (
            .O(N__33945),
            .I(comm_buf_6_7));
    InMux I__6536 (
            .O(N__33940),
            .I(n19325));
    CEMux I__6535 (
            .O(N__33937),
            .I(N__33933));
    CEMux I__6534 (
            .O(N__33936),
            .I(N__33930));
    LocalMux I__6533 (
            .O(N__33933),
            .I(N__33927));
    LocalMux I__6532 (
            .O(N__33930),
            .I(N__33924));
    Span4Mux_v I__6531 (
            .O(N__33927),
            .I(N__33918));
    Span4Mux_h I__6530 (
            .O(N__33924),
            .I(N__33918));
    CEMux I__6529 (
            .O(N__33923),
            .I(N__33915));
    Span4Mux_h I__6528 (
            .O(N__33918),
            .I(N__33911));
    LocalMux I__6527 (
            .O(N__33915),
            .I(N__33908));
    InMux I__6526 (
            .O(N__33914),
            .I(N__33905));
    Odrv4 I__6525 (
            .O(N__33911),
            .I(n11538));
    Odrv12 I__6524 (
            .O(N__33908),
            .I(n11538));
    LocalMux I__6523 (
            .O(N__33905),
            .I(n11538));
    SRMux I__6522 (
            .O(N__33898),
            .I(N__33895));
    LocalMux I__6521 (
            .O(N__33895),
            .I(N__33891));
    SRMux I__6520 (
            .O(N__33894),
            .I(N__33888));
    Span4Mux_h I__6519 (
            .O(N__33891),
            .I(N__33885));
    LocalMux I__6518 (
            .O(N__33888),
            .I(N__33882));
    Odrv4 I__6517 (
            .O(N__33885),
            .I(n14639));
    Odrv4 I__6516 (
            .O(N__33882),
            .I(n14639));
    CascadeMux I__6515 (
            .O(N__33877),
            .I(N__33874));
    InMux I__6514 (
            .O(N__33874),
            .I(N__33871));
    LocalMux I__6513 (
            .O(N__33871),
            .I(\SIG_DDS.tmp_buf_11 ));
    InMux I__6512 (
            .O(N__33868),
            .I(N__33865));
    LocalMux I__6511 (
            .O(N__33865),
            .I(N__33861));
    InMux I__6510 (
            .O(N__33864),
            .I(N__33858));
    Span4Mux_h I__6509 (
            .O(N__33861),
            .I(N__33854));
    LocalMux I__6508 (
            .O(N__33858),
            .I(N__33851));
    InMux I__6507 (
            .O(N__33857),
            .I(N__33848));
    Sp12to4 I__6506 (
            .O(N__33854),
            .I(N__33843));
    Span12Mux_h I__6505 (
            .O(N__33851),
            .I(N__33843));
    LocalMux I__6504 (
            .O(N__33848),
            .I(buf_dds0_12));
    Odrv12 I__6503 (
            .O(N__33843),
            .I(buf_dds0_12));
    CascadeMux I__6502 (
            .O(N__33838),
            .I(N__33835));
    InMux I__6501 (
            .O(N__33835),
            .I(N__33832));
    LocalMux I__6500 (
            .O(N__33832),
            .I(\SIG_DDS.tmp_buf_12 ));
    CascadeMux I__6499 (
            .O(N__33829),
            .I(N__33826));
    InMux I__6498 (
            .O(N__33826),
            .I(N__33823));
    LocalMux I__6497 (
            .O(N__33823),
            .I(\SIG_DDS.tmp_buf_1 ));
    InMux I__6496 (
            .O(N__33820),
            .I(N__33815));
    InMux I__6495 (
            .O(N__33819),
            .I(N__33812));
    InMux I__6494 (
            .O(N__33818),
            .I(N__33809));
    LocalMux I__6493 (
            .O(N__33815),
            .I(\comm_spi.n22632 ));
    LocalMux I__6492 (
            .O(N__33812),
            .I(\comm_spi.n22632 ));
    LocalMux I__6491 (
            .O(N__33809),
            .I(\comm_spi.n22632 ));
    InMux I__6490 (
            .O(N__33802),
            .I(N__33799));
    LocalMux I__6489 (
            .O(N__33799),
            .I(\comm_spi.n14600 ));
    SRMux I__6488 (
            .O(N__33796),
            .I(N__33793));
    LocalMux I__6487 (
            .O(N__33793),
            .I(N__33790));
    Sp12to4 I__6486 (
            .O(N__33790),
            .I(N__33787));
    Odrv12 I__6485 (
            .O(N__33787),
            .I(\comm_spi.DOUT_7__N_739 ));
    CascadeMux I__6484 (
            .O(N__33784),
            .I(\ADC_VDC.genclk.n21172_cascade_ ));
    InMux I__6483 (
            .O(N__33781),
            .I(N__33777));
    InMux I__6482 (
            .O(N__33780),
            .I(N__33774));
    LocalMux I__6481 (
            .O(N__33777),
            .I(\ADC_VDC.genclk.n21166 ));
    LocalMux I__6480 (
            .O(N__33774),
            .I(\ADC_VDC.genclk.n21166 ));
    InMux I__6479 (
            .O(N__33769),
            .I(N__33766));
    LocalMux I__6478 (
            .O(N__33766),
            .I(N__33763));
    Odrv4 I__6477 (
            .O(N__33763),
            .I(\ADC_VDC.genclk.n28_adj_1400 ));
    InMux I__6476 (
            .O(N__33760),
            .I(N__33757));
    LocalMux I__6475 (
            .O(N__33757),
            .I(\ADC_VDC.genclk.n26_adj_1401 ));
    CascadeMux I__6474 (
            .O(N__33754),
            .I(N__33750));
    InMux I__6473 (
            .O(N__33753),
            .I(N__33747));
    InMux I__6472 (
            .O(N__33750),
            .I(N__33744));
    LocalMux I__6471 (
            .O(N__33747),
            .I(acadc_skipcnt_6));
    LocalMux I__6470 (
            .O(N__33744),
            .I(acadc_skipcnt_6));
    InMux I__6469 (
            .O(N__33739),
            .I(n19316));
    InMux I__6468 (
            .O(N__33736),
            .I(n19317));
    InMux I__6467 (
            .O(N__33733),
            .I(N__33730));
    LocalMux I__6466 (
            .O(N__33730),
            .I(N__33726));
    InMux I__6465 (
            .O(N__33729),
            .I(N__33723));
    Span4Mux_h I__6464 (
            .O(N__33726),
            .I(N__33720));
    LocalMux I__6463 (
            .O(N__33723),
            .I(acadc_skipcnt_8));
    Odrv4 I__6462 (
            .O(N__33720),
            .I(acadc_skipcnt_8));
    InMux I__6461 (
            .O(N__33715),
            .I(n19318));
    InMux I__6460 (
            .O(N__33712),
            .I(bfn_13_18_0_));
    InMux I__6459 (
            .O(N__33709),
            .I(n19320));
    InMux I__6458 (
            .O(N__33706),
            .I(n19321));
    InMux I__6457 (
            .O(N__33703),
            .I(n19322));
    InMux I__6456 (
            .O(N__33700),
            .I(N__33697));
    LocalMux I__6455 (
            .O(N__33697),
            .I(N__33693));
    InMux I__6454 (
            .O(N__33696),
            .I(N__33690));
    Span4Mux_h I__6453 (
            .O(N__33693),
            .I(N__33687));
    LocalMux I__6452 (
            .O(N__33690),
            .I(acadc_skipcnt_13));
    Odrv4 I__6451 (
            .O(N__33687),
            .I(acadc_skipcnt_13));
    InMux I__6450 (
            .O(N__33682),
            .I(n19323));
    InMux I__6449 (
            .O(N__33679),
            .I(n19324));
    InMux I__6448 (
            .O(N__33676),
            .I(N__33672));
    InMux I__6447 (
            .O(N__33675),
            .I(N__33669));
    LocalMux I__6446 (
            .O(N__33672),
            .I(N__33666));
    LocalMux I__6445 (
            .O(N__33669),
            .I(acadc_skipcnt_1));
    Odrv4 I__6444 (
            .O(N__33666),
            .I(acadc_skipcnt_1));
    InMux I__6443 (
            .O(N__33661),
            .I(bfn_13_17_0_));
    InMux I__6442 (
            .O(N__33658),
            .I(n19312));
    InMux I__6441 (
            .O(N__33655),
            .I(N__33651));
    InMux I__6440 (
            .O(N__33654),
            .I(N__33648));
    LocalMux I__6439 (
            .O(N__33651),
            .I(N__33645));
    LocalMux I__6438 (
            .O(N__33648),
            .I(N__33640));
    Span4Mux_v I__6437 (
            .O(N__33645),
            .I(N__33640));
    Odrv4 I__6436 (
            .O(N__33640),
            .I(acadc_skipcnt_3));
    InMux I__6435 (
            .O(N__33637),
            .I(n19313));
    CascadeMux I__6434 (
            .O(N__33634),
            .I(N__33631));
    InMux I__6433 (
            .O(N__33631),
            .I(N__33627));
    InMux I__6432 (
            .O(N__33630),
            .I(N__33624));
    LocalMux I__6431 (
            .O(N__33627),
            .I(N__33621));
    LocalMux I__6430 (
            .O(N__33624),
            .I(N__33616));
    Span4Mux_h I__6429 (
            .O(N__33621),
            .I(N__33616));
    Odrv4 I__6428 (
            .O(N__33616),
            .I(acadc_skipcnt_4));
    InMux I__6427 (
            .O(N__33613),
            .I(n19314));
    InMux I__6426 (
            .O(N__33610),
            .I(N__33607));
    LocalMux I__6425 (
            .O(N__33607),
            .I(N__33603));
    InMux I__6424 (
            .O(N__33606),
            .I(N__33600));
    Span4Mux_h I__6423 (
            .O(N__33603),
            .I(N__33597));
    LocalMux I__6422 (
            .O(N__33600),
            .I(acadc_skipcnt_5));
    Odrv4 I__6421 (
            .O(N__33597),
            .I(acadc_skipcnt_5));
    InMux I__6420 (
            .O(N__33592),
            .I(n19315));
    CascadeMux I__6419 (
            .O(N__33589),
            .I(n22198_cascade_));
    CascadeMux I__6418 (
            .O(N__33586),
            .I(n30_adj_1503_cascade_));
    InMux I__6417 (
            .O(N__33583),
            .I(N__33580));
    LocalMux I__6416 (
            .O(N__33580),
            .I(N__33577));
    Span4Mux_h I__6415 (
            .O(N__33577),
            .I(N__33574));
    Odrv4 I__6414 (
            .O(N__33574),
            .I(n19_adj_1501));
    CascadeMux I__6413 (
            .O(N__33571),
            .I(N__33568));
    InMux I__6412 (
            .O(N__33568),
            .I(N__33565));
    LocalMux I__6411 (
            .O(N__33565),
            .I(N__33562));
    Span4Mux_h I__6410 (
            .O(N__33562),
            .I(N__33559));
    Sp12to4 I__6409 (
            .O(N__33559),
            .I(N__33555));
    CascadeMux I__6408 (
            .O(N__33558),
            .I(N__33552));
    Span12Mux_v I__6407 (
            .O(N__33555),
            .I(N__33549));
    InMux I__6406 (
            .O(N__33552),
            .I(N__33546));
    Odrv12 I__6405 (
            .O(N__33549),
            .I(buf_readRTD_3));
    LocalMux I__6404 (
            .O(N__33546),
            .I(buf_readRTD_3));
    InMux I__6403 (
            .O(N__33541),
            .I(N__33538));
    LocalMux I__6402 (
            .O(N__33538),
            .I(N__33535));
    Span4Mux_h I__6401 (
            .O(N__33535),
            .I(N__33530));
    InMux I__6400 (
            .O(N__33534),
            .I(N__33527));
    InMux I__6399 (
            .O(N__33533),
            .I(N__33524));
    Span4Mux_h I__6398 (
            .O(N__33530),
            .I(N__33521));
    LocalMux I__6397 (
            .O(N__33527),
            .I(buf_adcdata_iac_11));
    LocalMux I__6396 (
            .O(N__33524),
            .I(buf_adcdata_iac_11));
    Odrv4 I__6395 (
            .O(N__33521),
            .I(buf_adcdata_iac_11));
    CascadeMux I__6394 (
            .O(N__33514),
            .I(n22009_cascade_));
    InMux I__6393 (
            .O(N__33511),
            .I(N__33508));
    LocalMux I__6392 (
            .O(N__33508),
            .I(N__33505));
    Odrv12 I__6391 (
            .O(N__33505),
            .I(n16_adj_1500));
    InMux I__6390 (
            .O(N__33502),
            .I(N__33499));
    LocalMux I__6389 (
            .O(N__33499),
            .I(n22012));
    CascadeMux I__6388 (
            .O(N__33496),
            .I(N__33493));
    InMux I__6387 (
            .O(N__33493),
            .I(N__33489));
    InMux I__6386 (
            .O(N__33492),
            .I(N__33486));
    LocalMux I__6385 (
            .O(N__33489),
            .I(acadc_skipcnt_0));
    LocalMux I__6384 (
            .O(N__33486),
            .I(acadc_skipcnt_0));
    SRMux I__6383 (
            .O(N__33481),
            .I(N__33478));
    LocalMux I__6382 (
            .O(N__33478),
            .I(N__33475));
    Span4Mux_h I__6381 (
            .O(N__33475),
            .I(N__33472));
    Odrv4 I__6380 (
            .O(N__33472),
            .I(n20757));
    InMux I__6379 (
            .O(N__33469),
            .I(N__33466));
    LocalMux I__6378 (
            .O(N__33466),
            .I(N__33463));
    Span4Mux_v I__6377 (
            .O(N__33463),
            .I(N__33458));
    InMux I__6376 (
            .O(N__33462),
            .I(N__33455));
    InMux I__6375 (
            .O(N__33461),
            .I(N__33452));
    Span4Mux_h I__6374 (
            .O(N__33458),
            .I(N__33449));
    LocalMux I__6373 (
            .O(N__33455),
            .I(buf_adcdata_iac_12));
    LocalMux I__6372 (
            .O(N__33452),
            .I(buf_adcdata_iac_12));
    Odrv4 I__6371 (
            .O(N__33449),
            .I(buf_adcdata_iac_12));
    CascadeMux I__6370 (
            .O(N__33442),
            .I(n22081_cascade_));
    CascadeMux I__6369 (
            .O(N__33439),
            .I(N__33435));
    InMux I__6368 (
            .O(N__33438),
            .I(N__33432));
    InMux I__6367 (
            .O(N__33435),
            .I(N__33429));
    LocalMux I__6366 (
            .O(N__33432),
            .I(N__33426));
    LocalMux I__6365 (
            .O(N__33429),
            .I(data_idxvec_4));
    Odrv4 I__6364 (
            .O(N__33426),
            .I(data_idxvec_4));
    InMux I__6363 (
            .O(N__33421),
            .I(N__33418));
    LocalMux I__6362 (
            .O(N__33418),
            .I(N__33415));
    Span4Mux_h I__6361 (
            .O(N__33415),
            .I(N__33412));
    Odrv4 I__6360 (
            .O(N__33412),
            .I(n21261));
    CascadeMux I__6359 (
            .O(N__33409),
            .I(n26_adj_1484_cascade_));
    CascadeMux I__6358 (
            .O(N__33406),
            .I(n22159_cascade_));
    InMux I__6357 (
            .O(N__33403),
            .I(N__33400));
    LocalMux I__6356 (
            .O(N__33400),
            .I(n22084));
    CascadeMux I__6355 (
            .O(N__33397),
            .I(n22162_cascade_));
    CascadeMux I__6354 (
            .O(N__33394),
            .I(n30_adj_1493_cascade_));
    InMux I__6353 (
            .O(N__33391),
            .I(N__33387));
    InMux I__6352 (
            .O(N__33390),
            .I(N__33384));
    LocalMux I__6351 (
            .O(N__33387),
            .I(N__33381));
    LocalMux I__6350 (
            .O(N__33384),
            .I(data_idxvec_3));
    Odrv4 I__6349 (
            .O(N__33381),
            .I(data_idxvec_3));
    InMux I__6348 (
            .O(N__33376),
            .I(N__33373));
    LocalMux I__6347 (
            .O(N__33373),
            .I(N__33370));
    Span4Mux_h I__6346 (
            .O(N__33370),
            .I(N__33367));
    Span4Mux_h I__6345 (
            .O(N__33367),
            .I(N__33364));
    Odrv4 I__6344 (
            .O(N__33364),
            .I(n21285));
    CascadeMux I__6343 (
            .O(N__33361),
            .I(n26_adj_1502_cascade_));
    CascadeMux I__6342 (
            .O(N__33358),
            .I(n22195_cascade_));
    InMux I__6341 (
            .O(N__33355),
            .I(N__33350));
    InMux I__6340 (
            .O(N__33354),
            .I(N__33345));
    InMux I__6339 (
            .O(N__33353),
            .I(N__33345));
    LocalMux I__6338 (
            .O(N__33350),
            .I(acadc_skipCount_3));
    LocalMux I__6337 (
            .O(N__33345),
            .I(acadc_skipCount_3));
    CascadeMux I__6336 (
            .O(N__33340),
            .I(N__33337));
    InMux I__6335 (
            .O(N__33337),
            .I(N__33333));
    InMux I__6334 (
            .O(N__33336),
            .I(N__33330));
    LocalMux I__6333 (
            .O(N__33333),
            .I(data_idxvec_2));
    LocalMux I__6332 (
            .O(N__33330),
            .I(data_idxvec_2));
    CascadeMux I__6331 (
            .O(N__33325),
            .I(n26_adj_1506_cascade_));
    InMux I__6330 (
            .O(N__33322),
            .I(N__33319));
    LocalMux I__6329 (
            .O(N__33319),
            .I(N__33316));
    Span4Mux_v I__6328 (
            .O(N__33316),
            .I(N__33313));
    Span4Mux_h I__6327 (
            .O(N__33313),
            .I(N__33310));
    Span4Mux_h I__6326 (
            .O(N__33310),
            .I(N__33307));
    Odrv4 I__6325 (
            .O(N__33307),
            .I(buf_data_iac_10));
    CascadeMux I__6324 (
            .O(N__33304),
            .I(n20816_cascade_));
    InMux I__6323 (
            .O(N__33301),
            .I(N__33298));
    LocalMux I__6322 (
            .O(N__33298),
            .I(N__33295));
    Span4Mux_v I__6321 (
            .O(N__33295),
            .I(N__33292));
    Span4Mux_h I__6320 (
            .O(N__33292),
            .I(N__33289));
    Odrv4 I__6319 (
            .O(N__33289),
            .I(n20845));
    CascadeMux I__6318 (
            .O(N__33286),
            .I(n22087_cascade_));
    CascadeMux I__6317 (
            .O(N__33283),
            .I(n22090_cascade_));
    InMux I__6316 (
            .O(N__33280),
            .I(N__33277));
    LocalMux I__6315 (
            .O(N__33277),
            .I(N__33274));
    Odrv12 I__6314 (
            .O(N__33274),
            .I(n19_adj_1505));
    InMux I__6313 (
            .O(N__33271),
            .I(N__33268));
    LocalMux I__6312 (
            .O(N__33268),
            .I(N__33265));
    Span4Mux_v I__6311 (
            .O(N__33265),
            .I(N__33262));
    Span4Mux_h I__6310 (
            .O(N__33262),
            .I(N__33258));
    CascadeMux I__6309 (
            .O(N__33261),
            .I(N__33255));
    Span4Mux_h I__6308 (
            .O(N__33258),
            .I(N__33252));
    InMux I__6307 (
            .O(N__33255),
            .I(N__33249));
    Odrv4 I__6306 (
            .O(N__33252),
            .I(buf_readRTD_2));
    LocalMux I__6305 (
            .O(N__33249),
            .I(buf_readRTD_2));
    InMux I__6304 (
            .O(N__33244),
            .I(N__33241));
    LocalMux I__6303 (
            .O(N__33241),
            .I(n20846));
    InMux I__6302 (
            .O(N__33238),
            .I(N__33235));
    LocalMux I__6301 (
            .O(N__33235),
            .I(n20815));
    InMux I__6300 (
            .O(N__33232),
            .I(N__33229));
    LocalMux I__6299 (
            .O(N__33229),
            .I(N__33226));
    Span4Mux_v I__6298 (
            .O(N__33226),
            .I(N__33223));
    Span4Mux_h I__6297 (
            .O(N__33223),
            .I(N__33220));
    Odrv4 I__6296 (
            .O(N__33220),
            .I(n19));
    CascadeMux I__6295 (
            .O(N__33217),
            .I(N__33214));
    InMux I__6294 (
            .O(N__33214),
            .I(N__33211));
    LocalMux I__6293 (
            .O(N__33211),
            .I(N__33208));
    Span4Mux_v I__6292 (
            .O(N__33208),
            .I(N__33204));
    CascadeMux I__6291 (
            .O(N__33207),
            .I(N__33201));
    Sp12to4 I__6290 (
            .O(N__33204),
            .I(N__33198));
    InMux I__6289 (
            .O(N__33201),
            .I(N__33195));
    Odrv12 I__6288 (
            .O(N__33198),
            .I(buf_readRTD_4));
    LocalMux I__6287 (
            .O(N__33195),
            .I(buf_readRTD_4));
    InMux I__6286 (
            .O(N__33190),
            .I(N__33187));
    LocalMux I__6285 (
            .O(N__33187),
            .I(N__33184));
    Span4Mux_v I__6284 (
            .O(N__33184),
            .I(N__33181));
    Span4Mux_h I__6283 (
            .O(N__33181),
            .I(N__33178));
    Odrv4 I__6282 (
            .O(N__33178),
            .I(comm_buf_3_5));
    CascadeMux I__6281 (
            .O(N__33175),
            .I(n17331_cascade_));
    CascadeMux I__6280 (
            .O(N__33172),
            .I(n20903_cascade_));
    CascadeMux I__6279 (
            .O(N__33169),
            .I(n1_adj_1561_cascade_));
    CascadeMux I__6278 (
            .O(N__33166),
            .I(N__33163));
    InMux I__6277 (
            .O(N__33163),
            .I(N__33159));
    InMux I__6276 (
            .O(N__33162),
            .I(N__33156));
    LocalMux I__6275 (
            .O(N__33159),
            .I(N__33151));
    LocalMux I__6274 (
            .O(N__33156),
            .I(N__33151));
    Odrv12 I__6273 (
            .O(N__33151),
            .I(comm_buf_6_6));
    CascadeMux I__6272 (
            .O(N__33148),
            .I(N__33145));
    InMux I__6271 (
            .O(N__33145),
            .I(N__33142));
    LocalMux I__6270 (
            .O(N__33142),
            .I(N__33139));
    Span4Mux_v I__6269 (
            .O(N__33139),
            .I(N__33136));
    Odrv4 I__6268 (
            .O(N__33136),
            .I(comm_buf_3_6));
    InMux I__6267 (
            .O(N__33133),
            .I(N__33130));
    LocalMux I__6266 (
            .O(N__33130),
            .I(n2_adj_1562));
    InMux I__6265 (
            .O(N__33127),
            .I(N__33124));
    LocalMux I__6264 (
            .O(N__33124),
            .I(comm_buf_4_6));
    InMux I__6263 (
            .O(N__33121),
            .I(N__33118));
    LocalMux I__6262 (
            .O(N__33118),
            .I(n21051));
    CascadeMux I__6261 (
            .O(N__33115),
            .I(n4_adj_1563_cascade_));
    InMux I__6260 (
            .O(N__33112),
            .I(N__33109));
    LocalMux I__6259 (
            .O(N__33109),
            .I(n22093));
    SRMux I__6258 (
            .O(N__33106),
            .I(N__33103));
    LocalMux I__6257 (
            .O(N__33103),
            .I(n14763));
    CascadeMux I__6256 (
            .O(N__33100),
            .I(N__33097));
    InMux I__6255 (
            .O(N__33097),
            .I(N__33094));
    LocalMux I__6254 (
            .O(N__33094),
            .I(N__33091));
    Span4Mux_h I__6253 (
            .O(N__33091),
            .I(N__33088));
    Odrv4 I__6252 (
            .O(N__33088),
            .I(comm_buf_3_3));
    CascadeMux I__6251 (
            .O(N__33085),
            .I(n21979_cascade_));
    InMux I__6250 (
            .O(N__33082),
            .I(N__33079));
    LocalMux I__6249 (
            .O(N__33079),
            .I(comm_buf_4_3));
    InMux I__6248 (
            .O(N__33076),
            .I(N__33072));
    InMux I__6247 (
            .O(N__33075),
            .I(N__33069));
    LocalMux I__6246 (
            .O(N__33072),
            .I(N__33066));
    LocalMux I__6245 (
            .O(N__33069),
            .I(comm_buf_6_3));
    Odrv4 I__6244 (
            .O(N__33066),
            .I(comm_buf_6_3));
    CascadeMux I__6243 (
            .O(N__33061),
            .I(n4_adj_1567_cascade_));
    CascadeMux I__6242 (
            .O(N__33058),
            .I(n20783_cascade_));
    InMux I__6241 (
            .O(N__33055),
            .I(N__33052));
    LocalMux I__6240 (
            .O(N__33052),
            .I(n21982));
    SRMux I__6239 (
            .O(N__33049),
            .I(N__33046));
    LocalMux I__6238 (
            .O(N__33046),
            .I(N__33043));
    Odrv12 I__6237 (
            .O(N__33043),
            .I(\comm_spi.data_tx_7__N_762 ));
    CEMux I__6236 (
            .O(N__33040),
            .I(N__33037));
    LocalMux I__6235 (
            .O(N__33037),
            .I(n11727));
    InMux I__6234 (
            .O(N__33034),
            .I(N__33024));
    InMux I__6233 (
            .O(N__33033),
            .I(N__33024));
    InMux I__6232 (
            .O(N__33032),
            .I(N__33024));
    InMux I__6231 (
            .O(N__33031),
            .I(N__33021));
    LocalMux I__6230 (
            .O(N__33024),
            .I(\comm_spi.bit_cnt_1 ));
    LocalMux I__6229 (
            .O(N__33021),
            .I(\comm_spi.bit_cnt_1 ));
    CascadeMux I__6228 (
            .O(N__33016),
            .I(N__33012));
    InMux I__6227 (
            .O(N__33015),
            .I(N__33006));
    InMux I__6226 (
            .O(N__33012),
            .I(N__32997));
    InMux I__6225 (
            .O(N__33011),
            .I(N__32997));
    InMux I__6224 (
            .O(N__33010),
            .I(N__32997));
    InMux I__6223 (
            .O(N__33009),
            .I(N__32997));
    LocalMux I__6222 (
            .O(N__33006),
            .I(N__32994));
    LocalMux I__6221 (
            .O(N__32997),
            .I(\comm_spi.bit_cnt_0 ));
    Odrv4 I__6220 (
            .O(N__32994),
            .I(\comm_spi.bit_cnt_0 ));
    InMux I__6219 (
            .O(N__32989),
            .I(N__32984));
    InMux I__6218 (
            .O(N__32988),
            .I(N__32979));
    InMux I__6217 (
            .O(N__32987),
            .I(N__32979));
    LocalMux I__6216 (
            .O(N__32984),
            .I(N__32976));
    LocalMux I__6215 (
            .O(N__32979),
            .I(\comm_spi.bit_cnt_2 ));
    Odrv4 I__6214 (
            .O(N__32976),
            .I(\comm_spi.bit_cnt_2 ));
    CascadeMux I__6213 (
            .O(N__32971),
            .I(N__32968));
    InMux I__6212 (
            .O(N__32968),
            .I(N__32965));
    LocalMux I__6211 (
            .O(N__32965),
            .I(N__32962));
    Span4Mux_h I__6210 (
            .O(N__32962),
            .I(N__32959));
    Odrv4 I__6209 (
            .O(N__32959),
            .I(comm_buf_3_1));
    CascadeMux I__6208 (
            .O(N__32956),
            .I(n21991_cascade_));
    InMux I__6207 (
            .O(N__32953),
            .I(N__32948));
    InMux I__6206 (
            .O(N__32952),
            .I(N__32943));
    InMux I__6205 (
            .O(N__32951),
            .I(N__32943));
    LocalMux I__6204 (
            .O(N__32948),
            .I(\ADC_VDC.bit_cnt_6 ));
    LocalMux I__6203 (
            .O(N__32943),
            .I(\ADC_VDC.bit_cnt_6 ));
    InMux I__6202 (
            .O(N__32938),
            .I(\ADC_VDC.n19474 ));
    InMux I__6201 (
            .O(N__32935),
            .I(\ADC_VDC.n19475 ));
    InMux I__6200 (
            .O(N__32932),
            .I(N__32927));
    InMux I__6199 (
            .O(N__32931),
            .I(N__32924));
    InMux I__6198 (
            .O(N__32930),
            .I(N__32921));
    LocalMux I__6197 (
            .O(N__32927),
            .I(\ADC_VDC.bit_cnt_7 ));
    LocalMux I__6196 (
            .O(N__32924),
            .I(\ADC_VDC.bit_cnt_7 ));
    LocalMux I__6195 (
            .O(N__32921),
            .I(\ADC_VDC.bit_cnt_7 ));
    IoInMux I__6194 (
            .O(N__32914),
            .I(N__32909));
    ClkMux I__6193 (
            .O(N__32913),
            .I(N__32905));
    ClkMux I__6192 (
            .O(N__32912),
            .I(N__32900));
    LocalMux I__6191 (
            .O(N__32909),
            .I(N__32897));
    ClkMux I__6190 (
            .O(N__32908),
            .I(N__32890));
    LocalMux I__6189 (
            .O(N__32905),
            .I(N__32887));
    ClkMux I__6188 (
            .O(N__32904),
            .I(N__32881));
    ClkMux I__6187 (
            .O(N__32903),
            .I(N__32877));
    LocalMux I__6186 (
            .O(N__32900),
            .I(N__32874));
    IoSpan4Mux I__6185 (
            .O(N__32897),
            .I(N__32868));
    ClkMux I__6184 (
            .O(N__32896),
            .I(N__32865));
    ClkMux I__6183 (
            .O(N__32895),
            .I(N__32862));
    ClkMux I__6182 (
            .O(N__32894),
            .I(N__32858));
    ClkMux I__6181 (
            .O(N__32893),
            .I(N__32855));
    LocalMux I__6180 (
            .O(N__32890),
            .I(N__32850));
    Span4Mux_h I__6179 (
            .O(N__32887),
            .I(N__32850));
    ClkMux I__6178 (
            .O(N__32886),
            .I(N__32847));
    ClkMux I__6177 (
            .O(N__32885),
            .I(N__32843));
    ClkMux I__6176 (
            .O(N__32884),
            .I(N__32839));
    LocalMux I__6175 (
            .O(N__32881),
            .I(N__32836));
    ClkMux I__6174 (
            .O(N__32880),
            .I(N__32833));
    LocalMux I__6173 (
            .O(N__32877),
            .I(N__32830));
    Span4Mux_h I__6172 (
            .O(N__32874),
            .I(N__32827));
    ClkMux I__6171 (
            .O(N__32873),
            .I(N__32824));
    ClkMux I__6170 (
            .O(N__32872),
            .I(N__32821));
    ClkMux I__6169 (
            .O(N__32871),
            .I(N__32818));
    Span4Mux_s3_h I__6168 (
            .O(N__32868),
            .I(N__32815));
    LocalMux I__6167 (
            .O(N__32865),
            .I(N__32810));
    LocalMux I__6166 (
            .O(N__32862),
            .I(N__32810));
    ClkMux I__6165 (
            .O(N__32861),
            .I(N__32807));
    LocalMux I__6164 (
            .O(N__32858),
            .I(N__32801));
    LocalMux I__6163 (
            .O(N__32855),
            .I(N__32801));
    Span4Mux_h I__6162 (
            .O(N__32850),
            .I(N__32796));
    LocalMux I__6161 (
            .O(N__32847),
            .I(N__32796));
    ClkMux I__6160 (
            .O(N__32846),
            .I(N__32793));
    LocalMux I__6159 (
            .O(N__32843),
            .I(N__32790));
    ClkMux I__6158 (
            .O(N__32842),
            .I(N__32787));
    LocalMux I__6157 (
            .O(N__32839),
            .I(N__32784));
    Span4Mux_h I__6156 (
            .O(N__32836),
            .I(N__32779));
    LocalMux I__6155 (
            .O(N__32833),
            .I(N__32779));
    Span4Mux_h I__6154 (
            .O(N__32830),
            .I(N__32775));
    Span4Mux_v I__6153 (
            .O(N__32827),
            .I(N__32770));
    LocalMux I__6152 (
            .O(N__32824),
            .I(N__32770));
    LocalMux I__6151 (
            .O(N__32821),
            .I(N__32765));
    LocalMux I__6150 (
            .O(N__32818),
            .I(N__32765));
    Span4Mux_h I__6149 (
            .O(N__32815),
            .I(N__32762));
    Span4Mux_h I__6148 (
            .O(N__32810),
            .I(N__32757));
    LocalMux I__6147 (
            .O(N__32807),
            .I(N__32757));
    ClkMux I__6146 (
            .O(N__32806),
            .I(N__32754));
    Span4Mux_h I__6145 (
            .O(N__32801),
            .I(N__32751));
    Span4Mux_v I__6144 (
            .O(N__32796),
            .I(N__32746));
    LocalMux I__6143 (
            .O(N__32793),
            .I(N__32746));
    Span4Mux_v I__6142 (
            .O(N__32790),
            .I(N__32741));
    LocalMux I__6141 (
            .O(N__32787),
            .I(N__32741));
    Span4Mux_h I__6140 (
            .O(N__32784),
            .I(N__32736));
    Span4Mux_h I__6139 (
            .O(N__32779),
            .I(N__32736));
    ClkMux I__6138 (
            .O(N__32778),
            .I(N__32733));
    Span4Mux_v I__6137 (
            .O(N__32775),
            .I(N__32728));
    Span4Mux_h I__6136 (
            .O(N__32770),
            .I(N__32728));
    Span4Mux_h I__6135 (
            .O(N__32765),
            .I(N__32724));
    Span4Mux_h I__6134 (
            .O(N__32762),
            .I(N__32719));
    Span4Mux_v I__6133 (
            .O(N__32757),
            .I(N__32719));
    LocalMux I__6132 (
            .O(N__32754),
            .I(N__32716));
    Span4Mux_v I__6131 (
            .O(N__32751),
            .I(N__32711));
    Span4Mux_h I__6130 (
            .O(N__32746),
            .I(N__32711));
    Span4Mux_h I__6129 (
            .O(N__32741),
            .I(N__32704));
    Span4Mux_v I__6128 (
            .O(N__32736),
            .I(N__32704));
    LocalMux I__6127 (
            .O(N__32733),
            .I(N__32704));
    Span4Mux_v I__6126 (
            .O(N__32728),
            .I(N__32701));
    ClkMux I__6125 (
            .O(N__32727),
            .I(N__32698));
    Span4Mux_v I__6124 (
            .O(N__32724),
            .I(N__32693));
    Span4Mux_h I__6123 (
            .O(N__32719),
            .I(N__32693));
    Span4Mux_h I__6122 (
            .O(N__32716),
            .I(N__32688));
    Span4Mux_v I__6121 (
            .O(N__32711),
            .I(N__32688));
    Sp12to4 I__6120 (
            .O(N__32704),
            .I(N__32685));
    Span4Mux_h I__6119 (
            .O(N__32701),
            .I(N__32680));
    LocalMux I__6118 (
            .O(N__32698),
            .I(N__32680));
    Odrv4 I__6117 (
            .O(N__32693),
            .I(VDC_CLK));
    Odrv4 I__6116 (
            .O(N__32688),
            .I(VDC_CLK));
    Odrv12 I__6115 (
            .O(N__32685),
            .I(VDC_CLK));
    Odrv4 I__6114 (
            .O(N__32680),
            .I(VDC_CLK));
    SRMux I__6113 (
            .O(N__32671),
            .I(N__32668));
    LocalMux I__6112 (
            .O(N__32668),
            .I(N__32665));
    Span4Mux_h I__6111 (
            .O(N__32665),
            .I(N__32662));
    Odrv4 I__6110 (
            .O(N__32662),
            .I(\ADC_VDC.n18381 ));
    InMux I__6109 (
            .O(N__32659),
            .I(N__32656));
    LocalMux I__6108 (
            .O(N__32656),
            .I(N__32653));
    Span4Mux_v I__6107 (
            .O(N__32653),
            .I(N__32650));
    Span4Mux_h I__6106 (
            .O(N__32650),
            .I(N__32647));
    Span4Mux_h I__6105 (
            .O(N__32647),
            .I(N__32644));
    Odrv4 I__6104 (
            .O(N__32644),
            .I(buf_data_iac_6));
    InMux I__6103 (
            .O(N__32641),
            .I(N__32637));
    CascadeMux I__6102 (
            .O(N__32640),
            .I(N__32634));
    LocalMux I__6101 (
            .O(N__32637),
            .I(N__32629));
    InMux I__6100 (
            .O(N__32634),
            .I(N__32626));
    InMux I__6099 (
            .O(N__32633),
            .I(N__32622));
    InMux I__6098 (
            .O(N__32632),
            .I(N__32619));
    Span4Mux_v I__6097 (
            .O(N__32629),
            .I(N__32616));
    LocalMux I__6096 (
            .O(N__32626),
            .I(N__32613));
    InMux I__6095 (
            .O(N__32625),
            .I(N__32610));
    LocalMux I__6094 (
            .O(N__32622),
            .I(\ADC_VDC.bit_cnt_3 ));
    LocalMux I__6093 (
            .O(N__32619),
            .I(\ADC_VDC.bit_cnt_3 ));
    Odrv4 I__6092 (
            .O(N__32616),
            .I(\ADC_VDC.bit_cnt_3 ));
    Odrv4 I__6091 (
            .O(N__32613),
            .I(\ADC_VDC.bit_cnt_3 ));
    LocalMux I__6090 (
            .O(N__32610),
            .I(\ADC_VDC.bit_cnt_3 ));
    InMux I__6089 (
            .O(N__32599),
            .I(N__32596));
    LocalMux I__6088 (
            .O(N__32596),
            .I(N__32592));
    InMux I__6087 (
            .O(N__32595),
            .I(N__32586));
    Span4Mux_v I__6086 (
            .O(N__32592),
            .I(N__32583));
    InMux I__6085 (
            .O(N__32591),
            .I(N__32580));
    InMux I__6084 (
            .O(N__32590),
            .I(N__32575));
    InMux I__6083 (
            .O(N__32589),
            .I(N__32575));
    LocalMux I__6082 (
            .O(N__32586),
            .I(\ADC_VDC.bit_cnt_2 ));
    Odrv4 I__6081 (
            .O(N__32583),
            .I(\ADC_VDC.bit_cnt_2 ));
    LocalMux I__6080 (
            .O(N__32580),
            .I(\ADC_VDC.bit_cnt_2 ));
    LocalMux I__6079 (
            .O(N__32575),
            .I(\ADC_VDC.bit_cnt_2 ));
    InMux I__6078 (
            .O(N__32566),
            .I(N__32563));
    LocalMux I__6077 (
            .O(N__32563),
            .I(\ADC_VDC.n6_adj_1404 ));
    CascadeMux I__6076 (
            .O(N__32560),
            .I(\ADC_VDC.n11_cascade_ ));
    InMux I__6075 (
            .O(N__32557),
            .I(N__32554));
    LocalMux I__6074 (
            .O(N__32554),
            .I(\ADC_VDC.n17359 ));
    InMux I__6073 (
            .O(N__32551),
            .I(N__32548));
    LocalMux I__6072 (
            .O(N__32548),
            .I(N__32543));
    InMux I__6071 (
            .O(N__32547),
            .I(N__32538));
    InMux I__6070 (
            .O(N__32546),
            .I(N__32535));
    Span4Mux_h I__6069 (
            .O(N__32543),
            .I(N__32532));
    InMux I__6068 (
            .O(N__32542),
            .I(N__32527));
    InMux I__6067 (
            .O(N__32541),
            .I(N__32527));
    LocalMux I__6066 (
            .O(N__32538),
            .I(\ADC_VDC.bit_cnt_0 ));
    LocalMux I__6065 (
            .O(N__32535),
            .I(\ADC_VDC.bit_cnt_0 ));
    Odrv4 I__6064 (
            .O(N__32532),
            .I(\ADC_VDC.bit_cnt_0 ));
    LocalMux I__6063 (
            .O(N__32527),
            .I(\ADC_VDC.bit_cnt_0 ));
    InMux I__6062 (
            .O(N__32518),
            .I(bfn_13_6_0_));
    InMux I__6061 (
            .O(N__32515),
            .I(N__32512));
    LocalMux I__6060 (
            .O(N__32512),
            .I(N__32506));
    CascadeMux I__6059 (
            .O(N__32511),
            .I(N__32502));
    InMux I__6058 (
            .O(N__32510),
            .I(N__32499));
    InMux I__6057 (
            .O(N__32509),
            .I(N__32496));
    Span4Mux_h I__6056 (
            .O(N__32506),
            .I(N__32493));
    InMux I__6055 (
            .O(N__32505),
            .I(N__32488));
    InMux I__6054 (
            .O(N__32502),
            .I(N__32488));
    LocalMux I__6053 (
            .O(N__32499),
            .I(\ADC_VDC.bit_cnt_1 ));
    LocalMux I__6052 (
            .O(N__32496),
            .I(\ADC_VDC.bit_cnt_1 ));
    Odrv4 I__6051 (
            .O(N__32493),
            .I(\ADC_VDC.bit_cnt_1 ));
    LocalMux I__6050 (
            .O(N__32488),
            .I(\ADC_VDC.bit_cnt_1 ));
    InMux I__6049 (
            .O(N__32479),
            .I(\ADC_VDC.n19469 ));
    InMux I__6048 (
            .O(N__32476),
            .I(\ADC_VDC.n19470 ));
    InMux I__6047 (
            .O(N__32473),
            .I(\ADC_VDC.n19471 ));
    InMux I__6046 (
            .O(N__32470),
            .I(N__32467));
    LocalMux I__6045 (
            .O(N__32467),
            .I(N__32460));
    InMux I__6044 (
            .O(N__32466),
            .I(N__32457));
    InMux I__6043 (
            .O(N__32465),
            .I(N__32450));
    InMux I__6042 (
            .O(N__32464),
            .I(N__32450));
    InMux I__6041 (
            .O(N__32463),
            .I(N__32450));
    Span4Mux_h I__6040 (
            .O(N__32460),
            .I(N__32447));
    LocalMux I__6039 (
            .O(N__32457),
            .I(\ADC_VDC.bit_cnt_4 ));
    LocalMux I__6038 (
            .O(N__32450),
            .I(\ADC_VDC.bit_cnt_4 ));
    Odrv4 I__6037 (
            .O(N__32447),
            .I(\ADC_VDC.bit_cnt_4 ));
    InMux I__6036 (
            .O(N__32440),
            .I(\ADC_VDC.n19472 ));
    InMux I__6035 (
            .O(N__32437),
            .I(N__32432));
    InMux I__6034 (
            .O(N__32436),
            .I(N__32429));
    InMux I__6033 (
            .O(N__32435),
            .I(N__32426));
    LocalMux I__6032 (
            .O(N__32432),
            .I(\ADC_VDC.bit_cnt_5 ));
    LocalMux I__6031 (
            .O(N__32429),
            .I(\ADC_VDC.bit_cnt_5 ));
    LocalMux I__6030 (
            .O(N__32426),
            .I(\ADC_VDC.bit_cnt_5 ));
    InMux I__6029 (
            .O(N__32419),
            .I(\ADC_VDC.n19473 ));
    CascadeMux I__6028 (
            .O(N__32416),
            .I(\comm_spi.n22632_cascade_ ));
    CascadeMux I__6027 (
            .O(N__32413),
            .I(\comm_spi.imosi_cascade_ ));
    InMux I__6026 (
            .O(N__32410),
            .I(N__32404));
    InMux I__6025 (
            .O(N__32409),
            .I(N__32404));
    LocalMux I__6024 (
            .O(N__32404),
            .I(\comm_spi.imosi ));
    InMux I__6023 (
            .O(N__32401),
            .I(N__32398));
    LocalMux I__6022 (
            .O(N__32398),
            .I(\comm_spi.n14599 ));
    SRMux I__6021 (
            .O(N__32395),
            .I(N__32392));
    LocalMux I__6020 (
            .O(N__32392),
            .I(N__32389));
    Span4Mux_h I__6019 (
            .O(N__32389),
            .I(N__32386));
    Odrv4 I__6018 (
            .O(N__32386),
            .I(\comm_spi.DOUT_7__N_738 ));
    InMux I__6017 (
            .O(N__32383),
            .I(N__32379));
    InMux I__6016 (
            .O(N__32382),
            .I(N__32376));
    LocalMux I__6015 (
            .O(N__32379),
            .I(\ADC_VDC.genclk.n21167 ));
    LocalMux I__6014 (
            .O(N__32376),
            .I(\ADC_VDC.genclk.n21167 ));
    InMux I__6013 (
            .O(N__32371),
            .I(N__32367));
    CascadeMux I__6012 (
            .O(N__32370),
            .I(N__32363));
    LocalMux I__6011 (
            .O(N__32367),
            .I(N__32360));
    InMux I__6010 (
            .O(N__32366),
            .I(N__32355));
    InMux I__6009 (
            .O(N__32363),
            .I(N__32355));
    Odrv4 I__6008 (
            .O(N__32360),
            .I(buf_dds0_10));
    LocalMux I__6007 (
            .O(N__32355),
            .I(buf_dds0_10));
    InMux I__6006 (
            .O(N__32350),
            .I(N__32347));
    LocalMux I__6005 (
            .O(N__32347),
            .I(\SIG_DDS.tmp_buf_10 ));
    InMux I__6004 (
            .O(N__32344),
            .I(N__32341));
    LocalMux I__6003 (
            .O(N__32341),
            .I(N__32338));
    Span4Mux_h I__6002 (
            .O(N__32338),
            .I(N__32333));
    InMux I__6001 (
            .O(N__32337),
            .I(N__32330));
    InMux I__6000 (
            .O(N__32336),
            .I(N__32327));
    Odrv4 I__5999 (
            .O(N__32333),
            .I(buf_dds0_9));
    LocalMux I__5998 (
            .O(N__32330),
            .I(buf_dds0_9));
    LocalMux I__5997 (
            .O(N__32327),
            .I(buf_dds0_9));
    CascadeMux I__5996 (
            .O(N__32320),
            .I(N__32317));
    InMux I__5995 (
            .O(N__32317),
            .I(N__32314));
    LocalMux I__5994 (
            .O(N__32314),
            .I(\SIG_DDS.tmp_buf_9 ));
    InMux I__5993 (
            .O(N__32311),
            .I(N__32307));
    InMux I__5992 (
            .O(N__32310),
            .I(N__32304));
    LocalMux I__5991 (
            .O(N__32307),
            .I(N__32301));
    LocalMux I__5990 (
            .O(N__32304),
            .I(N__32297));
    Span4Mux_h I__5989 (
            .O(N__32301),
            .I(N__32294));
    InMux I__5988 (
            .O(N__32300),
            .I(N__32291));
    Span4Mux_v I__5987 (
            .O(N__32297),
            .I(N__32288));
    Odrv4 I__5986 (
            .O(N__32294),
            .I(buf_dds0_13));
    LocalMux I__5985 (
            .O(N__32291),
            .I(buf_dds0_13));
    Odrv4 I__5984 (
            .O(N__32288),
            .I(buf_dds0_13));
    CascadeMux I__5983 (
            .O(N__32281),
            .I(N__32278));
    InMux I__5982 (
            .O(N__32278),
            .I(N__32275));
    LocalMux I__5981 (
            .O(N__32275),
            .I(\SIG_DDS.tmp_buf_13 ));
    CascadeMux I__5980 (
            .O(N__32272),
            .I(N__32268));
    InMux I__5979 (
            .O(N__32271),
            .I(N__32265));
    InMux I__5978 (
            .O(N__32268),
            .I(N__32262));
    LocalMux I__5977 (
            .O(N__32265),
            .I(N__32259));
    LocalMux I__5976 (
            .O(N__32262),
            .I(N__32255));
    Span4Mux_v I__5975 (
            .O(N__32259),
            .I(N__32252));
    InMux I__5974 (
            .O(N__32258),
            .I(N__32249));
    Span4Mux_h I__5973 (
            .O(N__32255),
            .I(N__32246));
    Odrv4 I__5972 (
            .O(N__32252),
            .I(buf_dds0_14));
    LocalMux I__5971 (
            .O(N__32249),
            .I(buf_dds0_14));
    Odrv4 I__5970 (
            .O(N__32246),
            .I(buf_dds0_14));
    InMux I__5969 (
            .O(N__32239),
            .I(N__32235));
    InMux I__5968 (
            .O(N__32238),
            .I(N__32232));
    LocalMux I__5967 (
            .O(N__32235),
            .I(N__32228));
    LocalMux I__5966 (
            .O(N__32232),
            .I(N__32225));
    InMux I__5965 (
            .O(N__32231),
            .I(N__32222));
    Span4Mux_v I__5964 (
            .O(N__32228),
            .I(N__32219));
    Odrv4 I__5963 (
            .O(N__32225),
            .I(buf_dds0_1));
    LocalMux I__5962 (
            .O(N__32222),
            .I(buf_dds0_1));
    Odrv4 I__5961 (
            .O(N__32219),
            .I(buf_dds0_1));
    CascadeMux I__5960 (
            .O(N__32212),
            .I(N__32209));
    InMux I__5959 (
            .O(N__32209),
            .I(N__32206));
    LocalMux I__5958 (
            .O(N__32206),
            .I(\SIG_DDS.tmp_buf_7 ));
    CascadeMux I__5957 (
            .O(N__32203),
            .I(N__32200));
    InMux I__5956 (
            .O(N__32200),
            .I(N__32197));
    LocalMux I__5955 (
            .O(N__32197),
            .I(\SIG_DDS.tmp_buf_8 ));
    InMux I__5954 (
            .O(N__32194),
            .I(N__32191));
    LocalMux I__5953 (
            .O(N__32191),
            .I(\comm_spi.n22629 ));
    CascadeMux I__5952 (
            .O(N__32188),
            .I(\comm_spi.n22629_cascade_ ));
    CascadeMux I__5951 (
            .O(N__32185),
            .I(N__32182));
    InMux I__5950 (
            .O(N__32182),
            .I(N__32173));
    InMux I__5949 (
            .O(N__32181),
            .I(N__32173));
    InMux I__5948 (
            .O(N__32180),
            .I(N__32170));
    InMux I__5947 (
            .O(N__32179),
            .I(N__32165));
    InMux I__5946 (
            .O(N__32178),
            .I(N__32165));
    LocalMux I__5945 (
            .O(N__32173),
            .I(N__32152));
    LocalMux I__5944 (
            .O(N__32170),
            .I(N__32147));
    LocalMux I__5943 (
            .O(N__32165),
            .I(N__32147));
    InMux I__5942 (
            .O(N__32164),
            .I(N__32138));
    InMux I__5941 (
            .O(N__32163),
            .I(N__32138));
    InMux I__5940 (
            .O(N__32162),
            .I(N__32138));
    InMux I__5939 (
            .O(N__32161),
            .I(N__32138));
    InMux I__5938 (
            .O(N__32160),
            .I(N__32131));
    InMux I__5937 (
            .O(N__32159),
            .I(N__32131));
    InMux I__5936 (
            .O(N__32158),
            .I(N__32131));
    InMux I__5935 (
            .O(N__32157),
            .I(N__32128));
    InMux I__5934 (
            .O(N__32156),
            .I(N__32125));
    InMux I__5933 (
            .O(N__32155),
            .I(N__32122));
    Span4Mux_v I__5932 (
            .O(N__32152),
            .I(N__32117));
    Span4Mux_v I__5931 (
            .O(N__32147),
            .I(N__32117));
    LocalMux I__5930 (
            .O(N__32138),
            .I(N__32108));
    LocalMux I__5929 (
            .O(N__32131),
            .I(N__32108));
    LocalMux I__5928 (
            .O(N__32128),
            .I(N__32108));
    LocalMux I__5927 (
            .O(N__32125),
            .I(N__32108));
    LocalMux I__5926 (
            .O(N__32122),
            .I(eis_end_N_716));
    Odrv4 I__5925 (
            .O(N__32117),
            .I(eis_end_N_716));
    Odrv12 I__5924 (
            .O(N__32108),
            .I(eis_end_N_716));
    InMux I__5923 (
            .O(N__32101),
            .I(N__32096));
    InMux I__5922 (
            .O(N__32100),
            .I(N__32091));
    SRMux I__5921 (
            .O(N__32099),
            .I(N__32088));
    LocalMux I__5920 (
            .O(N__32096),
            .I(N__32084));
    InMux I__5919 (
            .O(N__32095),
            .I(N__32079));
    InMux I__5918 (
            .O(N__32094),
            .I(N__32079));
    LocalMux I__5917 (
            .O(N__32091),
            .I(N__32074));
    LocalMux I__5916 (
            .O(N__32088),
            .I(N__32074));
    CascadeMux I__5915 (
            .O(N__32087),
            .I(N__32071));
    Span4Mux_h I__5914 (
            .O(N__32084),
            .I(N__32064));
    LocalMux I__5913 (
            .O(N__32079),
            .I(N__32061));
    Sp12to4 I__5912 (
            .O(N__32074),
            .I(N__32058));
    InMux I__5911 (
            .O(N__32071),
            .I(N__32055));
    InMux I__5910 (
            .O(N__32070),
            .I(N__32052));
    InMux I__5909 (
            .O(N__32069),
            .I(N__32045));
    InMux I__5908 (
            .O(N__32068),
            .I(N__32045));
    InMux I__5907 (
            .O(N__32067),
            .I(N__32045));
    Odrv4 I__5906 (
            .O(N__32064),
            .I(acadc_rst));
    Odrv4 I__5905 (
            .O(N__32061),
            .I(acadc_rst));
    Odrv12 I__5904 (
            .O(N__32058),
            .I(acadc_rst));
    LocalMux I__5903 (
            .O(N__32055),
            .I(acadc_rst));
    LocalMux I__5902 (
            .O(N__32052),
            .I(acadc_rst));
    LocalMux I__5901 (
            .O(N__32045),
            .I(acadc_rst));
    InMux I__5900 (
            .O(N__32032),
            .I(N__32029));
    LocalMux I__5899 (
            .O(N__32029),
            .I(N__32026));
    Span4Mux_v I__5898 (
            .O(N__32026),
            .I(N__32023));
    Span4Mux_h I__5897 (
            .O(N__32023),
            .I(N__32020));
    Odrv4 I__5896 (
            .O(N__32020),
            .I(buf_data_iac_15));
    InMux I__5895 (
            .O(N__32017),
            .I(N__32013));
    InMux I__5894 (
            .O(N__32016),
            .I(N__32009));
    LocalMux I__5893 (
            .O(N__32013),
            .I(N__32006));
    InMux I__5892 (
            .O(N__32012),
            .I(N__32003));
    LocalMux I__5891 (
            .O(N__32009),
            .I(N__31998));
    Span4Mux_v I__5890 (
            .O(N__32006),
            .I(N__31998));
    LocalMux I__5889 (
            .O(N__32003),
            .I(N__31995));
    Odrv4 I__5888 (
            .O(N__31998),
            .I(buf_dds1_2));
    Odrv4 I__5887 (
            .O(N__31995),
            .I(buf_dds1_2));
    InMux I__5886 (
            .O(N__31990),
            .I(N__31987));
    LocalMux I__5885 (
            .O(N__31987),
            .I(N__31983));
    InMux I__5884 (
            .O(N__31986),
            .I(N__31980));
    Span4Mux_v I__5883 (
            .O(N__31983),
            .I(N__31976));
    LocalMux I__5882 (
            .O(N__31980),
            .I(N__31973));
    InMux I__5881 (
            .O(N__31979),
            .I(N__31970));
    Span4Mux_h I__5880 (
            .O(N__31976),
            .I(N__31965));
    Span4Mux_h I__5879 (
            .O(N__31973),
            .I(N__31965));
    LocalMux I__5878 (
            .O(N__31970),
            .I(buf_adcdata_iac_15));
    Odrv4 I__5877 (
            .O(N__31965),
            .I(buf_adcdata_iac_15));
    InMux I__5876 (
            .O(N__31960),
            .I(N__31957));
    LocalMux I__5875 (
            .O(N__31957),
            .I(N__31954));
    Span12Mux_v I__5874 (
            .O(N__31954),
            .I(N__31951));
    Odrv12 I__5873 (
            .O(N__31951),
            .I(n21961));
    CascadeMux I__5872 (
            .O(N__31948),
            .I(n16_adj_1621_cascade_));
    InMux I__5871 (
            .O(N__31945),
            .I(N__31942));
    LocalMux I__5870 (
            .O(N__31942),
            .I(N__31939));
    Span4Mux_v I__5869 (
            .O(N__31939),
            .I(N__31936));
    Odrv4 I__5868 (
            .O(N__31936),
            .I(n16_adj_1504));
    InMux I__5867 (
            .O(N__31933),
            .I(N__31928));
    InMux I__5866 (
            .O(N__31932),
            .I(N__31925));
    CascadeMux I__5865 (
            .O(N__31931),
            .I(N__31922));
    LocalMux I__5864 (
            .O(N__31928),
            .I(N__31917));
    LocalMux I__5863 (
            .O(N__31925),
            .I(N__31917));
    InMux I__5862 (
            .O(N__31922),
            .I(N__31914));
    Span4Mux_h I__5861 (
            .O(N__31917),
            .I(N__31911));
    LocalMux I__5860 (
            .O(N__31914),
            .I(buf_dds1_1));
    Odrv4 I__5859 (
            .O(N__31911),
            .I(buf_dds1_1));
    InMux I__5858 (
            .O(N__31906),
            .I(N__31899));
    InMux I__5857 (
            .O(N__31905),
            .I(N__31899));
    InMux I__5856 (
            .O(N__31904),
            .I(N__31896));
    LocalMux I__5855 (
            .O(N__31899),
            .I(acadc_skipCount_6));
    LocalMux I__5854 (
            .O(N__31896),
            .I(acadc_skipCount_6));
    InMux I__5853 (
            .O(N__31891),
            .I(N__31888));
    LocalMux I__5852 (
            .O(N__31888),
            .I(n17));
    InMux I__5851 (
            .O(N__31885),
            .I(N__31879));
    InMux I__5850 (
            .O(N__31884),
            .I(N__31876));
    InMux I__5849 (
            .O(N__31883),
            .I(N__31873));
    InMux I__5848 (
            .O(N__31882),
            .I(N__31870));
    LocalMux I__5847 (
            .O(N__31879),
            .I(acadc_dtrig_v));
    LocalMux I__5846 (
            .O(N__31876),
            .I(acadc_dtrig_v));
    LocalMux I__5845 (
            .O(N__31873),
            .I(acadc_dtrig_v));
    LocalMux I__5844 (
            .O(N__31870),
            .I(acadc_dtrig_v));
    InMux I__5843 (
            .O(N__31861),
            .I(N__31855));
    InMux I__5842 (
            .O(N__31860),
            .I(N__31852));
    InMux I__5841 (
            .O(N__31859),
            .I(N__31847));
    InMux I__5840 (
            .O(N__31858),
            .I(N__31847));
    LocalMux I__5839 (
            .O(N__31855),
            .I(acadc_dtrig_i));
    LocalMux I__5838 (
            .O(N__31852),
            .I(acadc_dtrig_i));
    LocalMux I__5837 (
            .O(N__31847),
            .I(acadc_dtrig_i));
    CascadeMux I__5836 (
            .O(N__31840),
            .I(iac_raw_buf_N_728_cascade_));
    InMux I__5835 (
            .O(N__31837),
            .I(N__31834));
    LocalMux I__5834 (
            .O(N__31834),
            .I(N__31831));
    Odrv4 I__5833 (
            .O(N__31831),
            .I(n21997));
    InMux I__5832 (
            .O(N__31828),
            .I(N__31824));
    InMux I__5831 (
            .O(N__31827),
            .I(N__31821));
    LocalMux I__5830 (
            .O(N__31824),
            .I(N__31815));
    LocalMux I__5829 (
            .O(N__31821),
            .I(N__31815));
    InMux I__5828 (
            .O(N__31820),
            .I(N__31812));
    Span4Mux_h I__5827 (
            .O(N__31815),
            .I(N__31809));
    LocalMux I__5826 (
            .O(N__31812),
            .I(buf_dds1_3));
    Odrv4 I__5825 (
            .O(N__31809),
            .I(buf_dds1_3));
    InMux I__5824 (
            .O(N__31804),
            .I(N__31801));
    LocalMux I__5823 (
            .O(N__31801),
            .I(N__31798));
    Span12Mux_h I__5822 (
            .O(N__31798),
            .I(N__31795));
    Odrv12 I__5821 (
            .O(N__31795),
            .I(n20624));
    CascadeMux I__5820 (
            .O(N__31792),
            .I(n12353_cascade_));
    CascadeMux I__5819 (
            .O(N__31789),
            .I(N__31786));
    InMux I__5818 (
            .O(N__31786),
            .I(N__31783));
    LocalMux I__5817 (
            .O(N__31783),
            .I(N__31780));
    Odrv4 I__5816 (
            .O(N__31780),
            .I(n35));
    SRMux I__5815 (
            .O(N__31777),
            .I(N__31773));
    SRMux I__5814 (
            .O(N__31776),
            .I(N__31770));
    LocalMux I__5813 (
            .O(N__31773),
            .I(N__31763));
    LocalMux I__5812 (
            .O(N__31770),
            .I(N__31760));
    SRMux I__5811 (
            .O(N__31769),
            .I(N__31757));
    SRMux I__5810 (
            .O(N__31768),
            .I(N__31754));
    SRMux I__5809 (
            .O(N__31767),
            .I(N__31747));
    SRMux I__5808 (
            .O(N__31766),
            .I(N__31744));
    Span4Mux_h I__5807 (
            .O(N__31763),
            .I(N__31741));
    Span4Mux_v I__5806 (
            .O(N__31760),
            .I(N__31736));
    LocalMux I__5805 (
            .O(N__31757),
            .I(N__31736));
    LocalMux I__5804 (
            .O(N__31754),
            .I(N__31733));
    SRMux I__5803 (
            .O(N__31753),
            .I(N__31730));
    SRMux I__5802 (
            .O(N__31752),
            .I(N__31727));
    SRMux I__5801 (
            .O(N__31751),
            .I(N__31723));
    SRMux I__5800 (
            .O(N__31750),
            .I(N__31720));
    LocalMux I__5799 (
            .O(N__31747),
            .I(N__31716));
    LocalMux I__5798 (
            .O(N__31744),
            .I(N__31713));
    Span4Mux_v I__5797 (
            .O(N__31741),
            .I(N__31708));
    Span4Mux_h I__5796 (
            .O(N__31736),
            .I(N__31708));
    Span4Mux_v I__5795 (
            .O(N__31733),
            .I(N__31703));
    LocalMux I__5794 (
            .O(N__31730),
            .I(N__31703));
    LocalMux I__5793 (
            .O(N__31727),
            .I(N__31700));
    SRMux I__5792 (
            .O(N__31726),
            .I(N__31697));
    LocalMux I__5791 (
            .O(N__31723),
            .I(N__31694));
    LocalMux I__5790 (
            .O(N__31720),
            .I(N__31691));
    SRMux I__5789 (
            .O(N__31719),
            .I(N__31688));
    Span4Mux_v I__5788 (
            .O(N__31716),
            .I(N__31685));
    Span4Mux_h I__5787 (
            .O(N__31713),
            .I(N__31682));
    Span4Mux_v I__5786 (
            .O(N__31708),
            .I(N__31677));
    Span4Mux_h I__5785 (
            .O(N__31703),
            .I(N__31677));
    Span4Mux_v I__5784 (
            .O(N__31700),
            .I(N__31672));
    LocalMux I__5783 (
            .O(N__31697),
            .I(N__31672));
    Span4Mux_v I__5782 (
            .O(N__31694),
            .I(N__31665));
    Span4Mux_v I__5781 (
            .O(N__31691),
            .I(N__31665));
    LocalMux I__5780 (
            .O(N__31688),
            .I(N__31665));
    Span4Mux_h I__5779 (
            .O(N__31685),
            .I(N__31662));
    Span4Mux_h I__5778 (
            .O(N__31682),
            .I(N__31659));
    Span4Mux_v I__5777 (
            .O(N__31677),
            .I(N__31654));
    Span4Mux_h I__5776 (
            .O(N__31672),
            .I(N__31654));
    Span4Mux_h I__5775 (
            .O(N__31665),
            .I(N__31651));
    Span4Mux_h I__5774 (
            .O(N__31662),
            .I(N__31648));
    Span4Mux_h I__5773 (
            .O(N__31659),
            .I(N__31641));
    Span4Mux_h I__5772 (
            .O(N__31654),
            .I(N__31641));
    Span4Mux_h I__5771 (
            .O(N__31651),
            .I(N__31641));
    Odrv4 I__5770 (
            .O(N__31648),
            .I(iac_raw_buf_N_726));
    Odrv4 I__5769 (
            .O(N__31641),
            .I(iac_raw_buf_N_726));
    CascadeMux I__5768 (
            .O(N__31636),
            .I(N__31633));
    CascadeBuf I__5767 (
            .O(N__31633),
            .I(N__31630));
    CascadeMux I__5766 (
            .O(N__31630),
            .I(N__31627));
    CascadeBuf I__5765 (
            .O(N__31627),
            .I(N__31624));
    CascadeMux I__5764 (
            .O(N__31624),
            .I(N__31621));
    CascadeBuf I__5763 (
            .O(N__31621),
            .I(N__31618));
    CascadeMux I__5762 (
            .O(N__31618),
            .I(N__31615));
    CascadeBuf I__5761 (
            .O(N__31615),
            .I(N__31612));
    CascadeMux I__5760 (
            .O(N__31612),
            .I(N__31609));
    CascadeBuf I__5759 (
            .O(N__31609),
            .I(N__31606));
    CascadeMux I__5758 (
            .O(N__31606),
            .I(N__31603));
    CascadeBuf I__5757 (
            .O(N__31603),
            .I(N__31600));
    CascadeMux I__5756 (
            .O(N__31600),
            .I(N__31597));
    CascadeBuf I__5755 (
            .O(N__31597),
            .I(N__31594));
    CascadeMux I__5754 (
            .O(N__31594),
            .I(N__31591));
    CascadeBuf I__5753 (
            .O(N__31591),
            .I(N__31588));
    CascadeMux I__5752 (
            .O(N__31588),
            .I(N__31584));
    CascadeMux I__5751 (
            .O(N__31587),
            .I(N__31581));
    CascadeBuf I__5750 (
            .O(N__31584),
            .I(N__31578));
    CascadeBuf I__5749 (
            .O(N__31581),
            .I(N__31575));
    CascadeMux I__5748 (
            .O(N__31578),
            .I(N__31572));
    CascadeMux I__5747 (
            .O(N__31575),
            .I(N__31569));
    InMux I__5746 (
            .O(N__31572),
            .I(N__31566));
    InMux I__5745 (
            .O(N__31569),
            .I(N__31563));
    LocalMux I__5744 (
            .O(N__31566),
            .I(N__31560));
    LocalMux I__5743 (
            .O(N__31563),
            .I(N__31557));
    Span4Mux_h I__5742 (
            .O(N__31560),
            .I(N__31554));
    Span4Mux_v I__5741 (
            .O(N__31557),
            .I(N__31551));
    Span4Mux_h I__5740 (
            .O(N__31554),
            .I(N__31548));
    Sp12to4 I__5739 (
            .O(N__31551),
            .I(N__31545));
    Span4Mux_v I__5738 (
            .O(N__31548),
            .I(N__31542));
    Odrv12 I__5737 (
            .O(N__31545),
            .I(data_index_9_N_212_0));
    Odrv4 I__5736 (
            .O(N__31542),
            .I(data_index_9_N_212_0));
    InMux I__5735 (
            .O(N__31537),
            .I(N__31534));
    LocalMux I__5734 (
            .O(N__31534),
            .I(N__31530));
    InMux I__5733 (
            .O(N__31533),
            .I(N__31526));
    Span4Mux_h I__5732 (
            .O(N__31530),
            .I(N__31523));
    InMux I__5731 (
            .O(N__31529),
            .I(N__31520));
    LocalMux I__5730 (
            .O(N__31526),
            .I(acadc_skipCount_8));
    Odrv4 I__5729 (
            .O(N__31523),
            .I(acadc_skipCount_8));
    LocalMux I__5728 (
            .O(N__31520),
            .I(acadc_skipCount_8));
    CascadeMux I__5727 (
            .O(N__31513),
            .I(n20_cascade_));
    InMux I__5726 (
            .O(N__31510),
            .I(N__31507));
    LocalMux I__5725 (
            .O(N__31507),
            .I(N__31504));
    Odrv4 I__5724 (
            .O(N__31504),
            .I(n14_adj_1498));
    InMux I__5723 (
            .O(N__31501),
            .I(N__31498));
    LocalMux I__5722 (
            .O(N__31498),
            .I(N__31495));
    Odrv4 I__5721 (
            .O(N__31495),
            .I(n18_adj_1587));
    CascadeMux I__5720 (
            .O(N__31492),
            .I(n26_adj_1604_cascade_));
    InMux I__5719 (
            .O(N__31489),
            .I(N__31483));
    InMux I__5718 (
            .O(N__31488),
            .I(N__31483));
    LocalMux I__5717 (
            .O(N__31483),
            .I(N__31480));
    Odrv4 I__5716 (
            .O(N__31480),
            .I(n31));
    CascadeMux I__5715 (
            .O(N__31477),
            .I(N__31474));
    CascadeBuf I__5714 (
            .O(N__31474),
            .I(N__31471));
    CascadeMux I__5713 (
            .O(N__31471),
            .I(N__31468));
    CascadeBuf I__5712 (
            .O(N__31468),
            .I(N__31465));
    CascadeMux I__5711 (
            .O(N__31465),
            .I(N__31462));
    CascadeBuf I__5710 (
            .O(N__31462),
            .I(N__31459));
    CascadeMux I__5709 (
            .O(N__31459),
            .I(N__31456));
    CascadeBuf I__5708 (
            .O(N__31456),
            .I(N__31453));
    CascadeMux I__5707 (
            .O(N__31453),
            .I(N__31450));
    CascadeBuf I__5706 (
            .O(N__31450),
            .I(N__31447));
    CascadeMux I__5705 (
            .O(N__31447),
            .I(N__31444));
    CascadeBuf I__5704 (
            .O(N__31444),
            .I(N__31441));
    CascadeMux I__5703 (
            .O(N__31441),
            .I(N__31438));
    CascadeBuf I__5702 (
            .O(N__31438),
            .I(N__31435));
    CascadeMux I__5701 (
            .O(N__31435),
            .I(N__31431));
    CascadeMux I__5700 (
            .O(N__31434),
            .I(N__31428));
    CascadeBuf I__5699 (
            .O(N__31431),
            .I(N__31425));
    CascadeBuf I__5698 (
            .O(N__31428),
            .I(N__31422));
    CascadeMux I__5697 (
            .O(N__31425),
            .I(N__31419));
    CascadeMux I__5696 (
            .O(N__31422),
            .I(N__31416));
    CascadeBuf I__5695 (
            .O(N__31419),
            .I(N__31413));
    InMux I__5694 (
            .O(N__31416),
            .I(N__31410));
    CascadeMux I__5693 (
            .O(N__31413),
            .I(N__31407));
    LocalMux I__5692 (
            .O(N__31410),
            .I(N__31404));
    InMux I__5691 (
            .O(N__31407),
            .I(N__31401));
    Span4Mux_v I__5690 (
            .O(N__31404),
            .I(N__31398));
    LocalMux I__5689 (
            .O(N__31401),
            .I(N__31395));
    Span4Mux_h I__5688 (
            .O(N__31398),
            .I(N__31392));
    Span4Mux_v I__5687 (
            .O(N__31395),
            .I(N__31389));
    Span4Mux_h I__5686 (
            .O(N__31392),
            .I(N__31384));
    Span4Mux_h I__5685 (
            .O(N__31389),
            .I(N__31384));
    Odrv4 I__5684 (
            .O(N__31384),
            .I(data_index_9_N_212_3));
    CascadeMux I__5683 (
            .O(N__31381),
            .I(N__31378));
    InMux I__5682 (
            .O(N__31378),
            .I(N__31373));
    InMux I__5681 (
            .O(N__31377),
            .I(N__31370));
    InMux I__5680 (
            .O(N__31376),
            .I(N__31367));
    LocalMux I__5679 (
            .O(N__31373),
            .I(N__31364));
    LocalMux I__5678 (
            .O(N__31370),
            .I(acadc_skipCount_5));
    LocalMux I__5677 (
            .O(N__31367),
            .I(acadc_skipCount_5));
    Odrv4 I__5676 (
            .O(N__31364),
            .I(acadc_skipCount_5));
    InMux I__5675 (
            .O(N__31357),
            .I(N__31353));
    InMux I__5674 (
            .O(N__31356),
            .I(N__31350));
    LocalMux I__5673 (
            .O(N__31353),
            .I(N__31347));
    LocalMux I__5672 (
            .O(N__31350),
            .I(data_idxvec_13));
    Odrv4 I__5671 (
            .O(N__31347),
            .I(data_idxvec_13));
    InMux I__5670 (
            .O(N__31342),
            .I(n19347));
    CascadeMux I__5669 (
            .O(N__31339),
            .I(N__31336));
    InMux I__5668 (
            .O(N__31336),
            .I(N__31333));
    LocalMux I__5667 (
            .O(N__31333),
            .I(N__31329));
    CascadeMux I__5666 (
            .O(N__31332),
            .I(N__31326));
    Span4Mux_h I__5665 (
            .O(N__31329),
            .I(N__31323));
    InMux I__5664 (
            .O(N__31326),
            .I(N__31320));
    Span4Mux_v I__5663 (
            .O(N__31323),
            .I(N__31317));
    LocalMux I__5662 (
            .O(N__31320),
            .I(data_idxvec_14));
    Odrv4 I__5661 (
            .O(N__31317),
            .I(data_idxvec_14));
    InMux I__5660 (
            .O(N__31312),
            .I(n19348));
    InMux I__5659 (
            .O(N__31309),
            .I(n19349));
    InMux I__5658 (
            .O(N__31306),
            .I(N__31303));
    LocalMux I__5657 (
            .O(N__31303),
            .I(N__31299));
    InMux I__5656 (
            .O(N__31302),
            .I(N__31296));
    Span4Mux_h I__5655 (
            .O(N__31299),
            .I(N__31293));
    LocalMux I__5654 (
            .O(N__31296),
            .I(data_idxvec_15));
    Odrv4 I__5653 (
            .O(N__31293),
            .I(data_idxvec_15));
    InMux I__5652 (
            .O(N__31288),
            .I(N__31284));
    InMux I__5651 (
            .O(N__31287),
            .I(N__31281));
    LocalMux I__5650 (
            .O(N__31284),
            .I(N__31278));
    LocalMux I__5649 (
            .O(N__31281),
            .I(data_idxvec_5));
    Odrv4 I__5648 (
            .O(N__31278),
            .I(data_idxvec_5));
    CascadeMux I__5647 (
            .O(N__31273),
            .I(n26_adj_1486_cascade_));
    CascadeMux I__5646 (
            .O(N__31270),
            .I(n22177_cascade_));
    InMux I__5645 (
            .O(N__31267),
            .I(N__31264));
    LocalMux I__5644 (
            .O(N__31264),
            .I(N__31261));
    Span4Mux_v I__5643 (
            .O(N__31261),
            .I(N__31258));
    Odrv4 I__5642 (
            .O(N__31258),
            .I(n22120));
    CascadeMux I__5641 (
            .O(N__31255),
            .I(n22180_cascade_));
    CascadeMux I__5640 (
            .O(N__31252),
            .I(n30_adj_1485_cascade_));
    InMux I__5639 (
            .O(N__31249),
            .I(N__31246));
    LocalMux I__5638 (
            .O(N__31246),
            .I(N__31243));
    Span4Mux_h I__5637 (
            .O(N__31243),
            .I(N__31240));
    Span4Mux_h I__5636 (
            .O(N__31240),
            .I(N__31237));
    Odrv4 I__5635 (
            .O(N__31237),
            .I(buf_data_iac_13));
    InMux I__5634 (
            .O(N__31234),
            .I(N__31231));
    LocalMux I__5633 (
            .O(N__31231),
            .I(n21036));
    InMux I__5632 (
            .O(N__31228),
            .I(n19338));
    InMux I__5631 (
            .O(N__31225),
            .I(n19339));
    InMux I__5630 (
            .O(N__31222),
            .I(N__31218));
    InMux I__5629 (
            .O(N__31221),
            .I(N__31215));
    LocalMux I__5628 (
            .O(N__31218),
            .I(N__31212));
    LocalMux I__5627 (
            .O(N__31215),
            .I(data_idxvec_6));
    Odrv4 I__5626 (
            .O(N__31212),
            .I(data_idxvec_6));
    InMux I__5625 (
            .O(N__31207),
            .I(n19340));
    InMux I__5624 (
            .O(N__31204),
            .I(n19341));
    InMux I__5623 (
            .O(N__31201),
            .I(bfn_12_13_0_));
    InMux I__5622 (
            .O(N__31198),
            .I(N__31195));
    LocalMux I__5621 (
            .O(N__31195),
            .I(N__31191));
    InMux I__5620 (
            .O(N__31194),
            .I(N__31188));
    Span4Mux_v I__5619 (
            .O(N__31191),
            .I(N__31185));
    LocalMux I__5618 (
            .O(N__31188),
            .I(data_idxvec_9));
    Odrv4 I__5617 (
            .O(N__31185),
            .I(data_idxvec_9));
    InMux I__5616 (
            .O(N__31180),
            .I(n19343));
    CascadeMux I__5615 (
            .O(N__31177),
            .I(N__31173));
    InMux I__5614 (
            .O(N__31176),
            .I(N__31170));
    InMux I__5613 (
            .O(N__31173),
            .I(N__31167));
    LocalMux I__5612 (
            .O(N__31170),
            .I(N__31164));
    LocalMux I__5611 (
            .O(N__31167),
            .I(N__31159));
    Span4Mux_v I__5610 (
            .O(N__31164),
            .I(N__31159));
    Odrv4 I__5609 (
            .O(N__31159),
            .I(data_idxvec_10));
    InMux I__5608 (
            .O(N__31156),
            .I(n19344));
    InMux I__5607 (
            .O(N__31153),
            .I(n19345));
    CascadeMux I__5606 (
            .O(N__31150),
            .I(N__31147));
    InMux I__5605 (
            .O(N__31147),
            .I(N__31143));
    CascadeMux I__5604 (
            .O(N__31146),
            .I(N__31140));
    LocalMux I__5603 (
            .O(N__31143),
            .I(N__31137));
    InMux I__5602 (
            .O(N__31140),
            .I(N__31134));
    Span4Mux_h I__5601 (
            .O(N__31137),
            .I(N__31131));
    LocalMux I__5600 (
            .O(N__31134),
            .I(data_idxvec_12));
    Odrv4 I__5599 (
            .O(N__31131),
            .I(data_idxvec_12));
    InMux I__5598 (
            .O(N__31126),
            .I(n19346));
    InMux I__5597 (
            .O(N__31123),
            .I(N__31120));
    LocalMux I__5596 (
            .O(N__31120),
            .I(N__31117));
    Span4Mux_h I__5595 (
            .O(N__31117),
            .I(N__31114));
    Span4Mux_v I__5594 (
            .O(N__31114),
            .I(N__31111));
    Span4Mux_h I__5593 (
            .O(N__31111),
            .I(N__31108));
    Odrv4 I__5592 (
            .O(N__31108),
            .I(buf_data_vac_13));
    InMux I__5591 (
            .O(N__31105),
            .I(N__31102));
    LocalMux I__5590 (
            .O(N__31102),
            .I(N__31099));
    Span4Mux_h I__5589 (
            .O(N__31099),
            .I(N__31096));
    Span4Mux_v I__5588 (
            .O(N__31096),
            .I(N__31093));
    Span4Mux_h I__5587 (
            .O(N__31093),
            .I(N__31090));
    Odrv4 I__5586 (
            .O(N__31090),
            .I(buf_data_vac_12));
    InMux I__5585 (
            .O(N__31087),
            .I(N__31084));
    LocalMux I__5584 (
            .O(N__31084),
            .I(N__31081));
    Span4Mux_h I__5583 (
            .O(N__31081),
            .I(N__31078));
    Span4Mux_h I__5582 (
            .O(N__31078),
            .I(N__31075));
    Span4Mux_v I__5581 (
            .O(N__31075),
            .I(N__31072));
    Odrv4 I__5580 (
            .O(N__31072),
            .I(buf_data_vac_11));
    InMux I__5579 (
            .O(N__31069),
            .I(N__31066));
    LocalMux I__5578 (
            .O(N__31066),
            .I(N__31063));
    Span4Mux_v I__5577 (
            .O(N__31063),
            .I(N__31060));
    Span4Mux_v I__5576 (
            .O(N__31060),
            .I(N__31057));
    Span4Mux_h I__5575 (
            .O(N__31057),
            .I(N__31054));
    Span4Mux_h I__5574 (
            .O(N__31054),
            .I(N__31051));
    Odrv4 I__5573 (
            .O(N__31051),
            .I(buf_data_vac_10));
    InMux I__5572 (
            .O(N__31048),
            .I(N__31045));
    LocalMux I__5571 (
            .O(N__31045),
            .I(N__31042));
    Span4Mux_h I__5570 (
            .O(N__31042),
            .I(N__31039));
    Span4Mux_v I__5569 (
            .O(N__31039),
            .I(N__31036));
    Span4Mux_v I__5568 (
            .O(N__31036),
            .I(N__31033));
    Span4Mux_h I__5567 (
            .O(N__31033),
            .I(N__31030));
    Odrv4 I__5566 (
            .O(N__31030),
            .I(buf_data_vac_9));
    InMux I__5565 (
            .O(N__31027),
            .I(N__31024));
    LocalMux I__5564 (
            .O(N__31024),
            .I(N__31021));
    Span4Mux_h I__5563 (
            .O(N__31021),
            .I(N__31018));
    Span4Mux_h I__5562 (
            .O(N__31018),
            .I(N__31015));
    Odrv4 I__5561 (
            .O(N__31015),
            .I(n14_adj_1516));
    InMux I__5560 (
            .O(N__31012),
            .I(bfn_12_12_0_));
    InMux I__5559 (
            .O(N__31009),
            .I(n19335));
    InMux I__5558 (
            .O(N__31006),
            .I(n19336));
    InMux I__5557 (
            .O(N__31003),
            .I(n19337));
    InMux I__5556 (
            .O(N__31000),
            .I(N__30994));
    InMux I__5555 (
            .O(N__30999),
            .I(N__30994));
    LocalMux I__5554 (
            .O(N__30994),
            .I(N__30986));
    CascadeMux I__5553 (
            .O(N__30993),
            .I(N__30983));
    InMux I__5552 (
            .O(N__30992),
            .I(N__30980));
    InMux I__5551 (
            .O(N__30991),
            .I(N__30977));
    InMux I__5550 (
            .O(N__30990),
            .I(N__30972));
    InMux I__5549 (
            .O(N__30989),
            .I(N__30972));
    Sp12to4 I__5548 (
            .O(N__30986),
            .I(N__30969));
    InMux I__5547 (
            .O(N__30983),
            .I(N__30966));
    LocalMux I__5546 (
            .O(N__30980),
            .I(N__30959));
    LocalMux I__5545 (
            .O(N__30977),
            .I(N__30959));
    LocalMux I__5544 (
            .O(N__30972),
            .I(N__30959));
    Span12Mux_v I__5543 (
            .O(N__30969),
            .I(N__30956));
    LocalMux I__5542 (
            .O(N__30966),
            .I(N__30953));
    Span4Mux_h I__5541 (
            .O(N__30959),
            .I(N__30950));
    Odrv12 I__5540 (
            .O(N__30956),
            .I(n14490));
    Odrv4 I__5539 (
            .O(N__30953),
            .I(n14490));
    Odrv4 I__5538 (
            .O(N__30950),
            .I(n14490));
    InMux I__5537 (
            .O(N__30943),
            .I(N__30940));
    LocalMux I__5536 (
            .O(N__30940),
            .I(N__30936));
    InMux I__5535 (
            .O(N__30939),
            .I(N__30933));
    Span4Mux_h I__5534 (
            .O(N__30936),
            .I(N__30925));
    LocalMux I__5533 (
            .O(N__30933),
            .I(N__30922));
    InMux I__5532 (
            .O(N__30932),
            .I(N__30917));
    InMux I__5531 (
            .O(N__30931),
            .I(N__30917));
    InMux I__5530 (
            .O(N__30930),
            .I(N__30912));
    InMux I__5529 (
            .O(N__30929),
            .I(N__30912));
    InMux I__5528 (
            .O(N__30928),
            .I(N__30909));
    Odrv4 I__5527 (
            .O(N__30925),
            .I(n11882));
    Odrv4 I__5526 (
            .O(N__30922),
            .I(n11882));
    LocalMux I__5525 (
            .O(N__30917),
            .I(n11882));
    LocalMux I__5524 (
            .O(N__30912),
            .I(n11882));
    LocalMux I__5523 (
            .O(N__30909),
            .I(n11882));
    InMux I__5522 (
            .O(N__30898),
            .I(N__30895));
    LocalMux I__5521 (
            .O(N__30895),
            .I(N__30892));
    Span4Mux_v I__5520 (
            .O(N__30892),
            .I(N__30889));
    Span4Mux_h I__5519 (
            .O(N__30889),
            .I(N__30886));
    Odrv4 I__5518 (
            .O(N__30886),
            .I(buf_data_iac_0));
    InMux I__5517 (
            .O(N__30883),
            .I(N__30880));
    LocalMux I__5516 (
            .O(N__30880),
            .I(N__30877));
    Span4Mux_v I__5515 (
            .O(N__30877),
            .I(N__30874));
    Odrv4 I__5514 (
            .O(N__30874),
            .I(n22_adj_1476));
    InMux I__5513 (
            .O(N__30871),
            .I(N__30868));
    LocalMux I__5512 (
            .O(N__30868),
            .I(N__30865));
    Span4Mux_h I__5511 (
            .O(N__30865),
            .I(N__30862));
    Span4Mux_v I__5510 (
            .O(N__30862),
            .I(N__30859));
    Span4Mux_v I__5509 (
            .O(N__30859),
            .I(N__30856));
    Span4Mux_h I__5508 (
            .O(N__30856),
            .I(N__30853));
    Odrv4 I__5507 (
            .O(N__30853),
            .I(buf_data_vac_8));
    InMux I__5506 (
            .O(N__30850),
            .I(N__30847));
    LocalMux I__5505 (
            .O(N__30847),
            .I(N__30844));
    Span4Mux_h I__5504 (
            .O(N__30844),
            .I(N__30841));
    Span4Mux_h I__5503 (
            .O(N__30841),
            .I(N__30838));
    Span4Mux_h I__5502 (
            .O(N__30838),
            .I(N__30835));
    Odrv4 I__5501 (
            .O(N__30835),
            .I(buf_data_vac_15));
    InMux I__5500 (
            .O(N__30832),
            .I(N__30829));
    LocalMux I__5499 (
            .O(N__30829),
            .I(N__30826));
    Span4Mux_v I__5498 (
            .O(N__30826),
            .I(N__30823));
    Span4Mux_h I__5497 (
            .O(N__30823),
            .I(N__30820));
    Span4Mux_h I__5496 (
            .O(N__30820),
            .I(N__30817));
    Odrv4 I__5495 (
            .O(N__30817),
            .I(buf_data_vac_14));
    InMux I__5494 (
            .O(N__30814),
            .I(N__30811));
    LocalMux I__5493 (
            .O(N__30811),
            .I(N__30807));
    InMux I__5492 (
            .O(N__30810),
            .I(N__30804));
    Span4Mux_v I__5491 (
            .O(N__30807),
            .I(N__30800));
    LocalMux I__5490 (
            .O(N__30804),
            .I(N__30797));
    InMux I__5489 (
            .O(N__30803),
            .I(N__30794));
    Span4Mux_h I__5488 (
            .O(N__30800),
            .I(N__30791));
    Span4Mux_h I__5487 (
            .O(N__30797),
            .I(N__30788));
    LocalMux I__5486 (
            .O(N__30794),
            .I(N__30785));
    Odrv4 I__5485 (
            .O(N__30791),
            .I(comm_buf_0_7));
    Odrv4 I__5484 (
            .O(N__30788),
            .I(comm_buf_0_7));
    Odrv4 I__5483 (
            .O(N__30785),
            .I(comm_buf_0_7));
    InMux I__5482 (
            .O(N__30778),
            .I(N__30775));
    LocalMux I__5481 (
            .O(N__30775),
            .I(\ADC_VDC.n10 ));
    InMux I__5480 (
            .O(N__30772),
            .I(N__30767));
    InMux I__5479 (
            .O(N__30771),
            .I(N__30764));
    InMux I__5478 (
            .O(N__30770),
            .I(N__30761));
    LocalMux I__5477 (
            .O(N__30767),
            .I(\ADC_VDC.n15 ));
    LocalMux I__5476 (
            .O(N__30764),
            .I(\ADC_VDC.n15 ));
    LocalMux I__5475 (
            .O(N__30761),
            .I(\ADC_VDC.n15 ));
    InMux I__5474 (
            .O(N__30754),
            .I(N__30751));
    LocalMux I__5473 (
            .O(N__30751),
            .I(N__30748));
    Odrv4 I__5472 (
            .O(N__30748),
            .I(\ADC_VDC.n19_adj_1405 ));
    CascadeMux I__5471 (
            .O(N__30745),
            .I(N__30741));
    InMux I__5470 (
            .O(N__30744),
            .I(N__30736));
    InMux I__5469 (
            .O(N__30741),
            .I(N__30729));
    InMux I__5468 (
            .O(N__30740),
            .I(N__30729));
    InMux I__5467 (
            .O(N__30739),
            .I(N__30729));
    LocalMux I__5466 (
            .O(N__30736),
            .I(wdtick_cnt_0));
    LocalMux I__5465 (
            .O(N__30729),
            .I(wdtick_cnt_0));
    InMux I__5464 (
            .O(N__30724),
            .I(N__30718));
    InMux I__5463 (
            .O(N__30723),
            .I(N__30711));
    InMux I__5462 (
            .O(N__30722),
            .I(N__30711));
    InMux I__5461 (
            .O(N__30721),
            .I(N__30711));
    LocalMux I__5460 (
            .O(N__30718),
            .I(wdtick_cnt_1));
    LocalMux I__5459 (
            .O(N__30711),
            .I(wdtick_cnt_1));
    CascadeMux I__5458 (
            .O(N__30706),
            .I(N__30703));
    InMux I__5457 (
            .O(N__30703),
            .I(N__30698));
    InMux I__5456 (
            .O(N__30702),
            .I(N__30693));
    InMux I__5455 (
            .O(N__30701),
            .I(N__30693));
    LocalMux I__5454 (
            .O(N__30698),
            .I(wdtick_cnt_2));
    LocalMux I__5453 (
            .O(N__30693),
            .I(wdtick_cnt_2));
    CascadeMux I__5452 (
            .O(N__30688),
            .I(\ADC_VDC.n20490_cascade_ ));
    CascadeMux I__5451 (
            .O(N__30685),
            .I(\ADC_VDC.n11251_cascade_ ));
    CascadeMux I__5450 (
            .O(N__30682),
            .I(\ADC_VDC.n20523_cascade_ ));
    InMux I__5449 (
            .O(N__30679),
            .I(N__30676));
    LocalMux I__5448 (
            .O(N__30676),
            .I(N__30673));
    Span4Mux_h I__5447 (
            .O(N__30673),
            .I(N__30670));
    Odrv4 I__5446 (
            .O(N__30670),
            .I(\ADC_VDC.n21178 ));
    InMux I__5445 (
            .O(N__30667),
            .I(N__30664));
    LocalMux I__5444 (
            .O(N__30664),
            .I(N__30660));
    InMux I__5443 (
            .O(N__30663),
            .I(N__30657));
    Span4Mux_h I__5442 (
            .O(N__30660),
            .I(N__30654));
    LocalMux I__5441 (
            .O(N__30657),
            .I(\ADC_VDC.n20490 ));
    Odrv4 I__5440 (
            .O(N__30654),
            .I(\ADC_VDC.n20490 ));
    InMux I__5439 (
            .O(N__30649),
            .I(N__30646));
    LocalMux I__5438 (
            .O(N__30646),
            .I(N__30643));
    Span4Mux_h I__5437 (
            .O(N__30643),
            .I(N__30640));
    Odrv4 I__5436 (
            .O(N__30640),
            .I(\ADC_VDC.n21025 ));
    InMux I__5435 (
            .O(N__30637),
            .I(N__30633));
    InMux I__5434 (
            .O(N__30636),
            .I(N__30630));
    LocalMux I__5433 (
            .O(N__30633),
            .I(\ADC_VDC.n7_adj_1403 ));
    LocalMux I__5432 (
            .O(N__30630),
            .I(\ADC_VDC.n7_adj_1403 ));
    InMux I__5431 (
            .O(N__30625),
            .I(N__30616));
    InMux I__5430 (
            .O(N__30624),
            .I(N__30616));
    InMux I__5429 (
            .O(N__30623),
            .I(N__30616));
    LocalMux I__5428 (
            .O(N__30616),
            .I(\ADC_VDC.n20712 ));
    InMux I__5427 (
            .O(N__30613),
            .I(N__30610));
    LocalMux I__5426 (
            .O(N__30610),
            .I(N__30607));
    Span4Mux_v I__5425 (
            .O(N__30607),
            .I(N__30604));
    Odrv4 I__5424 (
            .O(N__30604),
            .I(\ADC_VDC.n11662 ));
    InMux I__5423 (
            .O(N__30601),
            .I(N__30598));
    LocalMux I__5422 (
            .O(N__30598),
            .I(\ADC_VDC.n21028 ));
    InMux I__5421 (
            .O(N__30595),
            .I(N__30591));
    InMux I__5420 (
            .O(N__30594),
            .I(N__30588));
    LocalMux I__5419 (
            .O(N__30591),
            .I(\ADC_VDC.genclk.t0off_14 ));
    LocalMux I__5418 (
            .O(N__30588),
            .I(\ADC_VDC.genclk.t0off_14 ));
    CascadeMux I__5417 (
            .O(N__30583),
            .I(N__30580));
    InMux I__5416 (
            .O(N__30580),
            .I(N__30576));
    InMux I__5415 (
            .O(N__30579),
            .I(N__30573));
    LocalMux I__5414 (
            .O(N__30576),
            .I(\ADC_VDC.genclk.t0off_9 ));
    LocalMux I__5413 (
            .O(N__30573),
            .I(\ADC_VDC.genclk.t0off_9 ));
    CascadeMux I__5412 (
            .O(N__30568),
            .I(N__30564));
    InMux I__5411 (
            .O(N__30567),
            .I(N__30561));
    InMux I__5410 (
            .O(N__30564),
            .I(N__30558));
    LocalMux I__5409 (
            .O(N__30561),
            .I(\ADC_VDC.genclk.t0off_15 ));
    LocalMux I__5408 (
            .O(N__30558),
            .I(\ADC_VDC.genclk.t0off_15 ));
    CascadeMux I__5407 (
            .O(N__30553),
            .I(N__30550));
    InMux I__5406 (
            .O(N__30550),
            .I(N__30546));
    InMux I__5405 (
            .O(N__30549),
            .I(N__30543));
    LocalMux I__5404 (
            .O(N__30546),
            .I(\ADC_VDC.genclk.t0off_11 ));
    LocalMux I__5403 (
            .O(N__30543),
            .I(\ADC_VDC.genclk.t0off_11 ));
    InMux I__5402 (
            .O(N__30538),
            .I(N__30535));
    LocalMux I__5401 (
            .O(N__30535),
            .I(\ADC_VDC.genclk.n28 ));
    CEMux I__5400 (
            .O(N__30532),
            .I(N__30529));
    LocalMux I__5399 (
            .O(N__30529),
            .I(N__30525));
    CEMux I__5398 (
            .O(N__30528),
            .I(N__30522));
    Span4Mux_h I__5397 (
            .O(N__30525),
            .I(N__30519));
    LocalMux I__5396 (
            .O(N__30522),
            .I(N__30516));
    Odrv4 I__5395 (
            .O(N__30519),
            .I(\ADC_VDC.genclk.n11721 ));
    Odrv4 I__5394 (
            .O(N__30516),
            .I(\ADC_VDC.genclk.n11721 ));
    CascadeMux I__5393 (
            .O(N__30511),
            .I(\ADC_VDC.n10112_cascade_ ));
    CEMux I__5392 (
            .O(N__30508),
            .I(N__30505));
    LocalMux I__5391 (
            .O(N__30505),
            .I(N__30502));
    Odrv4 I__5390 (
            .O(N__30502),
            .I(\ADC_VDC.n12793 ));
    CEMux I__5389 (
            .O(N__30499),
            .I(N__30496));
    LocalMux I__5388 (
            .O(N__30496),
            .I(\ADC_VDC.n17 ));
    SRMux I__5387 (
            .O(N__30493),
            .I(N__30490));
    LocalMux I__5386 (
            .O(N__30490),
            .I(N__30487));
    Span4Mux_h I__5385 (
            .O(N__30487),
            .I(N__30484));
    Odrv4 I__5384 (
            .O(N__30484),
            .I(\ADC_VDC.n4 ));
    InMux I__5383 (
            .O(N__30481),
            .I(N__30478));
    LocalMux I__5382 (
            .O(N__30478),
            .I(\ADC_VDC.n12 ));
    InMux I__5381 (
            .O(N__30475),
            .I(N__30472));
    LocalMux I__5380 (
            .O(N__30472),
            .I(\ADC_VDC.n72 ));
    InMux I__5379 (
            .O(N__30469),
            .I(N__30466));
    LocalMux I__5378 (
            .O(N__30466),
            .I(\ADC_VDC.n20710 ));
    CascadeMux I__5377 (
            .O(N__30463),
            .I(N__30458));
    CascadeMux I__5376 (
            .O(N__30462),
            .I(N__30455));
    InMux I__5375 (
            .O(N__30461),
            .I(N__30451));
    InMux I__5374 (
            .O(N__30458),
            .I(N__30448));
    InMux I__5373 (
            .O(N__30455),
            .I(N__30443));
    InMux I__5372 (
            .O(N__30454),
            .I(N__30443));
    LocalMux I__5371 (
            .O(N__30451),
            .I(N__30439));
    LocalMux I__5370 (
            .O(N__30448),
            .I(N__30436));
    LocalMux I__5369 (
            .O(N__30443),
            .I(N__30433));
    InMux I__5368 (
            .O(N__30442),
            .I(N__30430));
    Span4Mux_v I__5367 (
            .O(N__30439),
            .I(N__30427));
    Span4Mux_v I__5366 (
            .O(N__30436),
            .I(N__30422));
    Span4Mux_h I__5365 (
            .O(N__30433),
            .I(N__30422));
    LocalMux I__5364 (
            .O(N__30430),
            .I(eis_start));
    Odrv4 I__5363 (
            .O(N__30427),
            .I(eis_start));
    Odrv4 I__5362 (
            .O(N__30422),
            .I(eis_start));
    InMux I__5361 (
            .O(N__30415),
            .I(N__30412));
    LocalMux I__5360 (
            .O(N__30412),
            .I(n17357));
    CascadeMux I__5359 (
            .O(N__30409),
            .I(n11_adj_1620_cascade_));
    CEMux I__5358 (
            .O(N__30406),
            .I(N__30403));
    LocalMux I__5357 (
            .O(N__30403),
            .I(N__30400));
    Span4Mux_v I__5356 (
            .O(N__30400),
            .I(N__30397));
    Odrv4 I__5355 (
            .O(N__30397),
            .I(n11730));
    CascadeMux I__5354 (
            .O(N__30394),
            .I(N__30391));
    InMux I__5353 (
            .O(N__30391),
            .I(N__30387));
    InMux I__5352 (
            .O(N__30390),
            .I(N__30384));
    LocalMux I__5351 (
            .O(N__30387),
            .I(\ADC_VDC.genclk.t0off_6 ));
    LocalMux I__5350 (
            .O(N__30384),
            .I(\ADC_VDC.genclk.t0off_6 ));
    InMux I__5349 (
            .O(N__30379),
            .I(N__30375));
    InMux I__5348 (
            .O(N__30378),
            .I(N__30372));
    LocalMux I__5347 (
            .O(N__30375),
            .I(\ADC_VDC.genclk.t0off_1 ));
    LocalMux I__5346 (
            .O(N__30372),
            .I(\ADC_VDC.genclk.t0off_1 ));
    CascadeMux I__5345 (
            .O(N__30367),
            .I(N__30363));
    CascadeMux I__5344 (
            .O(N__30366),
            .I(N__30360));
    InMux I__5343 (
            .O(N__30363),
            .I(N__30357));
    InMux I__5342 (
            .O(N__30360),
            .I(N__30354));
    LocalMux I__5341 (
            .O(N__30357),
            .I(\ADC_VDC.genclk.t0off_4 ));
    LocalMux I__5340 (
            .O(N__30354),
            .I(\ADC_VDC.genclk.t0off_4 ));
    InMux I__5339 (
            .O(N__30349),
            .I(N__30345));
    InMux I__5338 (
            .O(N__30348),
            .I(N__30342));
    LocalMux I__5337 (
            .O(N__30345),
            .I(\ADC_VDC.genclk.t0off_0 ));
    LocalMux I__5336 (
            .O(N__30342),
            .I(\ADC_VDC.genclk.t0off_0 ));
    CascadeMux I__5335 (
            .O(N__30337),
            .I(\ADC_VDC.genclk.n21169_cascade_ ));
    InMux I__5334 (
            .O(N__30334),
            .I(N__30330));
    InMux I__5333 (
            .O(N__30333),
            .I(N__30327));
    LocalMux I__5332 (
            .O(N__30330),
            .I(\ADC_VDC.genclk.t0off_12 ));
    LocalMux I__5331 (
            .O(N__30327),
            .I(\ADC_VDC.genclk.t0off_12 ));
    CascadeMux I__5330 (
            .O(N__30322),
            .I(N__30319));
    InMux I__5329 (
            .O(N__30319),
            .I(N__30315));
    InMux I__5328 (
            .O(N__30318),
            .I(N__30312));
    LocalMux I__5327 (
            .O(N__30315),
            .I(\ADC_VDC.genclk.t0off_2 ));
    LocalMux I__5326 (
            .O(N__30312),
            .I(\ADC_VDC.genclk.t0off_2 ));
    CascadeMux I__5325 (
            .O(N__30307),
            .I(N__30303));
    InMux I__5324 (
            .O(N__30306),
            .I(N__30300));
    InMux I__5323 (
            .O(N__30303),
            .I(N__30297));
    LocalMux I__5322 (
            .O(N__30300),
            .I(\ADC_VDC.genclk.t0off_7 ));
    LocalMux I__5321 (
            .O(N__30297),
            .I(\ADC_VDC.genclk.t0off_7 ));
    InMux I__5320 (
            .O(N__30292),
            .I(N__30288));
    InMux I__5319 (
            .O(N__30291),
            .I(N__30285));
    LocalMux I__5318 (
            .O(N__30288),
            .I(\ADC_VDC.genclk.t0off_10 ));
    LocalMux I__5317 (
            .O(N__30285),
            .I(\ADC_VDC.genclk.t0off_10 ));
    InMux I__5316 (
            .O(N__30280),
            .I(N__30277));
    LocalMux I__5315 (
            .O(N__30277),
            .I(\ADC_VDC.genclk.n27 ));
    CascadeMux I__5314 (
            .O(N__30274),
            .I(N__30271));
    InMux I__5313 (
            .O(N__30271),
            .I(N__30267));
    InMux I__5312 (
            .O(N__30270),
            .I(N__30264));
    LocalMux I__5311 (
            .O(N__30267),
            .I(\ADC_VDC.genclk.t0off_13 ));
    LocalMux I__5310 (
            .O(N__30264),
            .I(\ADC_VDC.genclk.t0off_13 ));
    InMux I__5309 (
            .O(N__30259),
            .I(N__30255));
    InMux I__5308 (
            .O(N__30258),
            .I(N__30252));
    LocalMux I__5307 (
            .O(N__30255),
            .I(\ADC_VDC.genclk.t0off_8 ));
    LocalMux I__5306 (
            .O(N__30252),
            .I(\ADC_VDC.genclk.t0off_8 ));
    CascadeMux I__5305 (
            .O(N__30247),
            .I(N__30243));
    InMux I__5304 (
            .O(N__30246),
            .I(N__30240));
    InMux I__5303 (
            .O(N__30243),
            .I(N__30237));
    LocalMux I__5302 (
            .O(N__30240),
            .I(\ADC_VDC.genclk.t0off_5 ));
    LocalMux I__5301 (
            .O(N__30237),
            .I(\ADC_VDC.genclk.t0off_5 ));
    InMux I__5300 (
            .O(N__30232),
            .I(N__30228));
    InMux I__5299 (
            .O(N__30231),
            .I(N__30225));
    LocalMux I__5298 (
            .O(N__30228),
            .I(\ADC_VDC.genclk.t0off_3 ));
    LocalMux I__5297 (
            .O(N__30225),
            .I(\ADC_VDC.genclk.t0off_3 ));
    InMux I__5296 (
            .O(N__30220),
            .I(N__30217));
    LocalMux I__5295 (
            .O(N__30217),
            .I(N__30214));
    Sp12to4 I__5294 (
            .O(N__30214),
            .I(N__30211));
    Odrv12 I__5293 (
            .O(N__30211),
            .I(\ADC_VDC.genclk.n26 ));
    CascadeMux I__5292 (
            .O(N__30208),
            .I(n4_adj_1473_cascade_));
    InMux I__5291 (
            .O(N__30205),
            .I(N__30200));
    InMux I__5290 (
            .O(N__30204),
            .I(N__30197));
    InMux I__5289 (
            .O(N__30203),
            .I(N__30194));
    LocalMux I__5288 (
            .O(N__30200),
            .I(acadc_skipCount_13));
    LocalMux I__5287 (
            .O(N__30197),
            .I(acadc_skipCount_13));
    LocalMux I__5286 (
            .O(N__30194),
            .I(acadc_skipCount_13));
    InMux I__5285 (
            .O(N__30187),
            .I(N__30182));
    InMux I__5284 (
            .O(N__30186),
            .I(N__30179));
    InMux I__5283 (
            .O(N__30185),
            .I(N__30176));
    LocalMux I__5282 (
            .O(N__30182),
            .I(N__30173));
    LocalMux I__5281 (
            .O(N__30179),
            .I(N__30170));
    LocalMux I__5280 (
            .O(N__30176),
            .I(buf_dds1_10));
    Odrv4 I__5279 (
            .O(N__30173),
            .I(buf_dds1_10));
    Odrv4 I__5278 (
            .O(N__30170),
            .I(buf_dds1_10));
    InMux I__5277 (
            .O(N__30163),
            .I(N__30160));
    LocalMux I__5276 (
            .O(N__30160),
            .I(n22147));
    InMux I__5275 (
            .O(N__30157),
            .I(N__30154));
    LocalMux I__5274 (
            .O(N__30154),
            .I(N__30151));
    Span4Mux_v I__5273 (
            .O(N__30151),
            .I(N__30148));
    Odrv4 I__5272 (
            .O(N__30148),
            .I(n22150));
    CascadeMux I__5271 (
            .O(N__30145),
            .I(n20690_cascade_));
    InMux I__5270 (
            .O(N__30142),
            .I(N__30134));
    InMux I__5269 (
            .O(N__30141),
            .I(N__30134));
    InMux I__5268 (
            .O(N__30140),
            .I(N__30128));
    InMux I__5267 (
            .O(N__30139),
            .I(N__30128));
    LocalMux I__5266 (
            .O(N__30134),
            .I(N__30125));
    InMux I__5265 (
            .O(N__30133),
            .I(N__30122));
    LocalMux I__5264 (
            .O(N__30128),
            .I(N__30119));
    Span4Mux_h I__5263 (
            .O(N__30125),
            .I(N__30116));
    LocalMux I__5262 (
            .O(N__30122),
            .I(N__30111));
    Span4Mux_v I__5261 (
            .O(N__30119),
            .I(N__30111));
    Odrv4 I__5260 (
            .O(N__30116),
            .I(acadc_trig));
    Odrv4 I__5259 (
            .O(N__30111),
            .I(acadc_trig));
    InMux I__5258 (
            .O(N__30106),
            .I(N__30103));
    LocalMux I__5257 (
            .O(N__30103),
            .I(n20529));
    InMux I__5256 (
            .O(N__30100),
            .I(N__30096));
    CascadeMux I__5255 (
            .O(N__30099),
            .I(N__30093));
    LocalMux I__5254 (
            .O(N__30096),
            .I(N__30090));
    InMux I__5253 (
            .O(N__30093),
            .I(N__30087));
    Span4Mux_h I__5252 (
            .O(N__30090),
            .I(N__30084));
    LocalMux I__5251 (
            .O(N__30087),
            .I(eis_end));
    Odrv4 I__5250 (
            .O(N__30084),
            .I(eis_end));
    InMux I__5249 (
            .O(N__30079),
            .I(N__30075));
    InMux I__5248 (
            .O(N__30078),
            .I(N__30072));
    LocalMux I__5247 (
            .O(N__30075),
            .I(N__30069));
    LocalMux I__5246 (
            .O(N__30072),
            .I(N__30064));
    Span4Mux_v I__5245 (
            .O(N__30069),
            .I(N__30064));
    Span4Mux_h I__5244 (
            .O(N__30064),
            .I(N__30061));
    Odrv4 I__5243 (
            .O(N__30061),
            .I(n8_adj_1536));
    IoInMux I__5242 (
            .O(N__30058),
            .I(N__30055));
    LocalMux I__5241 (
            .O(N__30055),
            .I(N__30052));
    Span4Mux_s2_h I__5240 (
            .O(N__30052),
            .I(N__30049));
    Sp12to4 I__5239 (
            .O(N__30049),
            .I(N__30046));
    Span12Mux_v I__5238 (
            .O(N__30046),
            .I(N__30042));
    InMux I__5237 (
            .O(N__30045),
            .I(N__30038));
    Span12Mux_h I__5236 (
            .O(N__30042),
            .I(N__30035));
    InMux I__5235 (
            .O(N__30041),
            .I(N__30032));
    LocalMux I__5234 (
            .O(N__30038),
            .I(N__30029));
    Odrv12 I__5233 (
            .O(N__30035),
            .I(AMPV_POW));
    LocalMux I__5232 (
            .O(N__30032),
            .I(AMPV_POW));
    Odrv4 I__5231 (
            .O(N__30029),
            .I(AMPV_POW));
    InMux I__5230 (
            .O(N__30022),
            .I(N__30018));
    InMux I__5229 (
            .O(N__30021),
            .I(N__30015));
    LocalMux I__5228 (
            .O(N__30018),
            .I(N__30009));
    LocalMux I__5227 (
            .O(N__30015),
            .I(N__30006));
    CascadeMux I__5226 (
            .O(N__30014),
            .I(N__30000));
    CascadeMux I__5225 (
            .O(N__30013),
            .I(N__29996));
    CascadeMux I__5224 (
            .O(N__30012),
            .I(N__29991));
    Span4Mux_h I__5223 (
            .O(N__30009),
            .I(N__29987));
    Span4Mux_h I__5222 (
            .O(N__30006),
            .I(N__29984));
    InMux I__5221 (
            .O(N__30005),
            .I(N__29981));
    InMux I__5220 (
            .O(N__30004),
            .I(N__29974));
    InMux I__5219 (
            .O(N__30003),
            .I(N__29974));
    InMux I__5218 (
            .O(N__30000),
            .I(N__29974));
    InMux I__5217 (
            .O(N__29999),
            .I(N__29961));
    InMux I__5216 (
            .O(N__29996),
            .I(N__29961));
    InMux I__5215 (
            .O(N__29995),
            .I(N__29961));
    InMux I__5214 (
            .O(N__29994),
            .I(N__29961));
    InMux I__5213 (
            .O(N__29991),
            .I(N__29961));
    InMux I__5212 (
            .O(N__29990),
            .I(N__29961));
    Odrv4 I__5211 (
            .O(N__29987),
            .I(DTRIG_N_910));
    Odrv4 I__5210 (
            .O(N__29984),
            .I(DTRIG_N_910));
    LocalMux I__5209 (
            .O(N__29981),
            .I(DTRIG_N_910));
    LocalMux I__5208 (
            .O(N__29974),
            .I(DTRIG_N_910));
    LocalMux I__5207 (
            .O(N__29961),
            .I(DTRIG_N_910));
    InMux I__5206 (
            .O(N__29950),
            .I(N__29946));
    InMux I__5205 (
            .O(N__29949),
            .I(N__29943));
    LocalMux I__5204 (
            .O(N__29946),
            .I(N__29940));
    LocalMux I__5203 (
            .O(N__29943),
            .I(N__29937));
    Span4Mux_h I__5202 (
            .O(N__29940),
            .I(N__29924));
    Span4Mux_v I__5201 (
            .O(N__29937),
            .I(N__29921));
    InMux I__5200 (
            .O(N__29936),
            .I(N__29918));
    InMux I__5199 (
            .O(N__29935),
            .I(N__29909));
    InMux I__5198 (
            .O(N__29934),
            .I(N__29909));
    InMux I__5197 (
            .O(N__29933),
            .I(N__29909));
    InMux I__5196 (
            .O(N__29932),
            .I(N__29909));
    InMux I__5195 (
            .O(N__29931),
            .I(N__29898));
    InMux I__5194 (
            .O(N__29930),
            .I(N__29898));
    InMux I__5193 (
            .O(N__29929),
            .I(N__29898));
    InMux I__5192 (
            .O(N__29928),
            .I(N__29898));
    InMux I__5191 (
            .O(N__29927),
            .I(N__29898));
    Odrv4 I__5190 (
            .O(N__29924),
            .I(adc_state_1));
    Odrv4 I__5189 (
            .O(N__29921),
            .I(adc_state_1));
    LocalMux I__5188 (
            .O(N__29918),
            .I(adc_state_1));
    LocalMux I__5187 (
            .O(N__29909),
            .I(adc_state_1));
    LocalMux I__5186 (
            .O(N__29898),
            .I(adc_state_1));
    InMux I__5185 (
            .O(N__29887),
            .I(N__29883));
    InMux I__5184 (
            .O(N__29886),
            .I(N__29880));
    LocalMux I__5183 (
            .O(N__29883),
            .I(N__29876));
    LocalMux I__5182 (
            .O(N__29880),
            .I(N__29873));
    InMux I__5181 (
            .O(N__29879),
            .I(N__29870));
    Odrv4 I__5180 (
            .O(N__29876),
            .I(n10503));
    Odrv4 I__5179 (
            .O(N__29873),
            .I(n10503));
    LocalMux I__5178 (
            .O(N__29870),
            .I(n10503));
    InMux I__5177 (
            .O(N__29863),
            .I(N__29859));
    InMux I__5176 (
            .O(N__29862),
            .I(N__29851));
    LocalMux I__5175 (
            .O(N__29859),
            .I(N__29848));
    CascadeMux I__5174 (
            .O(N__29858),
            .I(N__29842));
    CascadeMux I__5173 (
            .O(N__29857),
            .I(N__29838));
    InMux I__5172 (
            .O(N__29856),
            .I(N__29830));
    InMux I__5171 (
            .O(N__29855),
            .I(N__29830));
    InMux I__5170 (
            .O(N__29854),
            .I(N__29830));
    LocalMux I__5169 (
            .O(N__29851),
            .I(N__29827));
    Span4Mux_v I__5168 (
            .O(N__29848),
            .I(N__29824));
    InMux I__5167 (
            .O(N__29847),
            .I(N__29819));
    InMux I__5166 (
            .O(N__29846),
            .I(N__29819));
    InMux I__5165 (
            .O(N__29845),
            .I(N__29808));
    InMux I__5164 (
            .O(N__29842),
            .I(N__29808));
    InMux I__5163 (
            .O(N__29841),
            .I(N__29808));
    InMux I__5162 (
            .O(N__29838),
            .I(N__29808));
    InMux I__5161 (
            .O(N__29837),
            .I(N__29808));
    LocalMux I__5160 (
            .O(N__29830),
            .I(N__29805));
    Odrv12 I__5159 (
            .O(N__29827),
            .I(DTRIG_N_910_adj_1444));
    Odrv4 I__5158 (
            .O(N__29824),
            .I(DTRIG_N_910_adj_1444));
    LocalMux I__5157 (
            .O(N__29819),
            .I(DTRIG_N_910_adj_1444));
    LocalMux I__5156 (
            .O(N__29808),
            .I(DTRIG_N_910_adj_1444));
    Odrv12 I__5155 (
            .O(N__29805),
            .I(DTRIG_N_910_adj_1444));
    InMux I__5154 (
            .O(N__29794),
            .I(N__29788));
    CascadeMux I__5153 (
            .O(N__29793),
            .I(N__29784));
    InMux I__5152 (
            .O(N__29792),
            .I(N__29776));
    InMux I__5151 (
            .O(N__29791),
            .I(N__29776));
    LocalMux I__5150 (
            .O(N__29788),
            .I(N__29773));
    InMux I__5149 (
            .O(N__29787),
            .I(N__29768));
    InMux I__5148 (
            .O(N__29784),
            .I(N__29768));
    InMux I__5147 (
            .O(N__29783),
            .I(N__29757));
    InMux I__5146 (
            .O(N__29782),
            .I(N__29757));
    InMux I__5145 (
            .O(N__29781),
            .I(N__29757));
    LocalMux I__5144 (
            .O(N__29776),
            .I(N__29754));
    Span4Mux_h I__5143 (
            .O(N__29773),
            .I(N__29749));
    LocalMux I__5142 (
            .O(N__29768),
            .I(N__29749));
    InMux I__5141 (
            .O(N__29767),
            .I(N__29742));
    InMux I__5140 (
            .O(N__29766),
            .I(N__29742));
    InMux I__5139 (
            .O(N__29765),
            .I(N__29742));
    InMux I__5138 (
            .O(N__29764),
            .I(N__29739));
    LocalMux I__5137 (
            .O(N__29757),
            .I(N__29736));
    Odrv4 I__5136 (
            .O(N__29754),
            .I(adc_state_1_adj_1410));
    Odrv4 I__5135 (
            .O(N__29749),
            .I(adc_state_1_adj_1410));
    LocalMux I__5134 (
            .O(N__29742),
            .I(adc_state_1_adj_1410));
    LocalMux I__5133 (
            .O(N__29739),
            .I(adc_state_1_adj_1410));
    Odrv4 I__5132 (
            .O(N__29736),
            .I(adc_state_1_adj_1410));
    IoInMux I__5131 (
            .O(N__29725),
            .I(N__29722));
    LocalMux I__5130 (
            .O(N__29722),
            .I(N__29719));
    Span4Mux_s2_h I__5129 (
            .O(N__29719),
            .I(N__29716));
    Sp12to4 I__5128 (
            .O(N__29716),
            .I(N__29712));
    InMux I__5127 (
            .O(N__29715),
            .I(N__29709));
    Span12Mux_v I__5126 (
            .O(N__29712),
            .I(N__29706));
    LocalMux I__5125 (
            .O(N__29709),
            .I(N__29702));
    Span12Mux_h I__5124 (
            .O(N__29706),
            .I(N__29699));
    InMux I__5123 (
            .O(N__29705),
            .I(N__29696));
    Span4Mux_v I__5122 (
            .O(N__29702),
            .I(N__29693));
    Odrv12 I__5121 (
            .O(N__29699),
            .I(VAC_OSR1));
    LocalMux I__5120 (
            .O(N__29696),
            .I(VAC_OSR1));
    Odrv4 I__5119 (
            .O(N__29693),
            .I(VAC_OSR1));
    CascadeMux I__5118 (
            .O(N__29686),
            .I(n21940_cascade_));
    CascadeMux I__5117 (
            .O(N__29683),
            .I(n30_adj_1490_cascade_));
    InMux I__5116 (
            .O(N__29680),
            .I(N__29677));
    LocalMux I__5115 (
            .O(N__29677),
            .I(n26_adj_1495));
    CascadeMux I__5114 (
            .O(N__29674),
            .I(N__29671));
    InMux I__5113 (
            .O(N__29671),
            .I(N__29668));
    LocalMux I__5112 (
            .O(N__29668),
            .I(N__29665));
    Span4Mux_h I__5111 (
            .O(N__29665),
            .I(N__29662));
    Odrv4 I__5110 (
            .O(N__29662),
            .I(n21109));
    CascadeMux I__5109 (
            .O(N__29659),
            .I(n22111_cascade_));
    InMux I__5108 (
            .O(N__29656),
            .I(N__29653));
    LocalMux I__5107 (
            .O(N__29653),
            .I(n22114));
    CascadeMux I__5106 (
            .O(N__29650),
            .I(n16539_cascade_));
    CascadeMux I__5105 (
            .O(N__29647),
            .I(n17_adj_1601_cascade_));
    InMux I__5104 (
            .O(N__29644),
            .I(N__29641));
    LocalMux I__5103 (
            .O(N__29641),
            .I(n16547));
    CascadeMux I__5102 (
            .O(N__29638),
            .I(n16547_cascade_));
    CascadeMux I__5101 (
            .O(N__29635),
            .I(n13_cascade_));
    InMux I__5100 (
            .O(N__29632),
            .I(N__29629));
    LocalMux I__5099 (
            .O(N__29629),
            .I(N__29626));
    Span12Mux_h I__5098 (
            .O(N__29626),
            .I(N__29623));
    Odrv12 I__5097 (
            .O(N__29623),
            .I(n19_adj_1482));
    CascadeMux I__5096 (
            .O(N__29620),
            .I(N__29617));
    InMux I__5095 (
            .O(N__29617),
            .I(N__29614));
    LocalMux I__5094 (
            .O(N__29614),
            .I(N__29611));
    Span4Mux_h I__5093 (
            .O(N__29611),
            .I(N__29608));
    Span4Mux_h I__5092 (
            .O(N__29608),
            .I(N__29604));
    CascadeMux I__5091 (
            .O(N__29607),
            .I(N__29601));
    Span4Mux_v I__5090 (
            .O(N__29604),
            .I(N__29598));
    InMux I__5089 (
            .O(N__29601),
            .I(N__29595));
    Odrv4 I__5088 (
            .O(N__29598),
            .I(buf_readRTD_6));
    LocalMux I__5087 (
            .O(N__29595),
            .I(buf_readRTD_6));
    CascadeMux I__5086 (
            .O(N__29590),
            .I(n21937_cascade_));
    InMux I__5085 (
            .O(N__29587),
            .I(N__29583));
    InMux I__5084 (
            .O(N__29586),
            .I(N__29580));
    LocalMux I__5083 (
            .O(N__29583),
            .I(N__29577));
    LocalMux I__5082 (
            .O(N__29580),
            .I(N__29573));
    Span4Mux_h I__5081 (
            .O(N__29577),
            .I(N__29570));
    InMux I__5080 (
            .O(N__29576),
            .I(N__29567));
    Span4Mux_h I__5079 (
            .O(N__29573),
            .I(N__29562));
    Span4Mux_h I__5078 (
            .O(N__29570),
            .I(N__29562));
    LocalMux I__5077 (
            .O(N__29567),
            .I(buf_adcdata_iac_14));
    Odrv4 I__5076 (
            .O(N__29562),
            .I(buf_adcdata_iac_14));
    InMux I__5075 (
            .O(N__29557),
            .I(N__29552));
    InMux I__5074 (
            .O(N__29556),
            .I(N__29549));
    InMux I__5073 (
            .O(N__29555),
            .I(N__29546));
    LocalMux I__5072 (
            .O(N__29552),
            .I(N__29543));
    LocalMux I__5071 (
            .O(N__29549),
            .I(buf_dds1_11));
    LocalMux I__5070 (
            .O(N__29546),
            .I(buf_dds1_11));
    Odrv4 I__5069 (
            .O(N__29543),
            .I(buf_dds1_11));
    InMux I__5068 (
            .O(N__29536),
            .I(N__29533));
    LocalMux I__5067 (
            .O(N__29533),
            .I(N__29530));
    Span12Mux_v I__5066 (
            .O(N__29530),
            .I(N__29527));
    Odrv12 I__5065 (
            .O(N__29527),
            .I(n22075));
    InMux I__5064 (
            .O(N__29524),
            .I(N__29521));
    LocalMux I__5063 (
            .O(N__29521),
            .I(N__29518));
    Span4Mux_h I__5062 (
            .O(N__29518),
            .I(N__29515));
    Span4Mux_h I__5061 (
            .O(N__29515),
            .I(N__29512));
    Odrv4 I__5060 (
            .O(N__29512),
            .I(n22078));
    InMux I__5059 (
            .O(N__29509),
            .I(N__29505));
    InMux I__5058 (
            .O(N__29508),
            .I(N__29502));
    LocalMux I__5057 (
            .O(N__29505),
            .I(N__29499));
    LocalMux I__5056 (
            .O(N__29502),
            .I(N__29493));
    Span4Mux_v I__5055 (
            .O(N__29499),
            .I(N__29493));
    InMux I__5054 (
            .O(N__29498),
            .I(N__29490));
    Span4Mux_v I__5053 (
            .O(N__29493),
            .I(N__29487));
    LocalMux I__5052 (
            .O(N__29490),
            .I(buf_dds1_5));
    Odrv4 I__5051 (
            .O(N__29487),
            .I(buf_dds1_5));
    InMux I__5050 (
            .O(N__29482),
            .I(N__29479));
    LocalMux I__5049 (
            .O(N__29479),
            .I(n7));
    InMux I__5048 (
            .O(N__29476),
            .I(N__29459));
    InMux I__5047 (
            .O(N__29475),
            .I(N__29459));
    InMux I__5046 (
            .O(N__29474),
            .I(N__29459));
    InMux I__5045 (
            .O(N__29473),
            .I(N__29459));
    InMux I__5044 (
            .O(N__29472),
            .I(N__29459));
    InMux I__5043 (
            .O(N__29471),
            .I(N__29454));
    InMux I__5042 (
            .O(N__29470),
            .I(N__29454));
    LocalMux I__5041 (
            .O(N__29459),
            .I(n12214));
    LocalMux I__5040 (
            .O(N__29454),
            .I(n12214));
    InMux I__5039 (
            .O(N__29449),
            .I(N__29440));
    InMux I__5038 (
            .O(N__29448),
            .I(N__29440));
    InMux I__5037 (
            .O(N__29447),
            .I(N__29440));
    LocalMux I__5036 (
            .O(N__29440),
            .I(comm_cmd_4));
    CascadeMux I__5035 (
            .O(N__29437),
            .I(N__29433));
    InMux I__5034 (
            .O(N__29436),
            .I(N__29425));
    InMux I__5033 (
            .O(N__29433),
            .I(N__29425));
    InMux I__5032 (
            .O(N__29432),
            .I(N__29425));
    LocalMux I__5031 (
            .O(N__29425),
            .I(comm_cmd_6));
    InMux I__5030 (
            .O(N__29422),
            .I(N__29417));
    InMux I__5029 (
            .O(N__29421),
            .I(N__29412));
    InMux I__5028 (
            .O(N__29420),
            .I(N__29412));
    LocalMux I__5027 (
            .O(N__29417),
            .I(comm_cmd_5));
    LocalMux I__5026 (
            .O(N__29412),
            .I(comm_cmd_5));
    CascadeMux I__5025 (
            .O(N__29407),
            .I(n8_adj_1522_cascade_));
    CascadeMux I__5024 (
            .O(N__29404),
            .I(n12214_cascade_));
    InMux I__5023 (
            .O(N__29401),
            .I(N__29398));
    LocalMux I__5022 (
            .O(N__29398),
            .I(N__29394));
    InMux I__5021 (
            .O(N__29397),
            .I(N__29390));
    Span4Mux_v I__5020 (
            .O(N__29394),
            .I(N__29387));
    InMux I__5019 (
            .O(N__29393),
            .I(N__29384));
    LocalMux I__5018 (
            .O(N__29390),
            .I(buf_dds1_13));
    Odrv4 I__5017 (
            .O(N__29387),
            .I(buf_dds1_13));
    LocalMux I__5016 (
            .O(N__29384),
            .I(buf_dds1_13));
    InMux I__5015 (
            .O(N__29377),
            .I(N__29374));
    LocalMux I__5014 (
            .O(N__29374),
            .I(N__29371));
    Span4Mux_v I__5013 (
            .O(N__29371),
            .I(N__29368));
    Span4Mux_h I__5012 (
            .O(N__29368),
            .I(N__29365));
    Span4Mux_v I__5011 (
            .O(N__29365),
            .I(N__29362));
    Span4Mux_v I__5010 (
            .O(N__29362),
            .I(N__29359));
    Odrv4 I__5009 (
            .O(N__29359),
            .I(THERMOSTAT));
    InMux I__5008 (
            .O(N__29356),
            .I(N__29353));
    LocalMux I__5007 (
            .O(N__29353),
            .I(N__29350));
    Odrv4 I__5006 (
            .O(N__29350),
            .I(buf_control_7));
    CascadeMux I__5005 (
            .O(N__29347),
            .I(n21050_cascade_));
    CEMux I__5004 (
            .O(N__29344),
            .I(N__29341));
    LocalMux I__5003 (
            .O(N__29341),
            .I(N__29338));
    Span4Mux_h I__5002 (
            .O(N__29338),
            .I(N__29335));
    Span4Mux_h I__5001 (
            .O(N__29335),
            .I(N__29332));
    Odrv4 I__5000 (
            .O(N__29332),
            .I(n11905));
    CascadeMux I__4999 (
            .O(N__29329),
            .I(N__29326));
    InMux I__4998 (
            .O(N__29326),
            .I(N__29322));
    CascadeMux I__4997 (
            .O(N__29325),
            .I(N__29319));
    LocalMux I__4996 (
            .O(N__29322),
            .I(N__29314));
    InMux I__4995 (
            .O(N__29319),
            .I(N__29311));
    CascadeMux I__4994 (
            .O(N__29318),
            .I(N__29308));
    InMux I__4993 (
            .O(N__29317),
            .I(N__29305));
    Sp12to4 I__4992 (
            .O(N__29314),
            .I(N__29300));
    LocalMux I__4991 (
            .O(N__29311),
            .I(N__29300));
    InMux I__4990 (
            .O(N__29308),
            .I(N__29297));
    LocalMux I__4989 (
            .O(N__29305),
            .I(N__29293));
    Span12Mux_v I__4988 (
            .O(N__29300),
            .I(N__29288));
    LocalMux I__4987 (
            .O(N__29297),
            .I(N__29288));
    InMux I__4986 (
            .O(N__29296),
            .I(N__29285));
    Span4Mux_v I__4985 (
            .O(N__29293),
            .I(N__29282));
    Odrv12 I__4984 (
            .O(N__29288),
            .I(buf_cfgRTD_6));
    LocalMux I__4983 (
            .O(N__29285),
            .I(buf_cfgRTD_6));
    Odrv4 I__4982 (
            .O(N__29282),
            .I(buf_cfgRTD_6));
    CascadeMux I__4981 (
            .O(N__29275),
            .I(n11882_cascade_));
    InMux I__4980 (
            .O(N__29272),
            .I(N__29268));
    InMux I__4979 (
            .O(N__29271),
            .I(N__29265));
    LocalMux I__4978 (
            .O(N__29268),
            .I(\ADC_VDC.avg_cnt_7 ));
    LocalMux I__4977 (
            .O(N__29265),
            .I(\ADC_VDC.avg_cnt_7 ));
    InMux I__4976 (
            .O(N__29260),
            .I(\ADC_VDC.n19405 ));
    CascadeMux I__4975 (
            .O(N__29257),
            .I(N__29254));
    InMux I__4974 (
            .O(N__29254),
            .I(N__29250));
    InMux I__4973 (
            .O(N__29253),
            .I(N__29247));
    LocalMux I__4972 (
            .O(N__29250),
            .I(N__29244));
    LocalMux I__4971 (
            .O(N__29247),
            .I(\ADC_VDC.avg_cnt_8 ));
    Odrv12 I__4970 (
            .O(N__29244),
            .I(\ADC_VDC.avg_cnt_8 ));
    InMux I__4969 (
            .O(N__29239),
            .I(bfn_11_8_0_));
    InMux I__4968 (
            .O(N__29236),
            .I(N__29232));
    InMux I__4967 (
            .O(N__29235),
            .I(N__29229));
    LocalMux I__4966 (
            .O(N__29232),
            .I(\ADC_VDC.avg_cnt_9 ));
    LocalMux I__4965 (
            .O(N__29229),
            .I(\ADC_VDC.avg_cnt_9 ));
    InMux I__4964 (
            .O(N__29224),
            .I(\ADC_VDC.n19407 ));
    InMux I__4963 (
            .O(N__29221),
            .I(N__29217));
    InMux I__4962 (
            .O(N__29220),
            .I(N__29214));
    LocalMux I__4961 (
            .O(N__29217),
            .I(\ADC_VDC.avg_cnt_10 ));
    LocalMux I__4960 (
            .O(N__29214),
            .I(\ADC_VDC.avg_cnt_10 ));
    InMux I__4959 (
            .O(N__29209),
            .I(\ADC_VDC.n19408 ));
    InMux I__4958 (
            .O(N__29206),
            .I(\ADC_VDC.n19409 ));
    InMux I__4957 (
            .O(N__29203),
            .I(N__29199));
    InMux I__4956 (
            .O(N__29202),
            .I(N__29196));
    LocalMux I__4955 (
            .O(N__29199),
            .I(\ADC_VDC.avg_cnt_11 ));
    LocalMux I__4954 (
            .O(N__29196),
            .I(\ADC_VDC.avg_cnt_11 ));
    CEMux I__4953 (
            .O(N__29191),
            .I(N__29187));
    CEMux I__4952 (
            .O(N__29190),
            .I(N__29183));
    LocalMux I__4951 (
            .O(N__29187),
            .I(N__29180));
    CEMux I__4950 (
            .O(N__29186),
            .I(N__29174));
    LocalMux I__4949 (
            .O(N__29183),
            .I(N__29169));
    Span4Mux_v I__4948 (
            .O(N__29180),
            .I(N__29169));
    CEMux I__4947 (
            .O(N__29179),
            .I(N__29166));
    CEMux I__4946 (
            .O(N__29178),
            .I(N__29163));
    CEMux I__4945 (
            .O(N__29177),
            .I(N__29159));
    LocalMux I__4944 (
            .O(N__29174),
            .I(N__29152));
    Span4Mux_v I__4943 (
            .O(N__29169),
            .I(N__29152));
    LocalMux I__4942 (
            .O(N__29166),
            .I(N__29152));
    LocalMux I__4941 (
            .O(N__29163),
            .I(N__29149));
    CEMux I__4940 (
            .O(N__29162),
            .I(N__29146));
    LocalMux I__4939 (
            .O(N__29159),
            .I(N__29143));
    Span4Mux_v I__4938 (
            .O(N__29152),
            .I(N__29140));
    Span4Mux_v I__4937 (
            .O(N__29149),
            .I(N__29135));
    LocalMux I__4936 (
            .O(N__29146),
            .I(N__29135));
    Span4Mux_h I__4935 (
            .O(N__29143),
            .I(N__29131));
    Span4Mux_h I__4934 (
            .O(N__29140),
            .I(N__29128));
    Span4Mux_h I__4933 (
            .O(N__29135),
            .I(N__29125));
    InMux I__4932 (
            .O(N__29134),
            .I(N__29122));
    Odrv4 I__4931 (
            .O(N__29131),
            .I(\ADC_VDC.n13060 ));
    Odrv4 I__4930 (
            .O(N__29128),
            .I(\ADC_VDC.n13060 ));
    Odrv4 I__4929 (
            .O(N__29125),
            .I(\ADC_VDC.n13060 ));
    LocalMux I__4928 (
            .O(N__29122),
            .I(\ADC_VDC.n13060 ));
    SRMux I__4927 (
            .O(N__29113),
            .I(N__29110));
    LocalMux I__4926 (
            .O(N__29110),
            .I(N__29105));
    SRMux I__4925 (
            .O(N__29109),
            .I(N__29100));
    SRMux I__4924 (
            .O(N__29108),
            .I(N__29096));
    Span4Mux_v I__4923 (
            .O(N__29105),
            .I(N__29092));
    SRMux I__4922 (
            .O(N__29104),
            .I(N__29089));
    SRMux I__4921 (
            .O(N__29103),
            .I(N__29086));
    LocalMux I__4920 (
            .O(N__29100),
            .I(N__29083));
    SRMux I__4919 (
            .O(N__29099),
            .I(N__29080));
    LocalMux I__4918 (
            .O(N__29096),
            .I(N__29077));
    SRMux I__4917 (
            .O(N__29095),
            .I(N__29074));
    Span4Mux_v I__4916 (
            .O(N__29092),
            .I(N__29069));
    LocalMux I__4915 (
            .O(N__29089),
            .I(N__29069));
    LocalMux I__4914 (
            .O(N__29086),
            .I(N__29066));
    Span4Mux_h I__4913 (
            .O(N__29083),
            .I(N__29061));
    LocalMux I__4912 (
            .O(N__29080),
            .I(N__29061));
    Span4Mux_h I__4911 (
            .O(N__29077),
            .I(N__29056));
    LocalMux I__4910 (
            .O(N__29074),
            .I(N__29056));
    Span4Mux_v I__4909 (
            .O(N__29069),
            .I(N__29051));
    Span4Mux_h I__4908 (
            .O(N__29066),
            .I(N__29051));
    Span4Mux_v I__4907 (
            .O(N__29061),
            .I(N__29048));
    Span4Mux_v I__4906 (
            .O(N__29056),
            .I(N__29045));
    Span4Mux_v I__4905 (
            .O(N__29051),
            .I(N__29042));
    Odrv4 I__4904 (
            .O(N__29048),
            .I(\ADC_VDC.n14900 ));
    Odrv4 I__4903 (
            .O(N__29045),
            .I(\ADC_VDC.n14900 ));
    Odrv4 I__4902 (
            .O(N__29042),
            .I(\ADC_VDC.n14900 ));
    CascadeMux I__4901 (
            .O(N__29035),
            .I(n23_adj_1510_cascade_));
    InMux I__4900 (
            .O(N__29032),
            .I(N__29029));
    LocalMux I__4899 (
            .O(N__29029),
            .I(N__29026));
    Span4Mux_v I__4898 (
            .O(N__29026),
            .I(N__29023));
    Span4Mux_h I__4897 (
            .O(N__29023),
            .I(N__29020));
    Odrv4 I__4896 (
            .O(N__29020),
            .I(n20833));
    InMux I__4895 (
            .O(N__29017),
            .I(N__29014));
    LocalMux I__4894 (
            .O(N__29014),
            .I(N__29011));
    Span4Mux_v I__4893 (
            .O(N__29011),
            .I(N__29008));
    Span4Mux_h I__4892 (
            .O(N__29008),
            .I(N__29005));
    Span4Mux_h I__4891 (
            .O(N__29005),
            .I(N__29002));
    Odrv4 I__4890 (
            .O(N__29002),
            .I(buf_data_iac_20));
    CascadeMux I__4889 (
            .O(N__28999),
            .I(N__28996));
    InMux I__4888 (
            .O(N__28996),
            .I(N__28993));
    LocalMux I__4887 (
            .O(N__28993),
            .I(N__28990));
    Span4Mux_h I__4886 (
            .O(N__28990),
            .I(N__28987));
    Span4Mux_v I__4885 (
            .O(N__28987),
            .I(N__28984));
    Odrv4 I__4884 (
            .O(N__28984),
            .I(n20810));
    InMux I__4883 (
            .O(N__28981),
            .I(N__28968));
    InMux I__4882 (
            .O(N__28980),
            .I(N__28968));
    InMux I__4881 (
            .O(N__28979),
            .I(N__28955));
    InMux I__4880 (
            .O(N__28978),
            .I(N__28955));
    InMux I__4879 (
            .O(N__28977),
            .I(N__28955));
    InMux I__4878 (
            .O(N__28976),
            .I(N__28955));
    InMux I__4877 (
            .O(N__28975),
            .I(N__28955));
    InMux I__4876 (
            .O(N__28974),
            .I(N__28955));
    SRMux I__4875 (
            .O(N__28973),
            .I(N__28944));
    LocalMux I__4874 (
            .O(N__28968),
            .I(N__28937));
    LocalMux I__4873 (
            .O(N__28955),
            .I(N__28934));
    InMux I__4872 (
            .O(N__28954),
            .I(N__28931));
    InMux I__4871 (
            .O(N__28953),
            .I(N__28916));
    InMux I__4870 (
            .O(N__28952),
            .I(N__28916));
    InMux I__4869 (
            .O(N__28951),
            .I(N__28916));
    InMux I__4868 (
            .O(N__28950),
            .I(N__28916));
    InMux I__4867 (
            .O(N__28949),
            .I(N__28916));
    InMux I__4866 (
            .O(N__28948),
            .I(N__28916));
    InMux I__4865 (
            .O(N__28947),
            .I(N__28916));
    LocalMux I__4864 (
            .O(N__28944),
            .I(N__28913));
    InMux I__4863 (
            .O(N__28943),
            .I(N__28910));
    CascadeMux I__4862 (
            .O(N__28942),
            .I(N__28904));
    InMux I__4861 (
            .O(N__28941),
            .I(N__28899));
    InMux I__4860 (
            .O(N__28940),
            .I(N__28899));
    Span4Mux_v I__4859 (
            .O(N__28937),
            .I(N__28892));
    Span4Mux_v I__4858 (
            .O(N__28934),
            .I(N__28892));
    LocalMux I__4857 (
            .O(N__28931),
            .I(N__28892));
    LocalMux I__4856 (
            .O(N__28916),
            .I(N__28889));
    Span4Mux_h I__4855 (
            .O(N__28913),
            .I(N__28884));
    LocalMux I__4854 (
            .O(N__28910),
            .I(N__28884));
    InMux I__4853 (
            .O(N__28909),
            .I(N__28881));
    CascadeMux I__4852 (
            .O(N__28908),
            .I(N__28877));
    CEMux I__4851 (
            .O(N__28907),
            .I(N__28873));
    InMux I__4850 (
            .O(N__28904),
            .I(N__28870));
    LocalMux I__4849 (
            .O(N__28899),
            .I(N__28867));
    Span4Mux_v I__4848 (
            .O(N__28892),
            .I(N__28860));
    Span4Mux_v I__4847 (
            .O(N__28889),
            .I(N__28860));
    Span4Mux_v I__4846 (
            .O(N__28884),
            .I(N__28855));
    LocalMux I__4845 (
            .O(N__28881),
            .I(N__28855));
    InMux I__4844 (
            .O(N__28880),
            .I(N__28852));
    InMux I__4843 (
            .O(N__28877),
            .I(N__28849));
    InMux I__4842 (
            .O(N__28876),
            .I(N__28846));
    LocalMux I__4841 (
            .O(N__28873),
            .I(N__28841));
    LocalMux I__4840 (
            .O(N__28870),
            .I(N__28841));
    Span4Mux_v I__4839 (
            .O(N__28867),
            .I(N__28838));
    InMux I__4838 (
            .O(N__28866),
            .I(N__28833));
    InMux I__4837 (
            .O(N__28865),
            .I(N__28833));
    Span4Mux_v I__4836 (
            .O(N__28860),
            .I(N__28830));
    Span4Mux_h I__4835 (
            .O(N__28855),
            .I(N__28827));
    LocalMux I__4834 (
            .O(N__28852),
            .I(dds_state_1_adj_1446));
    LocalMux I__4833 (
            .O(N__28849),
            .I(dds_state_1_adj_1446));
    LocalMux I__4832 (
            .O(N__28846),
            .I(dds_state_1_adj_1446));
    Odrv4 I__4831 (
            .O(N__28841),
            .I(dds_state_1_adj_1446));
    Odrv4 I__4830 (
            .O(N__28838),
            .I(dds_state_1_adj_1446));
    LocalMux I__4829 (
            .O(N__28833),
            .I(dds_state_1_adj_1446));
    Odrv4 I__4828 (
            .O(N__28830),
            .I(dds_state_1_adj_1446));
    Odrv4 I__4827 (
            .O(N__28827),
            .I(dds_state_1_adj_1446));
    InMux I__4826 (
            .O(N__28810),
            .I(N__28788));
    InMux I__4825 (
            .O(N__28809),
            .I(N__28788));
    InMux I__4824 (
            .O(N__28808),
            .I(N__28788));
    InMux I__4823 (
            .O(N__28807),
            .I(N__28777));
    InMux I__4822 (
            .O(N__28806),
            .I(N__28777));
    InMux I__4821 (
            .O(N__28805),
            .I(N__28777));
    InMux I__4820 (
            .O(N__28804),
            .I(N__28777));
    InMux I__4819 (
            .O(N__28803),
            .I(N__28777));
    InMux I__4818 (
            .O(N__28802),
            .I(N__28756));
    InMux I__4817 (
            .O(N__28801),
            .I(N__28756));
    InMux I__4816 (
            .O(N__28800),
            .I(N__28756));
    InMux I__4815 (
            .O(N__28799),
            .I(N__28756));
    InMux I__4814 (
            .O(N__28798),
            .I(N__28756));
    InMux I__4813 (
            .O(N__28797),
            .I(N__28756));
    InMux I__4812 (
            .O(N__28796),
            .I(N__28756));
    InMux I__4811 (
            .O(N__28795),
            .I(N__28756));
    LocalMux I__4810 (
            .O(N__28788),
            .I(N__28751));
    LocalMux I__4809 (
            .O(N__28777),
            .I(N__28751));
    InMux I__4808 (
            .O(N__28776),
            .I(N__28743));
    InMux I__4807 (
            .O(N__28775),
            .I(N__28740));
    InMux I__4806 (
            .O(N__28774),
            .I(N__28737));
    InMux I__4805 (
            .O(N__28773),
            .I(N__28733));
    LocalMux I__4804 (
            .O(N__28756),
            .I(N__28728));
    Span4Mux_v I__4803 (
            .O(N__28751),
            .I(N__28728));
    InMux I__4802 (
            .O(N__28750),
            .I(N__28725));
    InMux I__4801 (
            .O(N__28749),
            .I(N__28716));
    InMux I__4800 (
            .O(N__28748),
            .I(N__28716));
    InMux I__4799 (
            .O(N__28747),
            .I(N__28716));
    InMux I__4798 (
            .O(N__28746),
            .I(N__28716));
    LocalMux I__4797 (
            .O(N__28743),
            .I(N__28711));
    LocalMux I__4796 (
            .O(N__28740),
            .I(N__28711));
    LocalMux I__4795 (
            .O(N__28737),
            .I(N__28708));
    InMux I__4794 (
            .O(N__28736),
            .I(N__28705));
    LocalMux I__4793 (
            .O(N__28733),
            .I(N__28702));
    Span4Mux_v I__4792 (
            .O(N__28728),
            .I(N__28699));
    LocalMux I__4791 (
            .O(N__28725),
            .I(N__28694));
    LocalMux I__4790 (
            .O(N__28716),
            .I(N__28694));
    Span4Mux_v I__4789 (
            .O(N__28711),
            .I(N__28689));
    Span4Mux_h I__4788 (
            .O(N__28708),
            .I(N__28689));
    LocalMux I__4787 (
            .O(N__28705),
            .I(dds_state_2_adj_1445));
    Odrv12 I__4786 (
            .O(N__28702),
            .I(dds_state_2_adj_1445));
    Odrv4 I__4785 (
            .O(N__28699),
            .I(dds_state_2_adj_1445));
    Odrv4 I__4784 (
            .O(N__28694),
            .I(dds_state_2_adj_1445));
    Odrv4 I__4783 (
            .O(N__28689),
            .I(dds_state_2_adj_1445));
    CascadeMux I__4782 (
            .O(N__28678),
            .I(N__28674));
    CascadeMux I__4781 (
            .O(N__28677),
            .I(N__28671));
    InMux I__4780 (
            .O(N__28674),
            .I(N__28668));
    InMux I__4779 (
            .O(N__28671),
            .I(N__28665));
    LocalMux I__4778 (
            .O(N__28668),
            .I(N__28661));
    LocalMux I__4777 (
            .O(N__28665),
            .I(N__28658));
    CascadeMux I__4776 (
            .O(N__28664),
            .I(N__28655));
    Span4Mux_h I__4775 (
            .O(N__28661),
            .I(N__28649));
    Span4Mux_v I__4774 (
            .O(N__28658),
            .I(N__28649));
    InMux I__4773 (
            .O(N__28655),
            .I(N__28646));
    CascadeMux I__4772 (
            .O(N__28654),
            .I(N__28643));
    Span4Mux_v I__4771 (
            .O(N__28649),
            .I(N__28640));
    LocalMux I__4770 (
            .O(N__28646),
            .I(N__28637));
    InMux I__4769 (
            .O(N__28643),
            .I(N__28634));
    Span4Mux_v I__4768 (
            .O(N__28640),
            .I(N__28631));
    Span12Mux_h I__4767 (
            .O(N__28637),
            .I(N__28628));
    LocalMux I__4766 (
            .O(N__28634),
            .I(trig_dds1));
    Odrv4 I__4765 (
            .O(N__28631),
            .I(trig_dds1));
    Odrv12 I__4764 (
            .O(N__28628),
            .I(trig_dds1));
    InMux I__4763 (
            .O(N__28621),
            .I(N__28618));
    LocalMux I__4762 (
            .O(N__28618),
            .I(N__28614));
    InMux I__4761 (
            .O(N__28617),
            .I(N__28608));
    Span4Mux_h I__4760 (
            .O(N__28614),
            .I(N__28604));
    InMux I__4759 (
            .O(N__28613),
            .I(N__28601));
    InMux I__4758 (
            .O(N__28612),
            .I(N__28598));
    InMux I__4757 (
            .O(N__28611),
            .I(N__28595));
    LocalMux I__4756 (
            .O(N__28608),
            .I(N__28588));
    InMux I__4755 (
            .O(N__28607),
            .I(N__28585));
    Span4Mux_h I__4754 (
            .O(N__28604),
            .I(N__28582));
    LocalMux I__4753 (
            .O(N__28601),
            .I(N__28575));
    LocalMux I__4752 (
            .O(N__28598),
            .I(N__28575));
    LocalMux I__4751 (
            .O(N__28595),
            .I(N__28575));
    InMux I__4750 (
            .O(N__28594),
            .I(N__28566));
    InMux I__4749 (
            .O(N__28593),
            .I(N__28566));
    InMux I__4748 (
            .O(N__28592),
            .I(N__28566));
    InMux I__4747 (
            .O(N__28591),
            .I(N__28566));
    Odrv4 I__4746 (
            .O(N__28588),
            .I(dds_state_0_adj_1447));
    LocalMux I__4745 (
            .O(N__28585),
            .I(dds_state_0_adj_1447));
    Odrv4 I__4744 (
            .O(N__28582),
            .I(dds_state_0_adj_1447));
    Odrv4 I__4743 (
            .O(N__28575),
            .I(dds_state_0_adj_1447));
    LocalMux I__4742 (
            .O(N__28566),
            .I(dds_state_0_adj_1447));
    CEMux I__4741 (
            .O(N__28555),
            .I(N__28552));
    LocalMux I__4740 (
            .O(N__28552),
            .I(N__28548));
    CEMux I__4739 (
            .O(N__28551),
            .I(N__28545));
    Span4Mux_v I__4738 (
            .O(N__28548),
            .I(N__28540));
    LocalMux I__4737 (
            .O(N__28545),
            .I(N__28540));
    Span4Mux_v I__4736 (
            .O(N__28540),
            .I(N__28537));
    Span4Mux_h I__4735 (
            .O(N__28537),
            .I(N__28534));
    Odrv4 I__4734 (
            .O(N__28534),
            .I(\CLK_DDS.n12722 ));
    InMux I__4733 (
            .O(N__28531),
            .I(N__28527));
    InMux I__4732 (
            .O(N__28530),
            .I(N__28524));
    LocalMux I__4731 (
            .O(N__28527),
            .I(\ADC_VDC.avg_cnt_0 ));
    LocalMux I__4730 (
            .O(N__28524),
            .I(\ADC_VDC.avg_cnt_0 ));
    InMux I__4729 (
            .O(N__28519),
            .I(bfn_11_7_0_));
    CascadeMux I__4728 (
            .O(N__28516),
            .I(N__28512));
    InMux I__4727 (
            .O(N__28515),
            .I(N__28509));
    InMux I__4726 (
            .O(N__28512),
            .I(N__28506));
    LocalMux I__4725 (
            .O(N__28509),
            .I(\ADC_VDC.avg_cnt_1 ));
    LocalMux I__4724 (
            .O(N__28506),
            .I(\ADC_VDC.avg_cnt_1 ));
    InMux I__4723 (
            .O(N__28501),
            .I(\ADC_VDC.n19399 ));
    InMux I__4722 (
            .O(N__28498),
            .I(N__28494));
    InMux I__4721 (
            .O(N__28497),
            .I(N__28491));
    LocalMux I__4720 (
            .O(N__28494),
            .I(\ADC_VDC.avg_cnt_2 ));
    LocalMux I__4719 (
            .O(N__28491),
            .I(\ADC_VDC.avg_cnt_2 ));
    InMux I__4718 (
            .O(N__28486),
            .I(\ADC_VDC.n19400 ));
    CascadeMux I__4717 (
            .O(N__28483),
            .I(N__28479));
    InMux I__4716 (
            .O(N__28482),
            .I(N__28476));
    InMux I__4715 (
            .O(N__28479),
            .I(N__28473));
    LocalMux I__4714 (
            .O(N__28476),
            .I(\ADC_VDC.avg_cnt_3 ));
    LocalMux I__4713 (
            .O(N__28473),
            .I(\ADC_VDC.avg_cnt_3 ));
    InMux I__4712 (
            .O(N__28468),
            .I(\ADC_VDC.n19401 ));
    InMux I__4711 (
            .O(N__28465),
            .I(N__28461));
    InMux I__4710 (
            .O(N__28464),
            .I(N__28458));
    LocalMux I__4709 (
            .O(N__28461),
            .I(\ADC_VDC.avg_cnt_4 ));
    LocalMux I__4708 (
            .O(N__28458),
            .I(\ADC_VDC.avg_cnt_4 ));
    InMux I__4707 (
            .O(N__28453),
            .I(\ADC_VDC.n19402 ));
    InMux I__4706 (
            .O(N__28450),
            .I(N__28446));
    InMux I__4705 (
            .O(N__28449),
            .I(N__28443));
    LocalMux I__4704 (
            .O(N__28446),
            .I(\ADC_VDC.avg_cnt_5 ));
    LocalMux I__4703 (
            .O(N__28443),
            .I(\ADC_VDC.avg_cnt_5 ));
    InMux I__4702 (
            .O(N__28438),
            .I(\ADC_VDC.n19403 ));
    InMux I__4701 (
            .O(N__28435),
            .I(N__28431));
    InMux I__4700 (
            .O(N__28434),
            .I(N__28428));
    LocalMux I__4699 (
            .O(N__28431),
            .I(\ADC_VDC.avg_cnt_6 ));
    LocalMux I__4698 (
            .O(N__28428),
            .I(\ADC_VDC.avg_cnt_6 ));
    InMux I__4697 (
            .O(N__28423),
            .I(\ADC_VDC.n19404 ));
    InMux I__4696 (
            .O(N__28420),
            .I(N__28399));
    InMux I__4695 (
            .O(N__28419),
            .I(N__28399));
    InMux I__4694 (
            .O(N__28418),
            .I(N__28399));
    InMux I__4693 (
            .O(N__28417),
            .I(N__28399));
    InMux I__4692 (
            .O(N__28416),
            .I(N__28399));
    InMux I__4691 (
            .O(N__28415),
            .I(N__28399));
    InMux I__4690 (
            .O(N__28414),
            .I(N__28399));
    LocalMux I__4689 (
            .O(N__28399),
            .I(N__28394));
    CascadeMux I__4688 (
            .O(N__28398),
            .I(N__28391));
    InMux I__4687 (
            .O(N__28397),
            .I(N__28385));
    Span4Mux_v I__4686 (
            .O(N__28394),
            .I(N__28382));
    InMux I__4685 (
            .O(N__28391),
            .I(N__28373));
    InMux I__4684 (
            .O(N__28390),
            .I(N__28373));
    InMux I__4683 (
            .O(N__28389),
            .I(N__28373));
    InMux I__4682 (
            .O(N__28388),
            .I(N__28373));
    LocalMux I__4681 (
            .O(N__28385),
            .I(N__28354));
    Span4Mux_h I__4680 (
            .O(N__28382),
            .I(N__28354));
    LocalMux I__4679 (
            .O(N__28373),
            .I(N__28354));
    InMux I__4678 (
            .O(N__28372),
            .I(N__28337));
    InMux I__4677 (
            .O(N__28371),
            .I(N__28337));
    InMux I__4676 (
            .O(N__28370),
            .I(N__28337));
    InMux I__4675 (
            .O(N__28369),
            .I(N__28337));
    InMux I__4674 (
            .O(N__28368),
            .I(N__28337));
    InMux I__4673 (
            .O(N__28367),
            .I(N__28337));
    InMux I__4672 (
            .O(N__28366),
            .I(N__28337));
    InMux I__4671 (
            .O(N__28365),
            .I(N__28337));
    InMux I__4670 (
            .O(N__28364),
            .I(N__28330));
    InMux I__4669 (
            .O(N__28363),
            .I(N__28330));
    InMux I__4668 (
            .O(N__28362),
            .I(N__28330));
    InMux I__4667 (
            .O(N__28361),
            .I(N__28327));
    Span4Mux_v I__4666 (
            .O(N__28354),
            .I(N__28324));
    LocalMux I__4665 (
            .O(N__28337),
            .I(N__28321));
    LocalMux I__4664 (
            .O(N__28330),
            .I(N__28318));
    LocalMux I__4663 (
            .O(N__28327),
            .I(N__28315));
    Span4Mux_h I__4662 (
            .O(N__28324),
            .I(N__28312));
    Span4Mux_v I__4661 (
            .O(N__28321),
            .I(N__28307));
    Span4Mux_h I__4660 (
            .O(N__28318),
            .I(N__28307));
    Odrv12 I__4659 (
            .O(N__28315),
            .I(n13073));
    Odrv4 I__4658 (
            .O(N__28312),
            .I(n13073));
    Odrv4 I__4657 (
            .O(N__28307),
            .I(n13073));
    CascadeMux I__4656 (
            .O(N__28300),
            .I(\ADC_VDC.n20618_cascade_ ));
    CEMux I__4655 (
            .O(N__28297),
            .I(N__28294));
    LocalMux I__4654 (
            .O(N__28294),
            .I(N__28291));
    Span4Mux_v I__4653 (
            .O(N__28291),
            .I(N__28288));
    Odrv4 I__4652 (
            .O(N__28288),
            .I(\ADC_VDC.n47 ));
    InMux I__4651 (
            .O(N__28285),
            .I(N__28282));
    LocalMux I__4650 (
            .O(N__28282),
            .I(N__28279));
    Odrv4 I__4649 (
            .O(N__28279),
            .I(\ADC_VDC.n20702 ));
    InMux I__4648 (
            .O(N__28276),
            .I(N__28273));
    LocalMux I__4647 (
            .O(N__28273),
            .I(N__28270));
    Span4Mux_v I__4646 (
            .O(N__28270),
            .I(N__28267));
    Odrv4 I__4645 (
            .O(N__28267),
            .I(\ADC_VDC.n20 ));
    InMux I__4644 (
            .O(N__28264),
            .I(\ADC_VDC.genclk.n19416 ));
    InMux I__4643 (
            .O(N__28261),
            .I(bfn_11_4_0_));
    InMux I__4642 (
            .O(N__28258),
            .I(\ADC_VDC.genclk.n19418 ));
    InMux I__4641 (
            .O(N__28255),
            .I(\ADC_VDC.genclk.n19419 ));
    InMux I__4640 (
            .O(N__28252),
            .I(\ADC_VDC.genclk.n19420 ));
    InMux I__4639 (
            .O(N__28249),
            .I(\ADC_VDC.genclk.n19421 ));
    InMux I__4638 (
            .O(N__28246),
            .I(\ADC_VDC.genclk.n19422 ));
    InMux I__4637 (
            .O(N__28243),
            .I(\ADC_VDC.genclk.n19423 ));
    InMux I__4636 (
            .O(N__28240),
            .I(\ADC_VDC.genclk.n19424 ));
    InMux I__4635 (
            .O(N__28237),
            .I(N__28234));
    LocalMux I__4634 (
            .O(N__28234),
            .I(N__28231));
    Span4Mux_h I__4633 (
            .O(N__28231),
            .I(N__28228));
    Odrv4 I__4632 (
            .O(N__28228),
            .I(n16_adj_1489));
    IoInMux I__4631 (
            .O(N__28225),
            .I(N__28222));
    LocalMux I__4630 (
            .O(N__28222),
            .I(N__28219));
    IoSpan4Mux I__4629 (
            .O(N__28219),
            .I(N__28216));
    Span4Mux_s3_v I__4628 (
            .O(N__28216),
            .I(N__28213));
    Span4Mux_v I__4627 (
            .O(N__28213),
            .I(N__28208));
    InMux I__4626 (
            .O(N__28212),
            .I(N__28205));
    InMux I__4625 (
            .O(N__28211),
            .I(N__28202));
    Odrv4 I__4624 (
            .O(N__28208),
            .I(IAC_OSR0));
    LocalMux I__4623 (
            .O(N__28205),
            .I(IAC_OSR0));
    LocalMux I__4622 (
            .O(N__28202),
            .I(IAC_OSR0));
    InMux I__4621 (
            .O(N__28195),
            .I(bfn_11_3_0_));
    InMux I__4620 (
            .O(N__28192),
            .I(\ADC_VDC.genclk.n19410 ));
    InMux I__4619 (
            .O(N__28189),
            .I(\ADC_VDC.genclk.n19411 ));
    InMux I__4618 (
            .O(N__28186),
            .I(\ADC_VDC.genclk.n19412 ));
    InMux I__4617 (
            .O(N__28183),
            .I(\ADC_VDC.genclk.n19413 ));
    InMux I__4616 (
            .O(N__28180),
            .I(\ADC_VDC.genclk.n19414 ));
    InMux I__4615 (
            .O(N__28177),
            .I(\ADC_VDC.genclk.n19415 ));
    InMux I__4614 (
            .O(N__28174),
            .I(N__28171));
    LocalMux I__4613 (
            .O(N__28171),
            .I(N__28168));
    Span4Mux_v I__4612 (
            .O(N__28168),
            .I(N__28165));
    Odrv4 I__4611 (
            .O(N__28165),
            .I(n23_adj_1513));
    CascadeMux I__4610 (
            .O(N__28162),
            .I(N__28158));
    CascadeMux I__4609 (
            .O(N__28161),
            .I(N__28154));
    InMux I__4608 (
            .O(N__28158),
            .I(N__28151));
    InMux I__4607 (
            .O(N__28157),
            .I(N__28146));
    InMux I__4606 (
            .O(N__28154),
            .I(N__28146));
    LocalMux I__4605 (
            .O(N__28151),
            .I(N__28143));
    LocalMux I__4604 (
            .O(N__28146),
            .I(cmd_rdadctmp_28));
    Odrv4 I__4603 (
            .O(N__28143),
            .I(cmd_rdadctmp_28));
    InMux I__4602 (
            .O(N__28138),
            .I(N__28135));
    LocalMux I__4601 (
            .O(N__28135),
            .I(N__28131));
    CascadeMux I__4600 (
            .O(N__28134),
            .I(N__28128));
    Span4Mux_h I__4599 (
            .O(N__28131),
            .I(N__28125));
    InMux I__4598 (
            .O(N__28128),
            .I(N__28122));
    Sp12to4 I__4597 (
            .O(N__28125),
            .I(N__28118));
    LocalMux I__4596 (
            .O(N__28122),
            .I(N__28115));
    InMux I__4595 (
            .O(N__28121),
            .I(N__28112));
    Span12Mux_v I__4594 (
            .O(N__28118),
            .I(N__28109));
    Span4Mux_v I__4593 (
            .O(N__28115),
            .I(N__28106));
    LocalMux I__4592 (
            .O(N__28112),
            .I(buf_adcdata_iac_20));
    Odrv12 I__4591 (
            .O(N__28109),
            .I(buf_adcdata_iac_20));
    Odrv4 I__4590 (
            .O(N__28106),
            .I(buf_adcdata_iac_20));
    IoInMux I__4589 (
            .O(N__28099),
            .I(N__28096));
    LocalMux I__4588 (
            .O(N__28096),
            .I(N__28093));
    IoSpan4Mux I__4587 (
            .O(N__28093),
            .I(N__28090));
    Span4Mux_s0_v I__4586 (
            .O(N__28090),
            .I(N__28087));
    Span4Mux_v I__4585 (
            .O(N__28087),
            .I(N__28082));
    CascadeMux I__4584 (
            .O(N__28086),
            .I(N__28079));
    InMux I__4583 (
            .O(N__28085),
            .I(N__28076));
    Span4Mux_v I__4582 (
            .O(N__28082),
            .I(N__28073));
    InMux I__4581 (
            .O(N__28079),
            .I(N__28070));
    LocalMux I__4580 (
            .O(N__28076),
            .I(N__28067));
    Odrv4 I__4579 (
            .O(N__28073),
            .I(IAC_FLT1));
    LocalMux I__4578 (
            .O(N__28070),
            .I(IAC_FLT1));
    Odrv4 I__4577 (
            .O(N__28067),
            .I(IAC_FLT1));
    IoInMux I__4576 (
            .O(N__28060),
            .I(N__28057));
    LocalMux I__4575 (
            .O(N__28057),
            .I(N__28054));
    Span4Mux_s1_v I__4574 (
            .O(N__28054),
            .I(N__28051));
    Span4Mux_h I__4573 (
            .O(N__28051),
            .I(N__28047));
    InMux I__4572 (
            .O(N__28050),
            .I(N__28043));
    Span4Mux_v I__4571 (
            .O(N__28047),
            .I(N__28040));
    InMux I__4570 (
            .O(N__28046),
            .I(N__28037));
    LocalMux I__4569 (
            .O(N__28043),
            .I(N__28034));
    Odrv4 I__4568 (
            .O(N__28040),
            .I(IAC_OSR1));
    LocalMux I__4567 (
            .O(N__28037),
            .I(IAC_OSR1));
    Odrv4 I__4566 (
            .O(N__28034),
            .I(IAC_OSR1));
    IoInMux I__4565 (
            .O(N__28027),
            .I(N__28024));
    LocalMux I__4564 (
            .O(N__28024),
            .I(N__28021));
    IoSpan4Mux I__4563 (
            .O(N__28021),
            .I(N__28018));
    Span4Mux_s1_v I__4562 (
            .O(N__28018),
            .I(N__28015));
    Span4Mux_v I__4561 (
            .O(N__28015),
            .I(N__28010));
    InMux I__4560 (
            .O(N__28014),
            .I(N__28007));
    InMux I__4559 (
            .O(N__28013),
            .I(N__28004));
    Odrv4 I__4558 (
            .O(N__28010),
            .I(IAC_FLT0));
    LocalMux I__4557 (
            .O(N__28007),
            .I(IAC_FLT0));
    LocalMux I__4556 (
            .O(N__28004),
            .I(IAC_FLT0));
    InMux I__4555 (
            .O(N__27997),
            .I(N__27994));
    LocalMux I__4554 (
            .O(N__27994),
            .I(N__27989));
    CascadeMux I__4553 (
            .O(N__27993),
            .I(N__27986));
    CascadeMux I__4552 (
            .O(N__27992),
            .I(N__27983));
    Span4Mux_v I__4551 (
            .O(N__27989),
            .I(N__27980));
    InMux I__4550 (
            .O(N__27986),
            .I(N__27977));
    InMux I__4549 (
            .O(N__27983),
            .I(N__27974));
    Span4Mux_h I__4548 (
            .O(N__27980),
            .I(N__27971));
    LocalMux I__4547 (
            .O(N__27977),
            .I(buf_adcdata_iac_16));
    LocalMux I__4546 (
            .O(N__27974),
            .I(buf_adcdata_iac_16));
    Odrv4 I__4545 (
            .O(N__27971),
            .I(buf_adcdata_iac_16));
    InMux I__4544 (
            .O(N__27964),
            .I(N__27960));
    InMux I__4543 (
            .O(N__27963),
            .I(N__27956));
    LocalMux I__4542 (
            .O(N__27960),
            .I(N__27953));
    InMux I__4541 (
            .O(N__27959),
            .I(N__27950));
    LocalMux I__4540 (
            .O(N__27956),
            .I(buf_dds1_8));
    Odrv12 I__4539 (
            .O(N__27953),
            .I(buf_dds1_8));
    LocalMux I__4538 (
            .O(N__27950),
            .I(buf_dds1_8));
    CascadeMux I__4537 (
            .O(N__27943),
            .I(n22189_cascade_));
    CascadeMux I__4536 (
            .O(N__27940),
            .I(N__27937));
    InMux I__4535 (
            .O(N__27937),
            .I(N__27934));
    LocalMux I__4534 (
            .O(N__27934),
            .I(N__27931));
    Span4Mux_v I__4533 (
            .O(N__27931),
            .I(N__27928));
    Span4Mux_v I__4532 (
            .O(N__27928),
            .I(N__27925));
    Odrv4 I__4531 (
            .O(N__27925),
            .I(n20769));
    InMux I__4530 (
            .O(N__27922),
            .I(N__27917));
    InMux I__4529 (
            .O(N__27921),
            .I(N__27914));
    InMux I__4528 (
            .O(N__27920),
            .I(N__27911));
    LocalMux I__4527 (
            .O(N__27917),
            .I(N__27908));
    LocalMux I__4526 (
            .O(N__27914),
            .I(buf_dds1_15));
    LocalMux I__4525 (
            .O(N__27911),
            .I(buf_dds1_15));
    Odrv4 I__4524 (
            .O(N__27908),
            .I(buf_dds1_15));
    InMux I__4523 (
            .O(N__27901),
            .I(N__27898));
    LocalMux I__4522 (
            .O(N__27898),
            .I(N__27895));
    Odrv4 I__4521 (
            .O(N__27895),
            .I(n22045));
    InMux I__4520 (
            .O(N__27892),
            .I(N__27889));
    LocalMux I__4519 (
            .O(N__27889),
            .I(N__27886));
    Span4Mux_h I__4518 (
            .O(N__27886),
            .I(N__27883));
    Odrv4 I__4517 (
            .O(N__27883),
            .I(n22048));
    IoInMux I__4516 (
            .O(N__27880),
            .I(N__27877));
    LocalMux I__4515 (
            .O(N__27877),
            .I(N__27874));
    Span4Mux_s1_h I__4514 (
            .O(N__27874),
            .I(N__27870));
    InMux I__4513 (
            .O(N__27873),
            .I(N__27867));
    Sp12to4 I__4512 (
            .O(N__27870),
            .I(N__27864));
    LocalMux I__4511 (
            .O(N__27867),
            .I(N__27861));
    Span12Mux_s5_v I__4510 (
            .O(N__27864),
            .I(N__27858));
    Span4Mux_v I__4509 (
            .O(N__27861),
            .I(N__27854));
    Span12Mux_h I__4508 (
            .O(N__27858),
            .I(N__27851));
    InMux I__4507 (
            .O(N__27857),
            .I(N__27848));
    Span4Mux_h I__4506 (
            .O(N__27854),
            .I(N__27845));
    Odrv12 I__4505 (
            .O(N__27851),
            .I(VAC_FLT0));
    LocalMux I__4504 (
            .O(N__27848),
            .I(VAC_FLT0));
    Odrv4 I__4503 (
            .O(N__27845),
            .I(VAC_FLT0));
    InMux I__4502 (
            .O(N__27838),
            .I(N__27835));
    LocalMux I__4501 (
            .O(N__27835),
            .I(N__27832));
    Span4Mux_h I__4500 (
            .O(N__27832),
            .I(N__27829));
    Odrv4 I__4499 (
            .O(N__27829),
            .I(n16_adj_1480));
    InMux I__4498 (
            .O(N__27826),
            .I(N__27821));
    InMux I__4497 (
            .O(N__27825),
            .I(N__27816));
    InMux I__4496 (
            .O(N__27824),
            .I(N__27816));
    LocalMux I__4495 (
            .O(N__27821),
            .I(buf_dds1_0));
    LocalMux I__4494 (
            .O(N__27816),
            .I(buf_dds1_0));
    InMux I__4493 (
            .O(N__27811),
            .I(N__27808));
    LocalMux I__4492 (
            .O(N__27808),
            .I(N__27805));
    Span4Mux_h I__4491 (
            .O(N__27805),
            .I(N__27802));
    Span4Mux_v I__4490 (
            .O(N__27802),
            .I(N__27797));
    CascadeMux I__4489 (
            .O(N__27801),
            .I(N__27794));
    InMux I__4488 (
            .O(N__27800),
            .I(N__27791));
    Span4Mux_v I__4487 (
            .O(N__27797),
            .I(N__27788));
    InMux I__4486 (
            .O(N__27794),
            .I(N__27785));
    LocalMux I__4485 (
            .O(N__27791),
            .I(buf_adcdata_iac_18));
    Odrv4 I__4484 (
            .O(N__27788),
            .I(buf_adcdata_iac_18));
    LocalMux I__4483 (
            .O(N__27785),
            .I(buf_adcdata_iac_18));
    CascadeMux I__4482 (
            .O(N__27778),
            .I(N__27774));
    InMux I__4481 (
            .O(N__27777),
            .I(N__27770));
    InMux I__4480 (
            .O(N__27774),
            .I(N__27767));
    InMux I__4479 (
            .O(N__27773),
            .I(N__27764));
    LocalMux I__4478 (
            .O(N__27770),
            .I(cmd_rdadctmp_25));
    LocalMux I__4477 (
            .O(N__27767),
            .I(cmd_rdadctmp_25));
    LocalMux I__4476 (
            .O(N__27764),
            .I(cmd_rdadctmp_25));
    InMux I__4475 (
            .O(N__27757),
            .I(N__27753));
    CascadeMux I__4474 (
            .O(N__27756),
            .I(N__27750));
    LocalMux I__4473 (
            .O(N__27753),
            .I(N__27747));
    InMux I__4472 (
            .O(N__27750),
            .I(N__27743));
    Span4Mux_h I__4471 (
            .O(N__27747),
            .I(N__27740));
    InMux I__4470 (
            .O(N__27746),
            .I(N__27737));
    LocalMux I__4469 (
            .O(N__27743),
            .I(cmd_rdadctmp_26));
    Odrv4 I__4468 (
            .O(N__27740),
            .I(cmd_rdadctmp_26));
    LocalMux I__4467 (
            .O(N__27737),
            .I(cmd_rdadctmp_26));
    CascadeMux I__4466 (
            .O(N__27730),
            .I(N__27727));
    InMux I__4465 (
            .O(N__27727),
            .I(N__27723));
    InMux I__4464 (
            .O(N__27726),
            .I(N__27720));
    LocalMux I__4463 (
            .O(N__27723),
            .I(N__27717));
    LocalMux I__4462 (
            .O(N__27720),
            .I(N__27714));
    Span4Mux_v I__4461 (
            .O(N__27717),
            .I(N__27709));
    Span4Mux_h I__4460 (
            .O(N__27714),
            .I(N__27709));
    Odrv4 I__4459 (
            .O(N__27709),
            .I(tmp_buf_15_adj_1448));
    CascadeMux I__4458 (
            .O(N__27706),
            .I(N__27703));
    InMux I__4457 (
            .O(N__27703),
            .I(N__27700));
    LocalMux I__4456 (
            .O(N__27700),
            .I(\CLK_DDS.tmp_buf_0 ));
    CascadeMux I__4455 (
            .O(N__27697),
            .I(N__27694));
    InMux I__4454 (
            .O(N__27694),
            .I(N__27691));
    LocalMux I__4453 (
            .O(N__27691),
            .I(\CLK_DDS.tmp_buf_1 ));
    CascadeMux I__4452 (
            .O(N__27688),
            .I(N__27685));
    InMux I__4451 (
            .O(N__27685),
            .I(N__27682));
    LocalMux I__4450 (
            .O(N__27682),
            .I(\CLK_DDS.tmp_buf_2 ));
    CascadeMux I__4449 (
            .O(N__27679),
            .I(N__27676));
    InMux I__4448 (
            .O(N__27676),
            .I(N__27673));
    LocalMux I__4447 (
            .O(N__27673),
            .I(N__27670));
    Odrv4 I__4446 (
            .O(N__27670),
            .I(\CLK_DDS.tmp_buf_3 ));
    CascadeMux I__4445 (
            .O(N__27667),
            .I(N__27664));
    InMux I__4444 (
            .O(N__27664),
            .I(N__27661));
    LocalMux I__4443 (
            .O(N__27661),
            .I(\CLK_DDS.tmp_buf_4 ));
    CascadeMux I__4442 (
            .O(N__27658),
            .I(N__27655));
    InMux I__4441 (
            .O(N__27655),
            .I(N__27652));
    LocalMux I__4440 (
            .O(N__27652),
            .I(\CLK_DDS.tmp_buf_5 ));
    CascadeMux I__4439 (
            .O(N__27649),
            .I(N__27646));
    InMux I__4438 (
            .O(N__27646),
            .I(N__27643));
    LocalMux I__4437 (
            .O(N__27643),
            .I(\CLK_DDS.tmp_buf_6 ));
    CascadeMux I__4436 (
            .O(N__27640),
            .I(N__27637));
    InMux I__4435 (
            .O(N__27637),
            .I(N__27634));
    LocalMux I__4434 (
            .O(N__27634),
            .I(N__27631));
    Odrv12 I__4433 (
            .O(N__27631),
            .I(\CLK_DDS.tmp_buf_7 ));
    CascadeMux I__4432 (
            .O(N__27628),
            .I(N__27625));
    InMux I__4431 (
            .O(N__27625),
            .I(N__27622));
    LocalMux I__4430 (
            .O(N__27622),
            .I(\CLK_DDS.tmp_buf_9 ));
    InMux I__4429 (
            .O(N__27619),
            .I(N__27616));
    LocalMux I__4428 (
            .O(N__27616),
            .I(\CLK_DDS.tmp_buf_8 ));
    InMux I__4427 (
            .O(N__27613),
            .I(N__27610));
    LocalMux I__4426 (
            .O(N__27610),
            .I(N__27605));
    InMux I__4425 (
            .O(N__27609),
            .I(N__27602));
    InMux I__4424 (
            .O(N__27608),
            .I(N__27599));
    Span4Mux_v I__4423 (
            .O(N__27605),
            .I(N__27596));
    LocalMux I__4422 (
            .O(N__27602),
            .I(buf_dds1_14));
    LocalMux I__4421 (
            .O(N__27599),
            .I(buf_dds1_14));
    Odrv4 I__4420 (
            .O(N__27596),
            .I(buf_dds1_14));
    InMux I__4419 (
            .O(N__27589),
            .I(N__27584));
    InMux I__4418 (
            .O(N__27588),
            .I(N__27581));
    InMux I__4417 (
            .O(N__27587),
            .I(N__27578));
    LocalMux I__4416 (
            .O(N__27584),
            .I(buf_dds1_12));
    LocalMux I__4415 (
            .O(N__27581),
            .I(buf_dds1_12));
    LocalMux I__4414 (
            .O(N__27578),
            .I(buf_dds1_12));
    InMux I__4413 (
            .O(N__27571),
            .I(N__27567));
    CascadeMux I__4412 (
            .O(N__27570),
            .I(N__27563));
    LocalMux I__4411 (
            .O(N__27567),
            .I(N__27560));
    InMux I__4410 (
            .O(N__27566),
            .I(N__27557));
    InMux I__4409 (
            .O(N__27563),
            .I(N__27554));
    Span4Mux_h I__4408 (
            .O(N__27560),
            .I(N__27551));
    LocalMux I__4407 (
            .O(N__27557),
            .I(buf_dds1_9));
    LocalMux I__4406 (
            .O(N__27554),
            .I(buf_dds1_9));
    Odrv4 I__4405 (
            .O(N__27551),
            .I(buf_dds1_9));
    CascadeMux I__4404 (
            .O(N__27544),
            .I(n22036_cascade_));
    InMux I__4403 (
            .O(N__27541),
            .I(N__27538));
    LocalMux I__4402 (
            .O(N__27538),
            .I(N__27535));
    Span4Mux_h I__4401 (
            .O(N__27535),
            .I(N__27532));
    Odrv4 I__4400 (
            .O(N__27532),
            .I(n22156));
    InMux I__4399 (
            .O(N__27529),
            .I(N__27526));
    LocalMux I__4398 (
            .O(N__27526),
            .I(n21910));
    CascadeMux I__4397 (
            .O(N__27523),
            .I(n20823_cascade_));
    CascadeMux I__4396 (
            .O(N__27520),
            .I(n30_adj_1514_cascade_));
    CEMux I__4395 (
            .O(N__27517),
            .I(N__27514));
    LocalMux I__4394 (
            .O(N__27514),
            .I(N__27509));
    CEMux I__4393 (
            .O(N__27513),
            .I(N__27506));
    CEMux I__4392 (
            .O(N__27512),
            .I(N__27501));
    Span4Mux_h I__4391 (
            .O(N__27509),
            .I(N__27496));
    LocalMux I__4390 (
            .O(N__27506),
            .I(N__27496));
    CEMux I__4389 (
            .O(N__27505),
            .I(N__27493));
    CEMux I__4388 (
            .O(N__27504),
            .I(N__27490));
    LocalMux I__4387 (
            .O(N__27501),
            .I(N__27487));
    Span4Mux_h I__4386 (
            .O(N__27496),
            .I(N__27484));
    LocalMux I__4385 (
            .O(N__27493),
            .I(N__27481));
    LocalMux I__4384 (
            .O(N__27490),
            .I(N__27478));
    Odrv4 I__4383 (
            .O(N__27487),
            .I(n11941));
    Odrv4 I__4382 (
            .O(N__27484),
            .I(n11941));
    Odrv12 I__4381 (
            .O(N__27481),
            .I(n11941));
    Odrv12 I__4380 (
            .O(N__27478),
            .I(n11941));
    SRMux I__4379 (
            .O(N__27469),
            .I(N__27466));
    LocalMux I__4378 (
            .O(N__27466),
            .I(N__27461));
    SRMux I__4377 (
            .O(N__27465),
            .I(N__27458));
    SRMux I__4376 (
            .O(N__27464),
            .I(N__27455));
    Span4Mux_v I__4375 (
            .O(N__27461),
            .I(N__27448));
    LocalMux I__4374 (
            .O(N__27458),
            .I(N__27448));
    LocalMux I__4373 (
            .O(N__27455),
            .I(N__27445));
    SRMux I__4372 (
            .O(N__27454),
            .I(N__27442));
    SRMux I__4371 (
            .O(N__27453),
            .I(N__27439));
    Span4Mux_h I__4370 (
            .O(N__27448),
            .I(N__27436));
    Span4Mux_h I__4369 (
            .O(N__27445),
            .I(N__27433));
    LocalMux I__4368 (
            .O(N__27442),
            .I(N__27430));
    LocalMux I__4367 (
            .O(N__27439),
            .I(N__27427));
    Odrv4 I__4366 (
            .O(N__27436),
            .I(n14735));
    Odrv4 I__4365 (
            .O(N__27433),
            .I(n14735));
    Odrv12 I__4364 (
            .O(N__27430),
            .I(n14735));
    Odrv12 I__4363 (
            .O(N__27427),
            .I(n14735));
    CascadeMux I__4362 (
            .O(N__27418),
            .I(N__27415));
    InMux I__4361 (
            .O(N__27415),
            .I(N__27412));
    LocalMux I__4360 (
            .O(N__27412),
            .I(\CLK_DDS.tmp_buf_10 ));
    CascadeMux I__4359 (
            .O(N__27409),
            .I(N__27406));
    InMux I__4358 (
            .O(N__27406),
            .I(N__27403));
    LocalMux I__4357 (
            .O(N__27403),
            .I(\CLK_DDS.tmp_buf_11 ));
    CascadeMux I__4356 (
            .O(N__27400),
            .I(N__27397));
    InMux I__4355 (
            .O(N__27397),
            .I(N__27394));
    LocalMux I__4354 (
            .O(N__27394),
            .I(\CLK_DDS.tmp_buf_12 ));
    CascadeMux I__4353 (
            .O(N__27391),
            .I(N__27388));
    InMux I__4352 (
            .O(N__27388),
            .I(N__27385));
    LocalMux I__4351 (
            .O(N__27385),
            .I(\CLK_DDS.tmp_buf_13 ));
    CascadeMux I__4350 (
            .O(N__27382),
            .I(N__27379));
    InMux I__4349 (
            .O(N__27379),
            .I(N__27376));
    LocalMux I__4348 (
            .O(N__27376),
            .I(\CLK_DDS.tmp_buf_14 ));
    InMux I__4347 (
            .O(N__27373),
            .I(N__27370));
    LocalMux I__4346 (
            .O(N__27370),
            .I(N__27367));
    Span4Mux_h I__4345 (
            .O(N__27367),
            .I(N__27364));
    Span4Mux_h I__4344 (
            .O(N__27364),
            .I(N__27361));
    Odrv4 I__4343 (
            .O(N__27361),
            .I(buf_data_iac_18));
    CascadeMux I__4342 (
            .O(N__27358),
            .I(n20794_cascade_));
    InMux I__4341 (
            .O(N__27355),
            .I(N__27352));
    LocalMux I__4340 (
            .O(N__27352),
            .I(n21922));
    CascadeMux I__4339 (
            .O(N__27349),
            .I(n20796_cascade_));
    InMux I__4338 (
            .O(N__27346),
            .I(N__27343));
    LocalMux I__4337 (
            .O(N__27343),
            .I(N__27340));
    Span4Mux_h I__4336 (
            .O(N__27340),
            .I(N__27337));
    Odrv4 I__4335 (
            .O(N__27337),
            .I(n21934));
    CascadeMux I__4334 (
            .O(N__27334),
            .I(n22213_cascade_));
    CascadeMux I__4333 (
            .O(N__27331),
            .I(n22216_cascade_));
    InMux I__4332 (
            .O(N__27328),
            .I(N__27325));
    LocalMux I__4331 (
            .O(N__27325),
            .I(N__27322));
    Span4Mux_h I__4330 (
            .O(N__27322),
            .I(N__27319));
    Span4Mux_h I__4329 (
            .O(N__27319),
            .I(N__27316));
    Odrv4 I__4328 (
            .O(N__27316),
            .I(n20937));
    CascadeMux I__4327 (
            .O(N__27313),
            .I(N__27310));
    InMux I__4326 (
            .O(N__27310),
            .I(N__27307));
    LocalMux I__4325 (
            .O(N__27307),
            .I(n20936));
    CascadeMux I__4324 (
            .O(N__27304),
            .I(n21907_cascade_));
    InMux I__4323 (
            .O(N__27301),
            .I(N__27297));
    CascadeMux I__4322 (
            .O(N__27300),
            .I(N__27294));
    LocalMux I__4321 (
            .O(N__27297),
            .I(N__27291));
    InMux I__4320 (
            .O(N__27294),
            .I(N__27288));
    Span12Mux_h I__4319 (
            .O(N__27291),
            .I(N__27284));
    LocalMux I__4318 (
            .O(N__27288),
            .I(N__27281));
    InMux I__4317 (
            .O(N__27287),
            .I(N__27278));
    Span12Mux_v I__4316 (
            .O(N__27284),
            .I(N__27275));
    Span4Mux_h I__4315 (
            .O(N__27281),
            .I(N__27272));
    LocalMux I__4314 (
            .O(N__27278),
            .I(buf_adcdata_iac_21));
    Odrv12 I__4313 (
            .O(N__27275),
            .I(buf_adcdata_iac_21));
    Odrv4 I__4312 (
            .O(N__27272),
            .I(buf_adcdata_iac_21));
    CascadeMux I__4311 (
            .O(N__27265),
            .I(n22033_cascade_));
    CascadeMux I__4310 (
            .O(N__27262),
            .I(n12_cascade_));
    CEMux I__4309 (
            .O(N__27259),
            .I(N__27256));
    LocalMux I__4308 (
            .O(N__27256),
            .I(n12116));
    CascadeMux I__4307 (
            .O(N__27253),
            .I(n12116_cascade_));
    SRMux I__4306 (
            .O(N__27250),
            .I(N__27247));
    LocalMux I__4305 (
            .O(N__27247),
            .I(N__27244));
    Span4Mux_h I__4304 (
            .O(N__27244),
            .I(N__27241));
    Odrv4 I__4303 (
            .O(N__27241),
            .I(n14756));
    CascadeMux I__4302 (
            .O(N__27238),
            .I(n25_adj_1592_cascade_));
    CascadeMux I__4301 (
            .O(N__27235),
            .I(n11944_cascade_));
    CascadeMux I__4300 (
            .O(N__27232),
            .I(n11941_cascade_));
    CascadeMux I__4299 (
            .O(N__27229),
            .I(n21919_cascade_));
    InMux I__4298 (
            .O(N__27226),
            .I(N__27223));
    LocalMux I__4297 (
            .O(N__27223),
            .I(N__27220));
    Span4Mux_h I__4296 (
            .O(N__27220),
            .I(N__27217));
    Span4Mux_v I__4295 (
            .O(N__27217),
            .I(N__27214));
    Span4Mux_v I__4294 (
            .O(N__27214),
            .I(N__27211));
    Odrv4 I__4293 (
            .O(N__27211),
            .I(buf_data_vac_23));
    InMux I__4292 (
            .O(N__27208),
            .I(N__27205));
    LocalMux I__4291 (
            .O(N__27205),
            .I(N__27202));
    Span4Mux_h I__4290 (
            .O(N__27202),
            .I(N__27199));
    Span4Mux_h I__4289 (
            .O(N__27199),
            .I(N__27196));
    Span4Mux_v I__4288 (
            .O(N__27196),
            .I(N__27193));
    Odrv4 I__4287 (
            .O(N__27193),
            .I(buf_data_vac_22));
    CascadeMux I__4286 (
            .O(N__27190),
            .I(N__27187));
    InMux I__4285 (
            .O(N__27187),
            .I(N__27184));
    LocalMux I__4284 (
            .O(N__27184),
            .I(N__27181));
    Span12Mux_h I__4283 (
            .O(N__27181),
            .I(N__27178));
    Odrv12 I__4282 (
            .O(N__27178),
            .I(buf_data_vac_21));
    InMux I__4281 (
            .O(N__27175),
            .I(N__27172));
    LocalMux I__4280 (
            .O(N__27172),
            .I(N__27169));
    Span4Mux_h I__4279 (
            .O(N__27169),
            .I(N__27166));
    Span4Mux_h I__4278 (
            .O(N__27166),
            .I(N__27163));
    Span4Mux_v I__4277 (
            .O(N__27163),
            .I(N__27160));
    Odrv4 I__4276 (
            .O(N__27160),
            .I(buf_data_vac_20));
    InMux I__4275 (
            .O(N__27157),
            .I(N__27154));
    LocalMux I__4274 (
            .O(N__27154),
            .I(N__27151));
    Odrv12 I__4273 (
            .O(N__27151),
            .I(buf_data_vac_19));
    InMux I__4272 (
            .O(N__27148),
            .I(N__27145));
    LocalMux I__4271 (
            .O(N__27145),
            .I(N__27142));
    Span4Mux_h I__4270 (
            .O(N__27142),
            .I(N__27139));
    Span4Mux_h I__4269 (
            .O(N__27139),
            .I(N__27136));
    Odrv4 I__4268 (
            .O(N__27136),
            .I(buf_data_vac_18));
    InMux I__4267 (
            .O(N__27133),
            .I(N__27130));
    LocalMux I__4266 (
            .O(N__27130),
            .I(N__27127));
    Span4Mux_v I__4265 (
            .O(N__27127),
            .I(N__27124));
    Span4Mux_h I__4264 (
            .O(N__27124),
            .I(N__27121));
    Odrv4 I__4263 (
            .O(N__27121),
            .I(buf_data_vac_17));
    CascadeMux I__4262 (
            .O(N__27118),
            .I(n21143_cascade_));
    InMux I__4261 (
            .O(N__27115),
            .I(N__27111));
    InMux I__4260 (
            .O(N__27114),
            .I(N__27108));
    LocalMux I__4259 (
            .O(N__27111),
            .I(cmd_rdadcbuf_18));
    LocalMux I__4258 (
            .O(N__27108),
            .I(cmd_rdadcbuf_18));
    InMux I__4257 (
            .O(N__27103),
            .I(N__27099));
    InMux I__4256 (
            .O(N__27102),
            .I(N__27096));
    LocalMux I__4255 (
            .O(N__27099),
            .I(cmd_rdadcbuf_17));
    LocalMux I__4254 (
            .O(N__27096),
            .I(cmd_rdadcbuf_17));
    CascadeMux I__4253 (
            .O(N__27091),
            .I(N__27088));
    InMux I__4252 (
            .O(N__27088),
            .I(N__27084));
    InMux I__4251 (
            .O(N__27087),
            .I(N__27081));
    LocalMux I__4250 (
            .O(N__27084),
            .I(cmd_rdadcbuf_16));
    LocalMux I__4249 (
            .O(N__27081),
            .I(cmd_rdadcbuf_16));
    InMux I__4248 (
            .O(N__27076),
            .I(N__27073));
    LocalMux I__4247 (
            .O(N__27073),
            .I(N__27070));
    Odrv12 I__4246 (
            .O(N__27070),
            .I(\ADC_VDC.n18394 ));
    InMux I__4245 (
            .O(N__27067),
            .I(N__27064));
    LocalMux I__4244 (
            .O(N__27064),
            .I(N__27061));
    Odrv4 I__4243 (
            .O(N__27061),
            .I(\ADC_VDC.cmd_rdadcbuf_35_N_1130_34 ));
    CascadeMux I__4242 (
            .O(N__27058),
            .I(\ADC_VDC.n21106_cascade_ ));
    InMux I__4241 (
            .O(N__27055),
            .I(N__27052));
    LocalMux I__4240 (
            .O(N__27052),
            .I(N__27049));
    Span4Mux_h I__4239 (
            .O(N__27049),
            .I(N__27044));
    InMux I__4238 (
            .O(N__27048),
            .I(N__27041));
    InMux I__4237 (
            .O(N__27047),
            .I(N__27038));
    Odrv4 I__4236 (
            .O(N__27044),
            .I(cmd_rdadcbuf_34));
    LocalMux I__4235 (
            .O(N__27041),
            .I(cmd_rdadcbuf_34));
    LocalMux I__4234 (
            .O(N__27038),
            .I(cmd_rdadcbuf_34));
    CEMux I__4233 (
            .O(N__27031),
            .I(N__27028));
    LocalMux I__4232 (
            .O(N__27028),
            .I(N__27025));
    Odrv4 I__4231 (
            .O(N__27025),
            .I(\ADC_VDC.n13020 ));
    InMux I__4230 (
            .O(N__27022),
            .I(N__27019));
    LocalMux I__4229 (
            .O(N__27019),
            .I(N__27016));
    Odrv12 I__4228 (
            .O(N__27016),
            .I(\ADC_VDC.n21 ));
    InMux I__4227 (
            .O(N__27013),
            .I(N__27010));
    LocalMux I__4226 (
            .O(N__27010),
            .I(N__27007));
    Odrv12 I__4225 (
            .O(N__27007),
            .I(\ADC_VDC.n19 ));
    InMux I__4224 (
            .O(N__27004),
            .I(N__27001));
    LocalMux I__4223 (
            .O(N__27001),
            .I(N__26998));
    Span4Mux_h I__4222 (
            .O(N__26998),
            .I(N__26995));
    Span4Mux_h I__4221 (
            .O(N__26995),
            .I(N__26992));
    Odrv4 I__4220 (
            .O(N__26992),
            .I(buf_data_vac_16));
    InMux I__4219 (
            .O(N__26989),
            .I(N__26985));
    CascadeMux I__4218 (
            .O(N__26988),
            .I(N__26981));
    LocalMux I__4217 (
            .O(N__26985),
            .I(N__26978));
    CascadeMux I__4216 (
            .O(N__26984),
            .I(N__26975));
    InMux I__4215 (
            .O(N__26981),
            .I(N__26972));
    Span4Mux_h I__4214 (
            .O(N__26978),
            .I(N__26969));
    InMux I__4213 (
            .O(N__26975),
            .I(N__26966));
    LocalMux I__4212 (
            .O(N__26972),
            .I(cmd_rdadctmp_10_adj_1462));
    Odrv4 I__4211 (
            .O(N__26969),
            .I(cmd_rdadctmp_10_adj_1462));
    LocalMux I__4210 (
            .O(N__26966),
            .I(cmd_rdadctmp_10_adj_1462));
    CascadeMux I__4209 (
            .O(N__26959),
            .I(N__26954));
    InMux I__4208 (
            .O(N__26958),
            .I(N__26949));
    InMux I__4207 (
            .O(N__26957),
            .I(N__26949));
    InMux I__4206 (
            .O(N__26954),
            .I(N__26946));
    LocalMux I__4205 (
            .O(N__26949),
            .I(cmd_rdadctmp_11_adj_1461));
    LocalMux I__4204 (
            .O(N__26946),
            .I(cmd_rdadctmp_11_adj_1461));
    CascadeMux I__4203 (
            .O(N__26941),
            .I(\ADC_VDC.n21673_cascade_ ));
    IoInMux I__4202 (
            .O(N__26938),
            .I(N__26935));
    LocalMux I__4201 (
            .O(N__26935),
            .I(N__26932));
    Span12Mux_s11_h I__4200 (
            .O(N__26932),
            .I(N__26928));
    InMux I__4199 (
            .O(N__26931),
            .I(N__26925));
    Odrv12 I__4198 (
            .O(N__26928),
            .I(VDC_SCLK));
    LocalMux I__4197 (
            .O(N__26925),
            .I(VDC_SCLK));
    InMux I__4196 (
            .O(N__26920),
            .I(N__26916));
    CascadeMux I__4195 (
            .O(N__26919),
            .I(N__26912));
    LocalMux I__4194 (
            .O(N__26916),
            .I(N__26909));
    InMux I__4193 (
            .O(N__26915),
            .I(N__26906));
    InMux I__4192 (
            .O(N__26912),
            .I(N__26903));
    Odrv4 I__4191 (
            .O(N__26909),
            .I(cmd_rdadctmp_19_adj_1453));
    LocalMux I__4190 (
            .O(N__26906),
            .I(cmd_rdadctmp_19_adj_1453));
    LocalMux I__4189 (
            .O(N__26903),
            .I(cmd_rdadctmp_19_adj_1453));
    CascadeMux I__4188 (
            .O(N__26896),
            .I(N__26892));
    CascadeMux I__4187 (
            .O(N__26895),
            .I(N__26885));
    InMux I__4186 (
            .O(N__26892),
            .I(N__26875));
    InMux I__4185 (
            .O(N__26891),
            .I(N__26864));
    InMux I__4184 (
            .O(N__26890),
            .I(N__26864));
    InMux I__4183 (
            .O(N__26889),
            .I(N__26864));
    InMux I__4182 (
            .O(N__26888),
            .I(N__26864));
    InMux I__4181 (
            .O(N__26885),
            .I(N__26864));
    CascadeMux I__4180 (
            .O(N__26884),
            .I(N__26861));
    CascadeMux I__4179 (
            .O(N__26883),
            .I(N__26858));
    CascadeMux I__4178 (
            .O(N__26882),
            .I(N__26855));
    CascadeMux I__4177 (
            .O(N__26881),
            .I(N__26852));
    CascadeMux I__4176 (
            .O(N__26880),
            .I(N__26847));
    CascadeMux I__4175 (
            .O(N__26879),
            .I(N__26843));
    CascadeMux I__4174 (
            .O(N__26878),
            .I(N__26838));
    LocalMux I__4173 (
            .O(N__26875),
            .I(N__26831));
    LocalMux I__4172 (
            .O(N__26864),
            .I(N__26831));
    InMux I__4171 (
            .O(N__26861),
            .I(N__26818));
    InMux I__4170 (
            .O(N__26858),
            .I(N__26818));
    InMux I__4169 (
            .O(N__26855),
            .I(N__26818));
    InMux I__4168 (
            .O(N__26852),
            .I(N__26818));
    InMux I__4167 (
            .O(N__26851),
            .I(N__26818));
    InMux I__4166 (
            .O(N__26850),
            .I(N__26818));
    InMux I__4165 (
            .O(N__26847),
            .I(N__26805));
    InMux I__4164 (
            .O(N__26846),
            .I(N__26805));
    InMux I__4163 (
            .O(N__26843),
            .I(N__26805));
    InMux I__4162 (
            .O(N__26842),
            .I(N__26805));
    InMux I__4161 (
            .O(N__26841),
            .I(N__26805));
    InMux I__4160 (
            .O(N__26838),
            .I(N__26805));
    CascadeMux I__4159 (
            .O(N__26837),
            .I(N__26802));
    CascadeMux I__4158 (
            .O(N__26836),
            .I(N__26799));
    Span4Mux_v I__4157 (
            .O(N__26831),
            .I(N__26792));
    LocalMux I__4156 (
            .O(N__26818),
            .I(N__26792));
    LocalMux I__4155 (
            .O(N__26805),
            .I(N__26789));
    InMux I__4154 (
            .O(N__26802),
            .I(N__26780));
    InMux I__4153 (
            .O(N__26799),
            .I(N__26780));
    InMux I__4152 (
            .O(N__26798),
            .I(N__26780));
    InMux I__4151 (
            .O(N__26797),
            .I(N__26780));
    Odrv4 I__4150 (
            .O(N__26792),
            .I(n12853));
    Odrv4 I__4149 (
            .O(N__26789),
            .I(n12853));
    LocalMux I__4148 (
            .O(N__26780),
            .I(n12853));
    CascadeMux I__4147 (
            .O(N__26773),
            .I(N__26770));
    InMux I__4146 (
            .O(N__26770),
            .I(N__26765));
    CascadeMux I__4145 (
            .O(N__26769),
            .I(N__26762));
    InMux I__4144 (
            .O(N__26768),
            .I(N__26759));
    LocalMux I__4143 (
            .O(N__26765),
            .I(N__26756));
    InMux I__4142 (
            .O(N__26762),
            .I(N__26753));
    LocalMux I__4141 (
            .O(N__26759),
            .I(cmd_rdadctmp_20_adj_1452));
    Odrv12 I__4140 (
            .O(N__26756),
            .I(cmd_rdadctmp_20_adj_1452));
    LocalMux I__4139 (
            .O(N__26753),
            .I(cmd_rdadctmp_20_adj_1452));
    InMux I__4138 (
            .O(N__26746),
            .I(N__26742));
    InMux I__4137 (
            .O(N__26745),
            .I(N__26739));
    LocalMux I__4136 (
            .O(N__26742),
            .I(cmd_rdadcbuf_23));
    LocalMux I__4135 (
            .O(N__26739),
            .I(cmd_rdadcbuf_23));
    InMux I__4134 (
            .O(N__26734),
            .I(N__26731));
    LocalMux I__4133 (
            .O(N__26731),
            .I(N__26728));
    Span4Mux_v I__4132 (
            .O(N__26728),
            .I(N__26724));
    CascadeMux I__4131 (
            .O(N__26727),
            .I(N__26721));
    Span4Mux_v I__4130 (
            .O(N__26724),
            .I(N__26718));
    InMux I__4129 (
            .O(N__26721),
            .I(N__26715));
    Odrv4 I__4128 (
            .O(N__26718),
            .I(buf_adcdata_vdc_12));
    LocalMux I__4127 (
            .O(N__26715),
            .I(buf_adcdata_vdc_12));
    InMux I__4126 (
            .O(N__26710),
            .I(N__26706));
    InMux I__4125 (
            .O(N__26709),
            .I(N__26703));
    LocalMux I__4124 (
            .O(N__26706),
            .I(cmd_rdadcbuf_22));
    LocalMux I__4123 (
            .O(N__26703),
            .I(cmd_rdadcbuf_22));
    InMux I__4122 (
            .O(N__26698),
            .I(N__26695));
    LocalMux I__4121 (
            .O(N__26695),
            .I(N__26692));
    Span4Mux_v I__4120 (
            .O(N__26692),
            .I(N__26688));
    CascadeMux I__4119 (
            .O(N__26691),
            .I(N__26685));
    Span4Mux_v I__4118 (
            .O(N__26688),
            .I(N__26682));
    InMux I__4117 (
            .O(N__26685),
            .I(N__26679));
    Odrv4 I__4116 (
            .O(N__26682),
            .I(buf_adcdata_vdc_11));
    LocalMux I__4115 (
            .O(N__26679),
            .I(buf_adcdata_vdc_11));
    CascadeMux I__4114 (
            .O(N__26674),
            .I(N__26671));
    InMux I__4113 (
            .O(N__26671),
            .I(N__26667));
    InMux I__4112 (
            .O(N__26670),
            .I(N__26664));
    LocalMux I__4111 (
            .O(N__26667),
            .I(cmd_rdadcbuf_15));
    LocalMux I__4110 (
            .O(N__26664),
            .I(cmd_rdadcbuf_15));
    InMux I__4109 (
            .O(N__26659),
            .I(N__26655));
    InMux I__4108 (
            .O(N__26658),
            .I(N__26652));
    LocalMux I__4107 (
            .O(N__26655),
            .I(cmd_rdadcbuf_20));
    LocalMux I__4106 (
            .O(N__26652),
            .I(cmd_rdadcbuf_20));
    InMux I__4105 (
            .O(N__26647),
            .I(N__26643));
    InMux I__4104 (
            .O(N__26646),
            .I(N__26640));
    LocalMux I__4103 (
            .O(N__26643),
            .I(cmd_rdadcbuf_19));
    LocalMux I__4102 (
            .O(N__26640),
            .I(cmd_rdadcbuf_19));
    InMux I__4101 (
            .O(N__26635),
            .I(N__26632));
    LocalMux I__4100 (
            .O(N__26632),
            .I(N__26629));
    Span4Mux_h I__4099 (
            .O(N__26629),
            .I(N__26625));
    CascadeMux I__4098 (
            .O(N__26628),
            .I(N__26622));
    Span4Mux_v I__4097 (
            .O(N__26625),
            .I(N__26619));
    InMux I__4096 (
            .O(N__26622),
            .I(N__26616));
    Odrv4 I__4095 (
            .O(N__26619),
            .I(buf_adcdata_vdc_8));
    LocalMux I__4094 (
            .O(N__26616),
            .I(buf_adcdata_vdc_8));
    CascadeMux I__4093 (
            .O(N__26611),
            .I(N__26606));
    InMux I__4092 (
            .O(N__26610),
            .I(N__26603));
    InMux I__4091 (
            .O(N__26609),
            .I(N__26600));
    InMux I__4090 (
            .O(N__26606),
            .I(N__26597));
    LocalMux I__4089 (
            .O(N__26603),
            .I(cmd_rdadctmp_0_adj_1472));
    LocalMux I__4088 (
            .O(N__26600),
            .I(cmd_rdadctmp_0_adj_1472));
    LocalMux I__4087 (
            .O(N__26597),
            .I(cmd_rdadctmp_0_adj_1472));
    CascadeMux I__4086 (
            .O(N__26590),
            .I(N__26587));
    InMux I__4085 (
            .O(N__26587),
            .I(N__26582));
    InMux I__4084 (
            .O(N__26586),
            .I(N__26577));
    InMux I__4083 (
            .O(N__26585),
            .I(N__26577));
    LocalMux I__4082 (
            .O(N__26582),
            .I(N__26574));
    LocalMux I__4081 (
            .O(N__26577),
            .I(cmd_rdadctmp_3_adj_1469));
    Odrv4 I__4080 (
            .O(N__26574),
            .I(cmd_rdadctmp_3_adj_1469));
    InMux I__4079 (
            .O(N__26569),
            .I(N__26565));
    CascadeMux I__4078 (
            .O(N__26568),
            .I(N__26561));
    LocalMux I__4077 (
            .O(N__26565),
            .I(N__26558));
    InMux I__4076 (
            .O(N__26564),
            .I(N__26555));
    InMux I__4075 (
            .O(N__26561),
            .I(N__26552));
    Odrv4 I__4074 (
            .O(N__26558),
            .I(cmd_rdadctmp_4_adj_1468));
    LocalMux I__4073 (
            .O(N__26555),
            .I(cmd_rdadctmp_4_adj_1468));
    LocalMux I__4072 (
            .O(N__26552),
            .I(cmd_rdadctmp_4_adj_1468));
    CEMux I__4071 (
            .O(N__26545),
            .I(N__26542));
    LocalMux I__4070 (
            .O(N__26542),
            .I(N__26539));
    Span4Mux_h I__4069 (
            .O(N__26539),
            .I(N__26536));
    Odrv4 I__4068 (
            .O(N__26536),
            .I(\ADC_VDC.n12885 ));
    CascadeMux I__4067 (
            .O(N__26533),
            .I(N__26529));
    InMux I__4066 (
            .O(N__26532),
            .I(N__26525));
    InMux I__4065 (
            .O(N__26529),
            .I(N__26522));
    InMux I__4064 (
            .O(N__26528),
            .I(N__26519));
    LocalMux I__4063 (
            .O(N__26525),
            .I(N__26514));
    LocalMux I__4062 (
            .O(N__26522),
            .I(N__26514));
    LocalMux I__4061 (
            .O(N__26519),
            .I(cmd_rdadctmp_7_adj_1465));
    Odrv4 I__4060 (
            .O(N__26514),
            .I(cmd_rdadctmp_7_adj_1465));
    InMux I__4059 (
            .O(N__26509),
            .I(N__26505));
    CascadeMux I__4058 (
            .O(N__26508),
            .I(N__26501));
    LocalMux I__4057 (
            .O(N__26505),
            .I(N__26498));
    InMux I__4056 (
            .O(N__26504),
            .I(N__26495));
    InMux I__4055 (
            .O(N__26501),
            .I(N__26492));
    Odrv4 I__4054 (
            .O(N__26498),
            .I(cmd_rdadctmp_8_adj_1464));
    LocalMux I__4053 (
            .O(N__26495),
            .I(cmd_rdadctmp_8_adj_1464));
    LocalMux I__4052 (
            .O(N__26492),
            .I(cmd_rdadctmp_8_adj_1464));
    CascadeMux I__4051 (
            .O(N__26485),
            .I(N__26482));
    InMux I__4050 (
            .O(N__26482),
            .I(N__26477));
    CascadeMux I__4049 (
            .O(N__26481),
            .I(N__26474));
    InMux I__4048 (
            .O(N__26480),
            .I(N__26471));
    LocalMux I__4047 (
            .O(N__26477),
            .I(N__26468));
    InMux I__4046 (
            .O(N__26474),
            .I(N__26465));
    LocalMux I__4045 (
            .O(N__26471),
            .I(cmd_rdadctmp_17_adj_1455));
    Odrv12 I__4044 (
            .O(N__26468),
            .I(cmd_rdadctmp_17_adj_1455));
    LocalMux I__4043 (
            .O(N__26465),
            .I(cmd_rdadctmp_17_adj_1455));
    CascadeMux I__4042 (
            .O(N__26458),
            .I(N__26455));
    InMux I__4041 (
            .O(N__26455),
            .I(N__26452));
    LocalMux I__4040 (
            .O(N__26452),
            .I(N__26447));
    CascadeMux I__4039 (
            .O(N__26451),
            .I(N__26444));
    InMux I__4038 (
            .O(N__26450),
            .I(N__26441));
    Span4Mux_h I__4037 (
            .O(N__26447),
            .I(N__26438));
    InMux I__4036 (
            .O(N__26444),
            .I(N__26435));
    LocalMux I__4035 (
            .O(N__26441),
            .I(cmd_rdadctmp_15_adj_1457));
    Odrv4 I__4034 (
            .O(N__26438),
            .I(cmd_rdadctmp_15_adj_1457));
    LocalMux I__4033 (
            .O(N__26435),
            .I(cmd_rdadctmp_15_adj_1457));
    CascadeMux I__4032 (
            .O(N__26428),
            .I(N__26423));
    InMux I__4031 (
            .O(N__26427),
            .I(N__26418));
    InMux I__4030 (
            .O(N__26426),
            .I(N__26418));
    InMux I__4029 (
            .O(N__26423),
            .I(N__26415));
    LocalMux I__4028 (
            .O(N__26418),
            .I(cmd_rdadctmp_16_adj_1456));
    LocalMux I__4027 (
            .O(N__26415),
            .I(cmd_rdadctmp_16_adj_1456));
    CascadeMux I__4026 (
            .O(N__26410),
            .I(N__26405));
    InMux I__4025 (
            .O(N__26409),
            .I(N__26402));
    InMux I__4024 (
            .O(N__26408),
            .I(N__26399));
    InMux I__4023 (
            .O(N__26405),
            .I(N__26396));
    LocalMux I__4022 (
            .O(N__26402),
            .I(cmd_rdadctmp_1_adj_1471));
    LocalMux I__4021 (
            .O(N__26399),
            .I(cmd_rdadctmp_1_adj_1471));
    LocalMux I__4020 (
            .O(N__26396),
            .I(cmd_rdadctmp_1_adj_1471));
    CascadeMux I__4019 (
            .O(N__26389),
            .I(N__26384));
    InMux I__4018 (
            .O(N__26388),
            .I(N__26381));
    InMux I__4017 (
            .O(N__26387),
            .I(N__26378));
    InMux I__4016 (
            .O(N__26384),
            .I(N__26375));
    LocalMux I__4015 (
            .O(N__26381),
            .I(N__26372));
    LocalMux I__4014 (
            .O(N__26378),
            .I(cmd_rdadctmp_2_adj_1470));
    LocalMux I__4013 (
            .O(N__26375),
            .I(cmd_rdadctmp_2_adj_1470));
    Odrv4 I__4012 (
            .O(N__26372),
            .I(cmd_rdadctmp_2_adj_1470));
    CascadeMux I__4011 (
            .O(N__26365),
            .I(N__26360));
    CascadeMux I__4010 (
            .O(N__26364),
            .I(N__26357));
    InMux I__4009 (
            .O(N__26363),
            .I(N__26354));
    InMux I__4008 (
            .O(N__26360),
            .I(N__26351));
    InMux I__4007 (
            .O(N__26357),
            .I(N__26348));
    LocalMux I__4006 (
            .O(N__26354),
            .I(N__26345));
    LocalMux I__4005 (
            .O(N__26351),
            .I(N__26342));
    LocalMux I__4004 (
            .O(N__26348),
            .I(cmd_rdadctmp_12_adj_1460));
    Odrv4 I__4003 (
            .O(N__26345),
            .I(cmd_rdadctmp_12_adj_1460));
    Odrv4 I__4002 (
            .O(N__26342),
            .I(cmd_rdadctmp_12_adj_1460));
    CascadeMux I__4001 (
            .O(N__26335),
            .I(\ADC_VDC.n31_cascade_ ));
    CascadeMux I__4000 (
            .O(N__26332),
            .I(\ADC_VDC.n21925_cascade_ ));
    InMux I__3999 (
            .O(N__26329),
            .I(N__26326));
    LocalMux I__3998 (
            .O(N__26326),
            .I(\ADC_VDC.n18397 ));
    CascadeMux I__3997 (
            .O(N__26323),
            .I(\ADC_VDC.n21928_cascade_ ));
    CEMux I__3996 (
            .O(N__26320),
            .I(N__26317));
    LocalMux I__3995 (
            .O(N__26317),
            .I(N__26314));
    Odrv4 I__3994 (
            .O(N__26314),
            .I(\ADC_VDC.n20514 ));
    CascadeMux I__3993 (
            .O(N__26311),
            .I(\ADC_VDC.n6_cascade_ ));
    InMux I__3992 (
            .O(N__26308),
            .I(N__26304));
    InMux I__3991 (
            .O(N__26307),
            .I(N__26301));
    LocalMux I__3990 (
            .O(N__26304),
            .I(\ADC_VDC.n10519 ));
    LocalMux I__3989 (
            .O(N__26301),
            .I(\ADC_VDC.n10519 ));
    CascadeMux I__3988 (
            .O(N__26296),
            .I(n12853_cascade_));
    CascadeMux I__3987 (
            .O(N__26293),
            .I(N__26289));
    CascadeMux I__3986 (
            .O(N__26292),
            .I(N__26286));
    InMux I__3985 (
            .O(N__26289),
            .I(N__26283));
    InMux I__3984 (
            .O(N__26286),
            .I(N__26280));
    LocalMux I__3983 (
            .O(N__26283),
            .I(cmd_rdadctmp_31));
    LocalMux I__3982 (
            .O(N__26280),
            .I(cmd_rdadctmp_31));
    InMux I__3981 (
            .O(N__26275),
            .I(N__26272));
    LocalMux I__3980 (
            .O(N__26272),
            .I(N__26269));
    Span4Mux_v I__3979 (
            .O(N__26269),
            .I(N__26266));
    Span4Mux_v I__3978 (
            .O(N__26266),
            .I(N__26263));
    Span4Mux_h I__3977 (
            .O(N__26263),
            .I(N__26259));
    CascadeMux I__3976 (
            .O(N__26262),
            .I(N__26255));
    Sp12to4 I__3975 (
            .O(N__26259),
            .I(N__26252));
    InMux I__3974 (
            .O(N__26258),
            .I(N__26247));
    InMux I__3973 (
            .O(N__26255),
            .I(N__26247));
    Odrv12 I__3972 (
            .O(N__26252),
            .I(buf_adcdata_iac_23));
    LocalMux I__3971 (
            .O(N__26247),
            .I(buf_adcdata_iac_23));
    IoInMux I__3970 (
            .O(N__26242),
            .I(N__26239));
    LocalMux I__3969 (
            .O(N__26239),
            .I(N__26236));
    Span4Mux_s0_v I__3968 (
            .O(N__26236),
            .I(N__26233));
    Span4Mux_v I__3967 (
            .O(N__26233),
            .I(N__26230));
    Span4Mux_v I__3966 (
            .O(N__26230),
            .I(N__26227));
    Sp12to4 I__3965 (
            .O(N__26227),
            .I(N__26224));
    Odrv12 I__3964 (
            .O(N__26224),
            .I(AC_ADC_SYNC));
    IoInMux I__3963 (
            .O(N__26221),
            .I(N__26218));
    LocalMux I__3962 (
            .O(N__26218),
            .I(N__26215));
    Span4Mux_s3_h I__3961 (
            .O(N__26215),
            .I(N__26212));
    Span4Mux_v I__3960 (
            .O(N__26212),
            .I(N__26209));
    Sp12to4 I__3959 (
            .O(N__26209),
            .I(N__26204));
    InMux I__3958 (
            .O(N__26208),
            .I(N__26199));
    InMux I__3957 (
            .O(N__26207),
            .I(N__26199));
    Odrv12 I__3956 (
            .O(N__26204),
            .I(VAC_FLT1));
    LocalMux I__3955 (
            .O(N__26199),
            .I(VAC_FLT1));
    IoInMux I__3954 (
            .O(N__26194),
            .I(N__26191));
    LocalMux I__3953 (
            .O(N__26191),
            .I(N__26188));
    Span4Mux_s3_v I__3952 (
            .O(N__26188),
            .I(N__26185));
    Span4Mux_h I__3951 (
            .O(N__26185),
            .I(N__26181));
    CascadeMux I__3950 (
            .O(N__26184),
            .I(N__26178));
    Span4Mux_v I__3949 (
            .O(N__26181),
            .I(N__26175));
    InMux I__3948 (
            .O(N__26178),
            .I(N__26172));
    Odrv4 I__3947 (
            .O(N__26175),
            .I(IAC_SCLK));
    LocalMux I__3946 (
            .O(N__26172),
            .I(IAC_SCLK));
    CascadeMux I__3945 (
            .O(N__26167),
            .I(\ADC_VDC.n18394_cascade_ ));
    InMux I__3944 (
            .O(N__26164),
            .I(N__26161));
    LocalMux I__3943 (
            .O(N__26161),
            .I(N__26158));
    Sp12to4 I__3942 (
            .O(N__26158),
            .I(N__26155));
    Odrv12 I__3941 (
            .O(N__26155),
            .I(EIS_SYNCCLK));
    IoInMux I__3940 (
            .O(N__26152),
            .I(N__26149));
    LocalMux I__3939 (
            .O(N__26149),
            .I(N__26145));
    IoInMux I__3938 (
            .O(N__26148),
            .I(N__26142));
    Span4Mux_s3_v I__3937 (
            .O(N__26145),
            .I(N__26139));
    LocalMux I__3936 (
            .O(N__26142),
            .I(N__26136));
    Span4Mux_h I__3935 (
            .O(N__26139),
            .I(N__26133));
    Span4Mux_s3_h I__3934 (
            .O(N__26136),
            .I(N__26130));
    Sp12to4 I__3933 (
            .O(N__26133),
            .I(N__26127));
    Span4Mux_v I__3932 (
            .O(N__26130),
            .I(N__26124));
    Span12Mux_s11_v I__3931 (
            .O(N__26127),
            .I(N__26119));
    Sp12to4 I__3930 (
            .O(N__26124),
            .I(N__26119));
    Span12Mux_v I__3929 (
            .O(N__26119),
            .I(N__26116));
    Odrv12 I__3928 (
            .O(N__26116),
            .I(IAC_CLK));
    IoInMux I__3927 (
            .O(N__26113),
            .I(N__26110));
    LocalMux I__3926 (
            .O(N__26110),
            .I(N__26107));
    Span4Mux_s3_h I__3925 (
            .O(N__26107),
            .I(N__26104));
    Span4Mux_v I__3924 (
            .O(N__26104),
            .I(N__26101));
    Span4Mux_v I__3923 (
            .O(N__26101),
            .I(N__26097));
    InMux I__3922 (
            .O(N__26100),
            .I(N__26093));
    Sp12to4 I__3921 (
            .O(N__26097),
            .I(N__26090));
    InMux I__3920 (
            .O(N__26096),
            .I(N__26087));
    LocalMux I__3919 (
            .O(N__26093),
            .I(N__26084));
    Odrv12 I__3918 (
            .O(N__26090),
            .I(VAC_OSR0));
    LocalMux I__3917 (
            .O(N__26087),
            .I(VAC_OSR0));
    Odrv4 I__3916 (
            .O(N__26084),
            .I(VAC_OSR0));
    InMux I__3915 (
            .O(N__26077),
            .I(N__26074));
    LocalMux I__3914 (
            .O(N__26074),
            .I(N__26071));
    Span4Mux_h I__3913 (
            .O(N__26071),
            .I(N__26066));
    CascadeMux I__3912 (
            .O(N__26070),
            .I(N__26063));
    InMux I__3911 (
            .O(N__26069),
            .I(N__26060));
    Span4Mux_v I__3910 (
            .O(N__26066),
            .I(N__26057));
    InMux I__3909 (
            .O(N__26063),
            .I(N__26054));
    LocalMux I__3908 (
            .O(N__26060),
            .I(buf_adcdata_iac_19));
    Odrv4 I__3907 (
            .O(N__26057),
            .I(buf_adcdata_iac_19));
    LocalMux I__3906 (
            .O(N__26054),
            .I(buf_adcdata_iac_19));
    InMux I__3905 (
            .O(N__26047),
            .I(N__26044));
    LocalMux I__3904 (
            .O(N__26044),
            .I(N__26041));
    Odrv12 I__3903 (
            .O(N__26041),
            .I(n11417));
    InMux I__3902 (
            .O(N__26038),
            .I(N__26035));
    LocalMux I__3901 (
            .O(N__26035),
            .I(N__26032));
    Span4Mux_v I__3900 (
            .O(N__26032),
            .I(N__26028));
    CascadeMux I__3899 (
            .O(N__26031),
            .I(N__26024));
    Span4Mux_h I__3898 (
            .O(N__26028),
            .I(N__26021));
    InMux I__3897 (
            .O(N__26027),
            .I(N__26016));
    InMux I__3896 (
            .O(N__26024),
            .I(N__26016));
    Odrv4 I__3895 (
            .O(N__26021),
            .I(buf_adcdata_iac_17));
    LocalMux I__3894 (
            .O(N__26016),
            .I(buf_adcdata_iac_17));
    CascadeMux I__3893 (
            .O(N__26011),
            .I(n22201_cascade_));
    CascadeMux I__3892 (
            .O(N__26008),
            .I(N__26005));
    InMux I__3891 (
            .O(N__26005),
            .I(N__26002));
    LocalMux I__3890 (
            .O(N__26002),
            .I(N__25999));
    Span4Mux_v I__3889 (
            .O(N__25999),
            .I(N__25996));
    Odrv4 I__3888 (
            .O(N__25996),
            .I(n20805));
    CascadeMux I__3887 (
            .O(N__25993),
            .I(N__25989));
    InMux I__3886 (
            .O(N__25992),
            .I(N__25986));
    InMux I__3885 (
            .O(N__25989),
            .I(N__25983));
    LocalMux I__3884 (
            .O(N__25986),
            .I(N__25977));
    LocalMux I__3883 (
            .O(N__25983),
            .I(N__25977));
    InMux I__3882 (
            .O(N__25982),
            .I(N__25974));
    Odrv12 I__3881 (
            .O(N__25977),
            .I(cmd_rdadctmp_24));
    LocalMux I__3880 (
            .O(N__25974),
            .I(cmd_rdadctmp_24));
    InMux I__3879 (
            .O(N__25969),
            .I(N__25965));
    InMux I__3878 (
            .O(N__25968),
            .I(N__25962));
    LocalMux I__3877 (
            .O(N__25965),
            .I(N__25958));
    LocalMux I__3876 (
            .O(N__25962),
            .I(N__25955));
    InMux I__3875 (
            .O(N__25961),
            .I(N__25952));
    Span4Mux_v I__3874 (
            .O(N__25958),
            .I(N__25949));
    Span4Mux_h I__3873 (
            .O(N__25955),
            .I(N__25946));
    LocalMux I__3872 (
            .O(N__25952),
            .I(buf_adcdata_iac_10));
    Odrv4 I__3871 (
            .O(N__25949),
            .I(buf_adcdata_iac_10));
    Odrv4 I__3870 (
            .O(N__25946),
            .I(buf_adcdata_iac_10));
    CascadeMux I__3869 (
            .O(N__25939),
            .I(N__25934));
    CascadeMux I__3868 (
            .O(N__25938),
            .I(N__25931));
    CascadeMux I__3867 (
            .O(N__25937),
            .I(N__25927));
    InMux I__3866 (
            .O(N__25934),
            .I(N__25920));
    InMux I__3865 (
            .O(N__25931),
            .I(N__25920));
    InMux I__3864 (
            .O(N__25930),
            .I(N__25920));
    InMux I__3863 (
            .O(N__25927),
            .I(N__25917));
    LocalMux I__3862 (
            .O(N__25920),
            .I(\SIG_DDS.bit_cnt_1 ));
    LocalMux I__3861 (
            .O(N__25917),
            .I(\SIG_DDS.bit_cnt_1 ));
    InMux I__3860 (
            .O(N__25912),
            .I(N__25905));
    InMux I__3859 (
            .O(N__25911),
            .I(N__25905));
    InMux I__3858 (
            .O(N__25910),
            .I(N__25902));
    LocalMux I__3857 (
            .O(N__25905),
            .I(\SIG_DDS.bit_cnt_2 ));
    LocalMux I__3856 (
            .O(N__25902),
            .I(\SIG_DDS.bit_cnt_2 ));
    InMux I__3855 (
            .O(N__25897),
            .I(N__25894));
    LocalMux I__3854 (
            .O(N__25894),
            .I(N__25890));
    InMux I__3853 (
            .O(N__25893),
            .I(N__25886));
    Span12Mux_v I__3852 (
            .O(N__25890),
            .I(N__25883));
    InMux I__3851 (
            .O(N__25889),
            .I(N__25880));
    LocalMux I__3850 (
            .O(N__25886),
            .I(buf_adcdata_vac_11));
    Odrv12 I__3849 (
            .O(N__25883),
            .I(buf_adcdata_vac_11));
    LocalMux I__3848 (
            .O(N__25880),
            .I(buf_adcdata_vac_11));
    CascadeMux I__3847 (
            .O(N__25873),
            .I(N__25869));
    CascadeMux I__3846 (
            .O(N__25872),
            .I(N__25866));
    InMux I__3845 (
            .O(N__25869),
            .I(N__25863));
    InMux I__3844 (
            .O(N__25866),
            .I(N__25860));
    LocalMux I__3843 (
            .O(N__25863),
            .I(N__25857));
    LocalMux I__3842 (
            .O(N__25860),
            .I(N__25853));
    Span4Mux_h I__3841 (
            .O(N__25857),
            .I(N__25850));
    InMux I__3840 (
            .O(N__25856),
            .I(N__25847));
    Odrv4 I__3839 (
            .O(N__25853),
            .I(cmd_rdadctmp_23));
    Odrv4 I__3838 (
            .O(N__25850),
            .I(cmd_rdadctmp_23));
    LocalMux I__3837 (
            .O(N__25847),
            .I(cmd_rdadctmp_23));
    CascadeMux I__3836 (
            .O(N__25840),
            .I(N__25837));
    InMux I__3835 (
            .O(N__25837),
            .I(N__25834));
    LocalMux I__3834 (
            .O(N__25834),
            .I(n8));
    InMux I__3833 (
            .O(N__25831),
            .I(N__25828));
    LocalMux I__3832 (
            .O(N__25828),
            .I(N__25825));
    Span4Mux_h I__3831 (
            .O(N__25825),
            .I(N__25822));
    Odrv4 I__3830 (
            .O(N__25822),
            .I(n22117));
    CascadeMux I__3829 (
            .O(N__25819),
            .I(N__25816));
    InMux I__3828 (
            .O(N__25816),
            .I(N__25813));
    LocalMux I__3827 (
            .O(N__25813),
            .I(N__25809));
    InMux I__3826 (
            .O(N__25812),
            .I(N__25805));
    Span4Mux_h I__3825 (
            .O(N__25809),
            .I(N__25802));
    InMux I__3824 (
            .O(N__25808),
            .I(N__25799));
    LocalMux I__3823 (
            .O(N__25805),
            .I(N__25796));
    Span4Mux_h I__3822 (
            .O(N__25802),
            .I(N__25793));
    LocalMux I__3821 (
            .O(N__25799),
            .I(buf_adcdata_iac_13));
    Odrv4 I__3820 (
            .O(N__25796),
            .I(buf_adcdata_iac_13));
    Odrv4 I__3819 (
            .O(N__25793),
            .I(buf_adcdata_iac_13));
    InMux I__3818 (
            .O(N__25786),
            .I(N__25782));
    InMux I__3817 (
            .O(N__25785),
            .I(N__25779));
    LocalMux I__3816 (
            .O(N__25782),
            .I(\SIG_DDS.bit_cnt_3 ));
    LocalMux I__3815 (
            .O(N__25779),
            .I(\SIG_DDS.bit_cnt_3 ));
    InMux I__3814 (
            .O(N__25774),
            .I(N__25771));
    LocalMux I__3813 (
            .O(N__25771),
            .I(N__25768));
    Odrv12 I__3812 (
            .O(N__25768),
            .I(\SIG_DDS.n21292 ));
    CascadeMux I__3811 (
            .O(N__25765),
            .I(n20624_cascade_));
    CascadeMux I__3810 (
            .O(N__25762),
            .I(\SIG_DDS.n10_cascade_ ));
    CascadeMux I__3809 (
            .O(N__25759),
            .I(N__25756));
    InMux I__3808 (
            .O(N__25756),
            .I(N__25753));
    LocalMux I__3807 (
            .O(N__25753),
            .I(N__25750));
    Span4Mux_v I__3806 (
            .O(N__25750),
            .I(N__25747));
    Span4Mux_h I__3805 (
            .O(N__25747),
            .I(N__25743));
    CascadeMux I__3804 (
            .O(N__25746),
            .I(N__25740));
    Span4Mux_v I__3803 (
            .O(N__25743),
            .I(N__25737));
    InMux I__3802 (
            .O(N__25740),
            .I(N__25734));
    Odrv4 I__3801 (
            .O(N__25737),
            .I(buf_readRTD_12));
    LocalMux I__3800 (
            .O(N__25734),
            .I(buf_readRTD_12));
    InMux I__3799 (
            .O(N__25729),
            .I(N__25726));
    LocalMux I__3798 (
            .O(N__25726),
            .I(n22006));
    CascadeMux I__3797 (
            .O(N__25723),
            .I(n22027_cascade_));
    InMux I__3796 (
            .O(N__25720),
            .I(N__25717));
    LocalMux I__3795 (
            .O(N__25717),
            .I(N__25714));
    Odrv4 I__3794 (
            .O(N__25714),
            .I(n22030));
    InMux I__3793 (
            .O(N__25711),
            .I(N__25707));
    InMux I__3792 (
            .O(N__25710),
            .I(N__25703));
    LocalMux I__3791 (
            .O(N__25707),
            .I(N__25700));
    CascadeMux I__3790 (
            .O(N__25706),
            .I(N__25697));
    LocalMux I__3789 (
            .O(N__25703),
            .I(N__25694));
    Span4Mux_v I__3788 (
            .O(N__25700),
            .I(N__25691));
    InMux I__3787 (
            .O(N__25697),
            .I(N__25688));
    Span4Mux_h I__3786 (
            .O(N__25694),
            .I(N__25685));
    Span4Mux_v I__3785 (
            .O(N__25691),
            .I(N__25682));
    LocalMux I__3784 (
            .O(N__25688),
            .I(buf_adcdata_vac_20));
    Odrv4 I__3783 (
            .O(N__25685),
            .I(buf_adcdata_vac_20));
    Odrv4 I__3782 (
            .O(N__25682),
            .I(buf_adcdata_vac_20));
    CascadeMux I__3781 (
            .O(N__25675),
            .I(N__25672));
    InMux I__3780 (
            .O(N__25672),
            .I(N__25669));
    LocalMux I__3779 (
            .O(N__25669),
            .I(N__25665));
    CascadeMux I__3778 (
            .O(N__25668),
            .I(N__25662));
    Span4Mux_v I__3777 (
            .O(N__25665),
            .I(N__25659));
    InMux I__3776 (
            .O(N__25662),
            .I(N__25656));
    Odrv4 I__3775 (
            .O(N__25659),
            .I(buf_adcdata_vdc_20));
    LocalMux I__3774 (
            .O(N__25656),
            .I(buf_adcdata_vdc_20));
    InMux I__3773 (
            .O(N__25651),
            .I(N__25648));
    LocalMux I__3772 (
            .O(N__25648),
            .I(n22207));
    InMux I__3771 (
            .O(N__25645),
            .I(N__25642));
    LocalMux I__3770 (
            .O(N__25642),
            .I(n20801));
    InMux I__3769 (
            .O(N__25639),
            .I(N__25636));
    LocalMux I__3768 (
            .O(N__25636),
            .I(N__25633));
    Span4Mux_h I__3767 (
            .O(N__25633),
            .I(N__25630));
    Span4Mux_h I__3766 (
            .O(N__25630),
            .I(N__25627));
    Odrv4 I__3765 (
            .O(N__25627),
            .I(buf_data_iac_17));
    CascadeMux I__3764 (
            .O(N__25624),
            .I(n20818_cascade_));
    InMux I__3763 (
            .O(N__25621),
            .I(N__25618));
    LocalMux I__3762 (
            .O(N__25618),
            .I(n20871));
    CascadeMux I__3761 (
            .O(N__25615),
            .I(n20820_cascade_));
    InMux I__3760 (
            .O(N__25612),
            .I(N__25609));
    LocalMux I__3759 (
            .O(N__25609),
            .I(n21967));
    InMux I__3758 (
            .O(N__25606),
            .I(N__25603));
    LocalMux I__3757 (
            .O(N__25603),
            .I(n21970));
    CascadeMux I__3756 (
            .O(N__25600),
            .I(n22003_cascade_));
    InMux I__3755 (
            .O(N__25597),
            .I(N__25594));
    LocalMux I__3754 (
            .O(N__25594),
            .I(N__25591));
    Odrv4 I__3753 (
            .O(N__25591),
            .I(n22060));
    InMux I__3752 (
            .O(N__25588),
            .I(N__25585));
    LocalMux I__3751 (
            .O(N__25585),
            .I(n22054));
    CascadeMux I__3750 (
            .O(N__25582),
            .I(n22015_cascade_));
    InMux I__3749 (
            .O(N__25579),
            .I(N__25575));
    InMux I__3748 (
            .O(N__25578),
            .I(N__25572));
    LocalMux I__3747 (
            .O(N__25575),
            .I(cmd_rdadcbuf_28));
    LocalMux I__3746 (
            .O(N__25572),
            .I(cmd_rdadcbuf_28));
    InMux I__3745 (
            .O(N__25567),
            .I(\ADC_VDC.n19391 ));
    InMux I__3744 (
            .O(N__25564),
            .I(N__25560));
    InMux I__3743 (
            .O(N__25563),
            .I(N__25557));
    LocalMux I__3742 (
            .O(N__25560),
            .I(cmd_rdadcbuf_29));
    LocalMux I__3741 (
            .O(N__25557),
            .I(cmd_rdadcbuf_29));
    InMux I__3740 (
            .O(N__25552),
            .I(\ADC_VDC.n19392 ));
    InMux I__3739 (
            .O(N__25549),
            .I(N__25545));
    InMux I__3738 (
            .O(N__25548),
            .I(N__25542));
    LocalMux I__3737 (
            .O(N__25545),
            .I(cmd_rdadcbuf_30));
    LocalMux I__3736 (
            .O(N__25542),
            .I(cmd_rdadcbuf_30));
    InMux I__3735 (
            .O(N__25537),
            .I(\ADC_VDC.n19393 ));
    InMux I__3734 (
            .O(N__25534),
            .I(N__25530));
    InMux I__3733 (
            .O(N__25533),
            .I(N__25527));
    LocalMux I__3732 (
            .O(N__25530),
            .I(cmd_rdadcbuf_31));
    LocalMux I__3731 (
            .O(N__25527),
            .I(cmd_rdadcbuf_31));
    InMux I__3730 (
            .O(N__25522),
            .I(\ADC_VDC.n19394 ));
    InMux I__3729 (
            .O(N__25519),
            .I(N__25515));
    InMux I__3728 (
            .O(N__25518),
            .I(N__25512));
    LocalMux I__3727 (
            .O(N__25515),
            .I(cmd_rdadcbuf_32));
    LocalMux I__3726 (
            .O(N__25512),
            .I(cmd_rdadcbuf_32));
    InMux I__3725 (
            .O(N__25507),
            .I(bfn_9_9_0_));
    InMux I__3724 (
            .O(N__25504),
            .I(N__25500));
    InMux I__3723 (
            .O(N__25503),
            .I(N__25497));
    LocalMux I__3722 (
            .O(N__25500),
            .I(cmd_rdadcbuf_33));
    LocalMux I__3721 (
            .O(N__25497),
            .I(cmd_rdadcbuf_33));
    InMux I__3720 (
            .O(N__25492),
            .I(\ADC_VDC.n19396 ));
    InMux I__3719 (
            .O(N__25489),
            .I(\ADC_VDC.n19397 ));
    InMux I__3718 (
            .O(N__25486),
            .I(N__25483));
    LocalMux I__3717 (
            .O(N__25483),
            .I(N__25480));
    Odrv4 I__3716 (
            .O(N__25480),
            .I(n20772));
    InMux I__3715 (
            .O(N__25477),
            .I(N__25474));
    LocalMux I__3714 (
            .O(N__25474),
            .I(n21943));
    CascadeMux I__3713 (
            .O(N__25471),
            .I(n21946_cascade_));
    InMux I__3712 (
            .O(N__25468),
            .I(\ADC_VDC.n19383 ));
    CascadeMux I__3711 (
            .O(N__25465),
            .I(N__25460));
    InMux I__3710 (
            .O(N__25464),
            .I(N__25457));
    InMux I__3709 (
            .O(N__25463),
            .I(N__25454));
    InMux I__3708 (
            .O(N__25460),
            .I(N__25451));
    LocalMux I__3707 (
            .O(N__25457),
            .I(cmd_rdadctmp_21_adj_1451));
    LocalMux I__3706 (
            .O(N__25454),
            .I(cmd_rdadctmp_21_adj_1451));
    LocalMux I__3705 (
            .O(N__25451),
            .I(cmd_rdadctmp_21_adj_1451));
    InMux I__3704 (
            .O(N__25444),
            .I(N__25440));
    InMux I__3703 (
            .O(N__25443),
            .I(N__25437));
    LocalMux I__3702 (
            .O(N__25440),
            .I(cmd_rdadcbuf_21));
    LocalMux I__3701 (
            .O(N__25437),
            .I(cmd_rdadcbuf_21));
    InMux I__3700 (
            .O(N__25432),
            .I(\ADC_VDC.n19384 ));
    InMux I__3699 (
            .O(N__25429),
            .I(N__25425));
    CascadeMux I__3698 (
            .O(N__25428),
            .I(N__25421));
    LocalMux I__3697 (
            .O(N__25425),
            .I(N__25418));
    InMux I__3696 (
            .O(N__25424),
            .I(N__25415));
    InMux I__3695 (
            .O(N__25421),
            .I(N__25412));
    Odrv4 I__3694 (
            .O(N__25418),
            .I(cmd_rdadctmp_22_adj_1450));
    LocalMux I__3693 (
            .O(N__25415),
            .I(cmd_rdadctmp_22_adj_1450));
    LocalMux I__3692 (
            .O(N__25412),
            .I(cmd_rdadctmp_22_adj_1450));
    InMux I__3691 (
            .O(N__25405),
            .I(\ADC_VDC.n19385 ));
    CascadeMux I__3690 (
            .O(N__25402),
            .I(N__25398));
    CascadeMux I__3689 (
            .O(N__25401),
            .I(N__25395));
    InMux I__3688 (
            .O(N__25398),
            .I(N__25392));
    InMux I__3687 (
            .O(N__25395),
            .I(N__25389));
    LocalMux I__3686 (
            .O(N__25392),
            .I(N__25386));
    LocalMux I__3685 (
            .O(N__25389),
            .I(\ADC_VDC.cmd_rdadctmp_23 ));
    Odrv4 I__3684 (
            .O(N__25386),
            .I(\ADC_VDC.cmd_rdadctmp_23 ));
    InMux I__3683 (
            .O(N__25381),
            .I(\ADC_VDC.n19386 ));
    InMux I__3682 (
            .O(N__25378),
            .I(N__25374));
    InMux I__3681 (
            .O(N__25377),
            .I(N__25371));
    LocalMux I__3680 (
            .O(N__25374),
            .I(cmd_rdadcbuf_24));
    LocalMux I__3679 (
            .O(N__25371),
            .I(cmd_rdadcbuf_24));
    InMux I__3678 (
            .O(N__25366),
            .I(bfn_9_8_0_));
    InMux I__3677 (
            .O(N__25363),
            .I(N__25359));
    InMux I__3676 (
            .O(N__25362),
            .I(N__25356));
    LocalMux I__3675 (
            .O(N__25359),
            .I(cmd_rdadcbuf_25));
    LocalMux I__3674 (
            .O(N__25356),
            .I(cmd_rdadcbuf_25));
    InMux I__3673 (
            .O(N__25351),
            .I(\ADC_VDC.n19388 ));
    InMux I__3672 (
            .O(N__25348),
            .I(N__25344));
    InMux I__3671 (
            .O(N__25347),
            .I(N__25341));
    LocalMux I__3670 (
            .O(N__25344),
            .I(cmd_rdadcbuf_26));
    LocalMux I__3669 (
            .O(N__25341),
            .I(cmd_rdadcbuf_26));
    InMux I__3668 (
            .O(N__25336),
            .I(\ADC_VDC.n19389 ));
    InMux I__3667 (
            .O(N__25333),
            .I(N__25329));
    InMux I__3666 (
            .O(N__25332),
            .I(N__25326));
    LocalMux I__3665 (
            .O(N__25329),
            .I(cmd_rdadcbuf_27));
    LocalMux I__3664 (
            .O(N__25326),
            .I(cmd_rdadcbuf_27));
    InMux I__3663 (
            .O(N__25321),
            .I(\ADC_VDC.n19390 ));
    InMux I__3662 (
            .O(N__25318),
            .I(N__25314));
    InMux I__3661 (
            .O(N__25317),
            .I(N__25311));
    LocalMux I__3660 (
            .O(N__25314),
            .I(cmd_rdadcbuf_11));
    LocalMux I__3659 (
            .O(N__25311),
            .I(cmd_rdadcbuf_11));
    InMux I__3658 (
            .O(N__25306),
            .I(\ADC_VDC.n19374 ));
    InMux I__3657 (
            .O(N__25303),
            .I(N__25299));
    InMux I__3656 (
            .O(N__25302),
            .I(N__25296));
    LocalMux I__3655 (
            .O(N__25299),
            .I(cmd_rdadcbuf_12));
    LocalMux I__3654 (
            .O(N__25296),
            .I(cmd_rdadcbuf_12));
    InMux I__3653 (
            .O(N__25291),
            .I(\ADC_VDC.n19375 ));
    CascadeMux I__3652 (
            .O(N__25288),
            .I(N__25283));
    InMux I__3651 (
            .O(N__25287),
            .I(N__25278));
    InMux I__3650 (
            .O(N__25286),
            .I(N__25278));
    InMux I__3649 (
            .O(N__25283),
            .I(N__25275));
    LocalMux I__3648 (
            .O(N__25278),
            .I(cmd_rdadctmp_13_adj_1459));
    LocalMux I__3647 (
            .O(N__25275),
            .I(cmd_rdadctmp_13_adj_1459));
    InMux I__3646 (
            .O(N__25270),
            .I(N__25267));
    LocalMux I__3645 (
            .O(N__25267),
            .I(N__25263));
    InMux I__3644 (
            .O(N__25266),
            .I(N__25260));
    Odrv4 I__3643 (
            .O(N__25263),
            .I(cmd_rdadcbuf_13));
    LocalMux I__3642 (
            .O(N__25260),
            .I(cmd_rdadcbuf_13));
    InMux I__3641 (
            .O(N__25255),
            .I(\ADC_VDC.n19376 ));
    CascadeMux I__3640 (
            .O(N__25252),
            .I(N__25249));
    InMux I__3639 (
            .O(N__25249),
            .I(N__25244));
    CascadeMux I__3638 (
            .O(N__25248),
            .I(N__25241));
    CascadeMux I__3637 (
            .O(N__25247),
            .I(N__25238));
    LocalMux I__3636 (
            .O(N__25244),
            .I(N__25235));
    InMux I__3635 (
            .O(N__25241),
            .I(N__25232));
    InMux I__3634 (
            .O(N__25238),
            .I(N__25229));
    Odrv4 I__3633 (
            .O(N__25235),
            .I(cmd_rdadctmp_14_adj_1458));
    LocalMux I__3632 (
            .O(N__25232),
            .I(cmd_rdadctmp_14_adj_1458));
    LocalMux I__3631 (
            .O(N__25229),
            .I(cmd_rdadctmp_14_adj_1458));
    InMux I__3630 (
            .O(N__25222),
            .I(N__25218));
    InMux I__3629 (
            .O(N__25221),
            .I(N__25215));
    LocalMux I__3628 (
            .O(N__25218),
            .I(cmd_rdadcbuf_14));
    LocalMux I__3627 (
            .O(N__25215),
            .I(cmd_rdadcbuf_14));
    InMux I__3626 (
            .O(N__25210),
            .I(\ADC_VDC.n19377 ));
    InMux I__3625 (
            .O(N__25207),
            .I(\ADC_VDC.n19378 ));
    InMux I__3624 (
            .O(N__25204),
            .I(bfn_9_7_0_));
    InMux I__3623 (
            .O(N__25201),
            .I(\ADC_VDC.n19380 ));
    CascadeMux I__3622 (
            .O(N__25198),
            .I(N__25194));
    CascadeMux I__3621 (
            .O(N__25197),
            .I(N__25190));
    InMux I__3620 (
            .O(N__25194),
            .I(N__25187));
    InMux I__3619 (
            .O(N__25193),
            .I(N__25184));
    InMux I__3618 (
            .O(N__25190),
            .I(N__25181));
    LocalMux I__3617 (
            .O(N__25187),
            .I(cmd_rdadctmp_18_adj_1454));
    LocalMux I__3616 (
            .O(N__25184),
            .I(cmd_rdadctmp_18_adj_1454));
    LocalMux I__3615 (
            .O(N__25181),
            .I(cmd_rdadctmp_18_adj_1454));
    InMux I__3614 (
            .O(N__25174),
            .I(\ADC_VDC.n19381 ));
    InMux I__3613 (
            .O(N__25171),
            .I(\ADC_VDC.n19382 ));
    InMux I__3612 (
            .O(N__25168),
            .I(N__25165));
    LocalMux I__3611 (
            .O(N__25165),
            .I(\ADC_VDC.cmd_rdadcbuf_3 ));
    InMux I__3610 (
            .O(N__25162),
            .I(\ADC_VDC.n19366 ));
    InMux I__3609 (
            .O(N__25159),
            .I(N__25156));
    LocalMux I__3608 (
            .O(N__25156),
            .I(\ADC_VDC.cmd_rdadcbuf_4 ));
    InMux I__3607 (
            .O(N__25153),
            .I(\ADC_VDC.n19367 ));
    CascadeMux I__3606 (
            .O(N__25150),
            .I(N__25145));
    InMux I__3605 (
            .O(N__25149),
            .I(N__25140));
    InMux I__3604 (
            .O(N__25148),
            .I(N__25140));
    InMux I__3603 (
            .O(N__25145),
            .I(N__25137));
    LocalMux I__3602 (
            .O(N__25140),
            .I(cmd_rdadctmp_5_adj_1467));
    LocalMux I__3601 (
            .O(N__25137),
            .I(cmd_rdadctmp_5_adj_1467));
    InMux I__3600 (
            .O(N__25132),
            .I(N__25129));
    LocalMux I__3599 (
            .O(N__25129),
            .I(\ADC_VDC.cmd_rdadcbuf_5 ));
    InMux I__3598 (
            .O(N__25126),
            .I(\ADC_VDC.n19368 ));
    CascadeMux I__3597 (
            .O(N__25123),
            .I(N__25118));
    InMux I__3596 (
            .O(N__25122),
            .I(N__25113));
    InMux I__3595 (
            .O(N__25121),
            .I(N__25113));
    InMux I__3594 (
            .O(N__25118),
            .I(N__25110));
    LocalMux I__3593 (
            .O(N__25113),
            .I(cmd_rdadctmp_6_adj_1466));
    LocalMux I__3592 (
            .O(N__25110),
            .I(cmd_rdadctmp_6_adj_1466));
    InMux I__3591 (
            .O(N__25105),
            .I(N__25102));
    LocalMux I__3590 (
            .O(N__25102),
            .I(\ADC_VDC.cmd_rdadcbuf_6 ));
    InMux I__3589 (
            .O(N__25099),
            .I(\ADC_VDC.n19369 ));
    InMux I__3588 (
            .O(N__25096),
            .I(N__25093));
    LocalMux I__3587 (
            .O(N__25093),
            .I(\ADC_VDC.cmd_rdadcbuf_7 ));
    InMux I__3586 (
            .O(N__25090),
            .I(\ADC_VDC.n19370 ));
    InMux I__3585 (
            .O(N__25087),
            .I(N__25084));
    LocalMux I__3584 (
            .O(N__25084),
            .I(\ADC_VDC.cmd_rdadcbuf_8 ));
    InMux I__3583 (
            .O(N__25081),
            .I(bfn_9_6_0_));
    InMux I__3582 (
            .O(N__25078),
            .I(N__25071));
    InMux I__3581 (
            .O(N__25077),
            .I(N__25071));
    InMux I__3580 (
            .O(N__25076),
            .I(N__25068));
    LocalMux I__3579 (
            .O(N__25071),
            .I(cmd_rdadctmp_9_adj_1463));
    LocalMux I__3578 (
            .O(N__25068),
            .I(cmd_rdadctmp_9_adj_1463));
    CascadeMux I__3577 (
            .O(N__25063),
            .I(N__25060));
    InMux I__3576 (
            .O(N__25060),
            .I(N__25057));
    LocalMux I__3575 (
            .O(N__25057),
            .I(\ADC_VDC.cmd_rdadcbuf_9 ));
    InMux I__3574 (
            .O(N__25054),
            .I(\ADC_VDC.n19372 ));
    InMux I__3573 (
            .O(N__25051),
            .I(N__25048));
    LocalMux I__3572 (
            .O(N__25048),
            .I(\ADC_VDC.cmd_rdadcbuf_10 ));
    InMux I__3571 (
            .O(N__25045),
            .I(\ADC_VDC.n19373 ));
    InMux I__3570 (
            .O(N__25042),
            .I(N__25038));
    InMux I__3569 (
            .O(N__25041),
            .I(N__25035));
    LocalMux I__3568 (
            .O(N__25038),
            .I(N__25032));
    LocalMux I__3567 (
            .O(N__25035),
            .I(\ADC_IAC.bit_cnt_5 ));
    Odrv4 I__3566 (
            .O(N__25032),
            .I(\ADC_IAC.bit_cnt_5 ));
    CascadeMux I__3565 (
            .O(N__25027),
            .I(\ADC_IAC.n20765_cascade_ ));
    CascadeMux I__3564 (
            .O(N__25024),
            .I(\ADC_IAC.n21007_cascade_ ));
    CEMux I__3563 (
            .O(N__25021),
            .I(N__25018));
    LocalMux I__3562 (
            .O(N__25018),
            .I(N__25015));
    Odrv4 I__3561 (
            .O(N__25015),
            .I(\ADC_IAC.n20670 ));
    CascadeMux I__3560 (
            .O(N__25012),
            .I(N__25009));
    InMux I__3559 (
            .O(N__25009),
            .I(N__25004));
    InMux I__3558 (
            .O(N__25008),
            .I(N__25001));
    InMux I__3557 (
            .O(N__25007),
            .I(N__24998));
    LocalMux I__3556 (
            .O(N__25004),
            .I(N__24990));
    LocalMux I__3555 (
            .O(N__25001),
            .I(N__24990));
    LocalMux I__3554 (
            .O(N__24998),
            .I(N__24990));
    CascadeMux I__3553 (
            .O(N__24997),
            .I(N__24986));
    Span4Mux_h I__3552 (
            .O(N__24990),
            .I(N__24983));
    InMux I__3551 (
            .O(N__24989),
            .I(N__24978));
    InMux I__3550 (
            .O(N__24986),
            .I(N__24978));
    Span4Mux_v I__3549 (
            .O(N__24983),
            .I(N__24975));
    LocalMux I__3548 (
            .O(N__24978),
            .I(N__24972));
    Span4Mux_v I__3547 (
            .O(N__24975),
            .I(N__24969));
    Span12Mux_h I__3546 (
            .O(N__24972),
            .I(N__24966));
    Span4Mux_h I__3545 (
            .O(N__24969),
            .I(N__24963));
    Odrv12 I__3544 (
            .O(N__24966),
            .I(IAC_DRDY));
    Odrv4 I__3543 (
            .O(N__24963),
            .I(IAC_DRDY));
    CascadeMux I__3542 (
            .O(N__24958),
            .I(\ADC_IAC.n17_cascade_ ));
    CEMux I__3541 (
            .O(N__24955),
            .I(N__24952));
    LocalMux I__3540 (
            .O(N__24952),
            .I(N__24949));
    Odrv4 I__3539 (
            .O(N__24949),
            .I(\ADC_IAC.n12 ));
    SRMux I__3538 (
            .O(N__24946),
            .I(N__24943));
    LocalMux I__3537 (
            .O(N__24943),
            .I(N__24940));
    Span4Mux_h I__3536 (
            .O(N__24940),
            .I(N__24937));
    Span4Mux_h I__3535 (
            .O(N__24937),
            .I(N__24934));
    Odrv4 I__3534 (
            .O(N__24934),
            .I(\ADC_VDC.n20345 ));
    InMux I__3533 (
            .O(N__24931),
            .I(N__24928));
    LocalMux I__3532 (
            .O(N__24928),
            .I(\ADC_VDC.cmd_rdadcbuf_0 ));
    InMux I__3531 (
            .O(N__24925),
            .I(N__24922));
    LocalMux I__3530 (
            .O(N__24922),
            .I(\ADC_VDC.cmd_rdadcbuf_1 ));
    InMux I__3529 (
            .O(N__24919),
            .I(\ADC_VDC.n19364 ));
    CascadeMux I__3528 (
            .O(N__24916),
            .I(N__24913));
    InMux I__3527 (
            .O(N__24913),
            .I(N__24910));
    LocalMux I__3526 (
            .O(N__24910),
            .I(\ADC_VDC.cmd_rdadcbuf_2 ));
    InMux I__3525 (
            .O(N__24907),
            .I(\ADC_VDC.n19365 ));
    CascadeMux I__3524 (
            .O(N__24904),
            .I(N__24900));
    InMux I__3523 (
            .O(N__24903),
            .I(N__24896));
    InMux I__3522 (
            .O(N__24900),
            .I(N__24891));
    InMux I__3521 (
            .O(N__24899),
            .I(N__24891));
    LocalMux I__3520 (
            .O(N__24896),
            .I(cmd_rdadctmp_30));
    LocalMux I__3519 (
            .O(N__24891),
            .I(cmd_rdadctmp_30));
    InMux I__3518 (
            .O(N__24886),
            .I(N__24882));
    InMux I__3517 (
            .O(N__24885),
            .I(N__24879));
    LocalMux I__3516 (
            .O(N__24882),
            .I(cmd_rdadctmp_4));
    LocalMux I__3515 (
            .O(N__24879),
            .I(cmd_rdadctmp_4));
    CascadeMux I__3514 (
            .O(N__24874),
            .I(N__24871));
    InMux I__3513 (
            .O(N__24871),
            .I(N__24867));
    InMux I__3512 (
            .O(N__24870),
            .I(N__24864));
    LocalMux I__3511 (
            .O(N__24867),
            .I(cmd_rdadctmp_2));
    LocalMux I__3510 (
            .O(N__24864),
            .I(cmd_rdadctmp_2));
    CascadeMux I__3509 (
            .O(N__24859),
            .I(N__24856));
    InMux I__3508 (
            .O(N__24856),
            .I(N__24850));
    InMux I__3507 (
            .O(N__24855),
            .I(N__24850));
    LocalMux I__3506 (
            .O(N__24850),
            .I(cmd_rdadctmp_3));
    IoInMux I__3505 (
            .O(N__24847),
            .I(N__24844));
    LocalMux I__3504 (
            .O(N__24844),
            .I(N__24841));
    Span4Mux_s0_v I__3503 (
            .O(N__24841),
            .I(N__24838));
    Sp12to4 I__3502 (
            .O(N__24838),
            .I(N__24834));
    CascadeMux I__3501 (
            .O(N__24837),
            .I(N__24831));
    Span12Mux_s11_h I__3500 (
            .O(N__24834),
            .I(N__24828));
    InMux I__3499 (
            .O(N__24831),
            .I(N__24825));
    Odrv12 I__3498 (
            .O(N__24828),
            .I(IAC_CS));
    LocalMux I__3497 (
            .O(N__24825),
            .I(IAC_CS));
    InMux I__3496 (
            .O(N__24820),
            .I(N__24817));
    LocalMux I__3495 (
            .O(N__24817),
            .I(n14_adj_1581));
    InMux I__3494 (
            .O(N__24814),
            .I(N__24811));
    LocalMux I__3493 (
            .O(N__24811),
            .I(\ADC_IAC.n20669 ));
    InMux I__3492 (
            .O(N__24808),
            .I(N__24804));
    InMux I__3491 (
            .O(N__24807),
            .I(N__24801));
    LocalMux I__3490 (
            .O(N__24804),
            .I(\ADC_IAC.bit_cnt_4 ));
    LocalMux I__3489 (
            .O(N__24801),
            .I(\ADC_IAC.bit_cnt_4 ));
    InMux I__3488 (
            .O(N__24796),
            .I(N__24792));
    InMux I__3487 (
            .O(N__24795),
            .I(N__24789));
    LocalMux I__3486 (
            .O(N__24792),
            .I(\ADC_IAC.bit_cnt_3 ));
    LocalMux I__3485 (
            .O(N__24789),
            .I(\ADC_IAC.bit_cnt_3 ));
    CascadeMux I__3484 (
            .O(N__24784),
            .I(N__24780));
    InMux I__3483 (
            .O(N__24783),
            .I(N__24777));
    InMux I__3482 (
            .O(N__24780),
            .I(N__24774));
    LocalMux I__3481 (
            .O(N__24777),
            .I(\ADC_IAC.bit_cnt_1 ));
    LocalMux I__3480 (
            .O(N__24774),
            .I(\ADC_IAC.bit_cnt_1 ));
    InMux I__3479 (
            .O(N__24769),
            .I(N__24765));
    InMux I__3478 (
            .O(N__24768),
            .I(N__24762));
    LocalMux I__3477 (
            .O(N__24765),
            .I(\ADC_IAC.bit_cnt_2 ));
    LocalMux I__3476 (
            .O(N__24762),
            .I(\ADC_IAC.bit_cnt_2 ));
    InMux I__3475 (
            .O(N__24757),
            .I(N__24753));
    InMux I__3474 (
            .O(N__24756),
            .I(N__24750));
    LocalMux I__3473 (
            .O(N__24753),
            .I(\ADC_IAC.bit_cnt_6 ));
    LocalMux I__3472 (
            .O(N__24750),
            .I(\ADC_IAC.bit_cnt_6 ));
    InMux I__3471 (
            .O(N__24745),
            .I(N__24741));
    InMux I__3470 (
            .O(N__24744),
            .I(N__24738));
    LocalMux I__3469 (
            .O(N__24741),
            .I(\ADC_IAC.bit_cnt_0 ));
    LocalMux I__3468 (
            .O(N__24738),
            .I(\ADC_IAC.bit_cnt_0 ));
    CascadeMux I__3467 (
            .O(N__24733),
            .I(\ADC_IAC.n20753_cascade_ ));
    InMux I__3466 (
            .O(N__24730),
            .I(N__24726));
    InMux I__3465 (
            .O(N__24729),
            .I(N__24723));
    LocalMux I__3464 (
            .O(N__24726),
            .I(\ADC_IAC.bit_cnt_7 ));
    LocalMux I__3463 (
            .O(N__24723),
            .I(\ADC_IAC.bit_cnt_7 ));
    CascadeMux I__3462 (
            .O(N__24718),
            .I(N__24715));
    InMux I__3461 (
            .O(N__24715),
            .I(N__24712));
    LocalMux I__3460 (
            .O(N__24712),
            .I(N__24708));
    InMux I__3459 (
            .O(N__24711),
            .I(N__24705));
    Odrv4 I__3458 (
            .O(N__24708),
            .I(cmd_rdadctmp_5));
    LocalMux I__3457 (
            .O(N__24705),
            .I(cmd_rdadctmp_5));
    InMux I__3456 (
            .O(N__24700),
            .I(N__24697));
    LocalMux I__3455 (
            .O(N__24697),
            .I(N__24694));
    Span4Mux_v I__3454 (
            .O(N__24694),
            .I(N__24691));
    Span4Mux_v I__3453 (
            .O(N__24691),
            .I(N__24687));
    InMux I__3452 (
            .O(N__24690),
            .I(N__24684));
    Span4Mux_v I__3451 (
            .O(N__24687),
            .I(N__24678));
    LocalMux I__3450 (
            .O(N__24684),
            .I(N__24678));
    InMux I__3449 (
            .O(N__24683),
            .I(N__24675));
    Span4Mux_h I__3448 (
            .O(N__24678),
            .I(N__24672));
    LocalMux I__3447 (
            .O(N__24675),
            .I(buf_adcdata_iac_22));
    Odrv4 I__3446 (
            .O(N__24672),
            .I(buf_adcdata_iac_22));
    InMux I__3445 (
            .O(N__24667),
            .I(N__24661));
    InMux I__3444 (
            .O(N__24666),
            .I(N__24661));
    LocalMux I__3443 (
            .O(N__24661),
            .I(cmd_rdadctmp_1));
    InMux I__3442 (
            .O(N__24658),
            .I(N__24654));
    InMux I__3441 (
            .O(N__24657),
            .I(N__24651));
    LocalMux I__3440 (
            .O(N__24654),
            .I(n20553));
    LocalMux I__3439 (
            .O(N__24651),
            .I(n20553));
    CascadeMux I__3438 (
            .O(N__24646),
            .I(N__24641));
    CascadeMux I__3437 (
            .O(N__24645),
            .I(N__24638));
    CascadeMux I__3436 (
            .O(N__24644),
            .I(N__24635));
    InMux I__3435 (
            .O(N__24641),
            .I(N__24632));
    InMux I__3434 (
            .O(N__24638),
            .I(N__24629));
    InMux I__3433 (
            .O(N__24635),
            .I(N__24626));
    LocalMux I__3432 (
            .O(N__24632),
            .I(N__24623));
    LocalMux I__3431 (
            .O(N__24629),
            .I(cmd_rdadctmp_29));
    LocalMux I__3430 (
            .O(N__24626),
            .I(cmd_rdadctmp_29));
    Odrv4 I__3429 (
            .O(N__24623),
            .I(cmd_rdadctmp_29));
    CascadeMux I__3428 (
            .O(N__24616),
            .I(N__24613));
    InMux I__3427 (
            .O(N__24613),
            .I(N__24608));
    InMux I__3426 (
            .O(N__24612),
            .I(N__24605));
    InMux I__3425 (
            .O(N__24611),
            .I(N__24602));
    LocalMux I__3424 (
            .O(N__24608),
            .I(cmd_rdadctmp_27));
    LocalMux I__3423 (
            .O(N__24605),
            .I(cmd_rdadctmp_27));
    LocalMux I__3422 (
            .O(N__24602),
            .I(cmd_rdadctmp_27));
    CascadeMux I__3421 (
            .O(N__24595),
            .I(N__24592));
    InMux I__3420 (
            .O(N__24592),
            .I(N__24589));
    LocalMux I__3419 (
            .O(N__24589),
            .I(N__24586));
    Span4Mux_v I__3418 (
            .O(N__24586),
            .I(N__24583));
    Sp12to4 I__3417 (
            .O(N__24583),
            .I(N__24580));
    Span12Mux_h I__3416 (
            .O(N__24580),
            .I(N__24577));
    Odrv12 I__3415 (
            .O(N__24577),
            .I(IAC_MISO));
    InMux I__3414 (
            .O(N__24574),
            .I(N__24570));
    InMux I__3413 (
            .O(N__24573),
            .I(N__24567));
    LocalMux I__3412 (
            .O(N__24570),
            .I(cmd_rdadctmp_0));
    LocalMux I__3411 (
            .O(N__24567),
            .I(cmd_rdadctmp_0));
    CascadeMux I__3410 (
            .O(N__24562),
            .I(N__24559));
    InMux I__3409 (
            .O(N__24559),
            .I(N__24553));
    InMux I__3408 (
            .O(N__24558),
            .I(N__24553));
    LocalMux I__3407 (
            .O(N__24553),
            .I(cmd_rdadctmp_6));
    CascadeMux I__3406 (
            .O(N__24550),
            .I(N__24547));
    CascadeBuf I__3405 (
            .O(N__24547),
            .I(N__24544));
    CascadeMux I__3404 (
            .O(N__24544),
            .I(N__24541));
    CascadeBuf I__3403 (
            .O(N__24541),
            .I(N__24538));
    CascadeMux I__3402 (
            .O(N__24538),
            .I(N__24535));
    CascadeBuf I__3401 (
            .O(N__24535),
            .I(N__24532));
    CascadeMux I__3400 (
            .O(N__24532),
            .I(N__24529));
    CascadeBuf I__3399 (
            .O(N__24529),
            .I(N__24526));
    CascadeMux I__3398 (
            .O(N__24526),
            .I(N__24523));
    CascadeBuf I__3397 (
            .O(N__24523),
            .I(N__24520));
    CascadeMux I__3396 (
            .O(N__24520),
            .I(N__24517));
    CascadeBuf I__3395 (
            .O(N__24517),
            .I(N__24514));
    CascadeMux I__3394 (
            .O(N__24514),
            .I(N__24510));
    CascadeMux I__3393 (
            .O(N__24513),
            .I(N__24507));
    CascadeBuf I__3392 (
            .O(N__24510),
            .I(N__24504));
    CascadeBuf I__3391 (
            .O(N__24507),
            .I(N__24501));
    CascadeMux I__3390 (
            .O(N__24504),
            .I(N__24498));
    CascadeMux I__3389 (
            .O(N__24501),
            .I(N__24495));
    CascadeBuf I__3388 (
            .O(N__24498),
            .I(N__24492));
    InMux I__3387 (
            .O(N__24495),
            .I(N__24489));
    CascadeMux I__3386 (
            .O(N__24492),
            .I(N__24486));
    LocalMux I__3385 (
            .O(N__24489),
            .I(N__24483));
    CascadeBuf I__3384 (
            .O(N__24486),
            .I(N__24480));
    Span4Mux_v I__3383 (
            .O(N__24483),
            .I(N__24477));
    CascadeMux I__3382 (
            .O(N__24480),
            .I(N__24474));
    Span4Mux_h I__3381 (
            .O(N__24477),
            .I(N__24471));
    InMux I__3380 (
            .O(N__24474),
            .I(N__24468));
    Span4Mux_h I__3379 (
            .O(N__24471),
            .I(N__24465));
    LocalMux I__3378 (
            .O(N__24468),
            .I(N__24462));
    Span4Mux_h I__3377 (
            .O(N__24465),
            .I(N__24457));
    Span4Mux_v I__3376 (
            .O(N__24462),
            .I(N__24457));
    Odrv4 I__3375 (
            .O(N__24457),
            .I(data_index_9_N_212_8));
    InMux I__3374 (
            .O(N__24454),
            .I(N__24450));
    CascadeMux I__3373 (
            .O(N__24453),
            .I(N__24447));
    LocalMux I__3372 (
            .O(N__24450),
            .I(N__24443));
    InMux I__3371 (
            .O(N__24447),
            .I(N__24438));
    InMux I__3370 (
            .O(N__24446),
            .I(N__24438));
    Odrv4 I__3369 (
            .O(N__24443),
            .I(cmd_rdadctmp_22));
    LocalMux I__3368 (
            .O(N__24438),
            .I(cmd_rdadctmp_22));
    InMux I__3367 (
            .O(N__24433),
            .I(N__24427));
    InMux I__3366 (
            .O(N__24432),
            .I(N__24427));
    LocalMux I__3365 (
            .O(N__24427),
            .I(n8_adj_1534));
    InMux I__3364 (
            .O(N__24424),
            .I(N__24421));
    LocalMux I__3363 (
            .O(N__24421),
            .I(N__24417));
    CascadeMux I__3362 (
            .O(N__24420),
            .I(N__24414));
    Span4Mux_v I__3361 (
            .O(N__24417),
            .I(N__24410));
    InMux I__3360 (
            .O(N__24414),
            .I(N__24407));
    InMux I__3359 (
            .O(N__24413),
            .I(N__24404));
    Span4Mux_h I__3358 (
            .O(N__24410),
            .I(N__24399));
    LocalMux I__3357 (
            .O(N__24407),
            .I(N__24399));
    LocalMux I__3356 (
            .O(N__24404),
            .I(buf_adcdata_iac_8));
    Odrv4 I__3355 (
            .O(N__24399),
            .I(buf_adcdata_iac_8));
    InMux I__3354 (
            .O(N__24394),
            .I(N__24391));
    LocalMux I__3353 (
            .O(N__24391),
            .I(N__24388));
    Span4Mux_v I__3352 (
            .O(N__24388),
            .I(N__24385));
    Span4Mux_h I__3351 (
            .O(N__24385),
            .I(N__24382));
    Sp12to4 I__3350 (
            .O(N__24382),
            .I(N__24379));
    Odrv12 I__3349 (
            .O(N__24379),
            .I(buf_data_iac_23));
    CascadeMux I__3348 (
            .O(N__24376),
            .I(n26_adj_1511_cascade_));
    CascadeMux I__3347 (
            .O(N__24373),
            .I(n20834_cascade_));
    CascadeMux I__3346 (
            .O(N__24370),
            .I(n22057_cascade_));
    InMux I__3345 (
            .O(N__24367),
            .I(N__24364));
    LocalMux I__3344 (
            .O(N__24364),
            .I(N__24361));
    Span4Mux_v I__3343 (
            .O(N__24361),
            .I(N__24358));
    Odrv4 I__3342 (
            .O(N__24358),
            .I(buf_data_iac_12));
    InMux I__3341 (
            .O(N__24355),
            .I(N__24352));
    LocalMux I__3340 (
            .O(N__24352),
            .I(N__24349));
    Odrv4 I__3339 (
            .O(N__24349),
            .I(n22135));
    InMux I__3338 (
            .O(N__24346),
            .I(N__24343));
    LocalMux I__3337 (
            .O(N__24343),
            .I(N__24339));
    InMux I__3336 (
            .O(N__24342),
            .I(N__24335));
    Span4Mux_v I__3335 (
            .O(N__24339),
            .I(N__24332));
    CascadeMux I__3334 (
            .O(N__24338),
            .I(N__24329));
    LocalMux I__3333 (
            .O(N__24335),
            .I(N__24326));
    Span4Mux_v I__3332 (
            .O(N__24332),
            .I(N__24323));
    InMux I__3331 (
            .O(N__24329),
            .I(N__24320));
    Span4Mux_v I__3330 (
            .O(N__24326),
            .I(N__24315));
    Span4Mux_v I__3329 (
            .O(N__24323),
            .I(N__24315));
    LocalMux I__3328 (
            .O(N__24320),
            .I(buf_adcdata_vac_23));
    Odrv4 I__3327 (
            .O(N__24315),
            .I(buf_adcdata_vac_23));
    InMux I__3326 (
            .O(N__24310),
            .I(N__24306));
    CascadeMux I__3325 (
            .O(N__24309),
            .I(N__24303));
    LocalMux I__3324 (
            .O(N__24306),
            .I(N__24300));
    InMux I__3323 (
            .O(N__24303),
            .I(N__24297));
    Odrv12 I__3322 (
            .O(N__24300),
            .I(buf_adcdata_vdc_23));
    LocalMux I__3321 (
            .O(N__24297),
            .I(buf_adcdata_vdc_23));
    InMux I__3320 (
            .O(N__24292),
            .I(N__24289));
    LocalMux I__3319 (
            .O(N__24289),
            .I(n20831));
    InMux I__3318 (
            .O(N__24286),
            .I(N__24283));
    LocalMux I__3317 (
            .O(N__24283),
            .I(N__24280));
    Span4Mux_h I__3316 (
            .O(N__24280),
            .I(N__24276));
    InMux I__3315 (
            .O(N__24279),
            .I(N__24273));
    Odrv4 I__3314 (
            .O(N__24276),
            .I(cmd_rdadctmp_7));
    LocalMux I__3313 (
            .O(N__24273),
            .I(cmd_rdadctmp_7));
    InMux I__3312 (
            .O(N__24268),
            .I(N__24265));
    LocalMux I__3311 (
            .O(N__24265),
            .I(N__24262));
    Span4Mux_v I__3310 (
            .O(N__24262),
            .I(N__24259));
    Odrv4 I__3309 (
            .O(N__24259),
            .I(n16_adj_1507));
    InMux I__3308 (
            .O(N__24256),
            .I(N__24252));
    InMux I__3307 (
            .O(N__24255),
            .I(N__24248));
    LocalMux I__3306 (
            .O(N__24252),
            .I(N__24245));
    InMux I__3305 (
            .O(N__24251),
            .I(N__24242));
    LocalMux I__3304 (
            .O(N__24248),
            .I(cmd_rdadctmp_24_adj_1419));
    Odrv4 I__3303 (
            .O(N__24245),
            .I(cmd_rdadctmp_24_adj_1419));
    LocalMux I__3302 (
            .O(N__24242),
            .I(cmd_rdadctmp_24_adj_1419));
    InMux I__3301 (
            .O(N__24235),
            .I(N__24231));
    InMux I__3300 (
            .O(N__24234),
            .I(N__24227));
    LocalMux I__3299 (
            .O(N__24231),
            .I(N__24224));
    InMux I__3298 (
            .O(N__24230),
            .I(N__24221));
    LocalMux I__3297 (
            .O(N__24227),
            .I(cmd_rdadctmp_25_adj_1418));
    Odrv4 I__3296 (
            .O(N__24224),
            .I(cmd_rdadctmp_25_adj_1418));
    LocalMux I__3295 (
            .O(N__24221),
            .I(cmd_rdadctmp_25_adj_1418));
    InMux I__3294 (
            .O(N__24214),
            .I(N__24211));
    LocalMux I__3293 (
            .O(N__24211),
            .I(N__24208));
    Odrv4 I__3292 (
            .O(N__24208),
            .I(n22039));
    InMux I__3291 (
            .O(N__24205),
            .I(N__24202));
    LocalMux I__3290 (
            .O(N__24202),
            .I(n22042));
    CascadeMux I__3289 (
            .O(N__24199),
            .I(N__24196));
    InMux I__3288 (
            .O(N__24196),
            .I(N__24191));
    CascadeMux I__3287 (
            .O(N__24195),
            .I(N__24188));
    CascadeMux I__3286 (
            .O(N__24194),
            .I(N__24185));
    LocalMux I__3285 (
            .O(N__24191),
            .I(N__24182));
    InMux I__3284 (
            .O(N__24188),
            .I(N__24179));
    InMux I__3283 (
            .O(N__24185),
            .I(N__24176));
    Span4Mux_v I__3282 (
            .O(N__24182),
            .I(N__24172));
    LocalMux I__3281 (
            .O(N__24179),
            .I(N__24167));
    LocalMux I__3280 (
            .O(N__24176),
            .I(N__24167));
    InMux I__3279 (
            .O(N__24175),
            .I(N__24163));
    Span4Mux_v I__3278 (
            .O(N__24172),
            .I(N__24160));
    Span4Mux_h I__3277 (
            .O(N__24167),
            .I(N__24157));
    InMux I__3276 (
            .O(N__24166),
            .I(N__24154));
    LocalMux I__3275 (
            .O(N__24163),
            .I(N__24151));
    Odrv4 I__3274 (
            .O(N__24160),
            .I(buf_cfgRTD_7));
    Odrv4 I__3273 (
            .O(N__24157),
            .I(buf_cfgRTD_7));
    LocalMux I__3272 (
            .O(N__24154),
            .I(buf_cfgRTD_7));
    Odrv4 I__3271 (
            .O(N__24151),
            .I(buf_cfgRTD_7));
    CascadeMux I__3270 (
            .O(N__24142),
            .I(N__24139));
    InMux I__3269 (
            .O(N__24139),
            .I(N__24135));
    CascadeMux I__3268 (
            .O(N__24138),
            .I(N__24132));
    LocalMux I__3267 (
            .O(N__24135),
            .I(N__24129));
    InMux I__3266 (
            .O(N__24132),
            .I(N__24125));
    Span4Mux_h I__3265 (
            .O(N__24129),
            .I(N__24122));
    InMux I__3264 (
            .O(N__24128),
            .I(N__24119));
    LocalMux I__3263 (
            .O(N__24125),
            .I(cmd_rdadctmp_20_adj_1423));
    Odrv4 I__3262 (
            .O(N__24122),
            .I(cmd_rdadctmp_20_adj_1423));
    LocalMux I__3261 (
            .O(N__24119),
            .I(cmd_rdadctmp_20_adj_1423));
    InMux I__3260 (
            .O(N__24112),
            .I(N__24107));
    InMux I__3259 (
            .O(N__24111),
            .I(N__24102));
    InMux I__3258 (
            .O(N__24110),
            .I(N__24102));
    LocalMux I__3257 (
            .O(N__24107),
            .I(cmd_rdadctmp_18_adj_1425));
    LocalMux I__3256 (
            .O(N__24102),
            .I(cmd_rdadctmp_18_adj_1425));
    InMux I__3255 (
            .O(N__24097),
            .I(N__24094));
    LocalMux I__3254 (
            .O(N__24094),
            .I(N__24091));
    Span4Mux_h I__3253 (
            .O(N__24091),
            .I(N__24086));
    InMux I__3252 (
            .O(N__24090),
            .I(N__24081));
    InMux I__3251 (
            .O(N__24089),
            .I(N__24081));
    Odrv4 I__3250 (
            .O(N__24086),
            .I(buf_adcdata_vac_12));
    LocalMux I__3249 (
            .O(N__24081),
            .I(buf_adcdata_vac_12));
    InMux I__3248 (
            .O(N__24076),
            .I(N__24073));
    LocalMux I__3247 (
            .O(N__24073),
            .I(N__24069));
    CascadeMux I__3246 (
            .O(N__24072),
            .I(N__24066));
    Span4Mux_v I__3245 (
            .O(N__24069),
            .I(N__24063));
    InMux I__3244 (
            .O(N__24066),
            .I(N__24060));
    Odrv4 I__3243 (
            .O(N__24063),
            .I(buf_adcdata_vdc_10));
    LocalMux I__3242 (
            .O(N__24060),
            .I(buf_adcdata_vdc_10));
    InMux I__3241 (
            .O(N__24055),
            .I(N__24052));
    LocalMux I__3240 (
            .O(N__24052),
            .I(N__24049));
    Span4Mux_v I__3239 (
            .O(N__24049),
            .I(N__24046));
    Span4Mux_h I__3238 (
            .O(N__24046),
            .I(N__24041));
    InMux I__3237 (
            .O(N__24045),
            .I(N__24036));
    InMux I__3236 (
            .O(N__24044),
            .I(N__24036));
    Odrv4 I__3235 (
            .O(N__24041),
            .I(buf_adcdata_vac_10));
    LocalMux I__3234 (
            .O(N__24036),
            .I(buf_adcdata_vac_10));
    CascadeMux I__3233 (
            .O(N__24031),
            .I(N__24027));
    CascadeMux I__3232 (
            .O(N__24030),
            .I(N__24024));
    InMux I__3231 (
            .O(N__24027),
            .I(N__24021));
    InMux I__3230 (
            .O(N__24024),
            .I(N__24017));
    LocalMux I__3229 (
            .O(N__24021),
            .I(N__24014));
    InMux I__3228 (
            .O(N__24020),
            .I(N__24011));
    LocalMux I__3227 (
            .O(N__24017),
            .I(cmd_rdadctmp_19_adj_1424));
    Odrv4 I__3226 (
            .O(N__24014),
            .I(cmd_rdadctmp_19_adj_1424));
    LocalMux I__3225 (
            .O(N__24011),
            .I(cmd_rdadctmp_19_adj_1424));
    CascadeMux I__3224 (
            .O(N__24004),
            .I(N__24001));
    InMux I__3223 (
            .O(N__24001),
            .I(N__23998));
    LocalMux I__3222 (
            .O(N__23998),
            .I(N__23995));
    Span4Mux_h I__3221 (
            .O(N__23995),
            .I(N__23992));
    Odrv4 I__3220 (
            .O(N__23992),
            .I(buf_data_iac_16));
    CascadeMux I__3219 (
            .O(N__23989),
            .I(n20781_cascade_));
    InMux I__3218 (
            .O(N__23986),
            .I(N__23982));
    CascadeMux I__3217 (
            .O(N__23985),
            .I(N__23979));
    LocalMux I__3216 (
            .O(N__23982),
            .I(N__23976));
    InMux I__3215 (
            .O(N__23979),
            .I(N__23973));
    Odrv12 I__3214 (
            .O(N__23976),
            .I(buf_adcdata_vdc_1));
    LocalMux I__3213 (
            .O(N__23973),
            .I(buf_adcdata_vdc_1));
    InMux I__3212 (
            .O(N__23968),
            .I(N__23965));
    LocalMux I__3211 (
            .O(N__23965),
            .I(N__23962));
    Span4Mux_v I__3210 (
            .O(N__23962),
            .I(N__23957));
    InMux I__3209 (
            .O(N__23961),
            .I(N__23954));
    InMux I__3208 (
            .O(N__23960),
            .I(N__23951));
    Span4Mux_h I__3207 (
            .O(N__23957),
            .I(N__23946));
    LocalMux I__3206 (
            .O(N__23954),
            .I(N__23946));
    LocalMux I__3205 (
            .O(N__23951),
            .I(buf_adcdata_vac_1));
    Odrv4 I__3204 (
            .O(N__23946),
            .I(buf_adcdata_vac_1));
    InMux I__3203 (
            .O(N__23941),
            .I(N__23938));
    LocalMux I__3202 (
            .O(N__23938),
            .I(n19_adj_1617));
    CascadeMux I__3201 (
            .O(N__23935),
            .I(n22171_cascade_));
    InMux I__3200 (
            .O(N__23932),
            .I(N__23929));
    LocalMux I__3199 (
            .O(N__23929),
            .I(N__23926));
    Odrv4 I__3198 (
            .O(N__23926),
            .I(n20775));
    InMux I__3197 (
            .O(N__23923),
            .I(N__23920));
    LocalMux I__3196 (
            .O(N__23920),
            .I(N__23917));
    Span4Mux_h I__3195 (
            .O(N__23917),
            .I(N__23914));
    Odrv4 I__3194 (
            .O(N__23914),
            .I(n20842));
    CascadeMux I__3193 (
            .O(N__23911),
            .I(N__23908));
    InMux I__3192 (
            .O(N__23908),
            .I(N__23905));
    LocalMux I__3191 (
            .O(N__23905),
            .I(N__23902));
    Odrv4 I__3190 (
            .O(N__23902),
            .I(n20843));
    CascadeMux I__3189 (
            .O(N__23899),
            .I(n22051_cascade_));
    InMux I__3188 (
            .O(N__23896),
            .I(N__23893));
    LocalMux I__3187 (
            .O(N__23893),
            .I(N__23890));
    Odrv4 I__3186 (
            .O(N__23890),
            .I(n20828));
    InMux I__3185 (
            .O(N__23887),
            .I(N__23884));
    LocalMux I__3184 (
            .O(N__23884),
            .I(N__23881));
    Odrv4 I__3183 (
            .O(N__23881),
            .I(n20814));
    InMux I__3182 (
            .O(N__23878),
            .I(N__23875));
    LocalMux I__3181 (
            .O(N__23875),
            .I(N__23871));
    CascadeMux I__3180 (
            .O(N__23874),
            .I(N__23868));
    Span4Mux_v I__3179 (
            .O(N__23871),
            .I(N__23865));
    InMux I__3178 (
            .O(N__23868),
            .I(N__23862));
    Odrv4 I__3177 (
            .O(N__23865),
            .I(buf_adcdata_vdc_18));
    LocalMux I__3176 (
            .O(N__23862),
            .I(buf_adcdata_vdc_18));
    InMux I__3175 (
            .O(N__23857),
            .I(N__23853));
    InMux I__3174 (
            .O(N__23856),
            .I(N__23849));
    LocalMux I__3173 (
            .O(N__23853),
            .I(N__23846));
    InMux I__3172 (
            .O(N__23852),
            .I(N__23843));
    LocalMux I__3171 (
            .O(N__23849),
            .I(N__23840));
    Span4Mux_v I__3170 (
            .O(N__23846),
            .I(N__23837));
    LocalMux I__3169 (
            .O(N__23843),
            .I(buf_adcdata_vac_18));
    Odrv4 I__3168 (
            .O(N__23840),
            .I(buf_adcdata_vac_18));
    Odrv4 I__3167 (
            .O(N__23837),
            .I(buf_adcdata_vac_18));
    CascadeMux I__3166 (
            .O(N__23830),
            .I(n21931_cascade_));
    InMux I__3165 (
            .O(N__23827),
            .I(N__23824));
    LocalMux I__3164 (
            .O(N__23824),
            .I(N__23820));
    CascadeMux I__3163 (
            .O(N__23823),
            .I(N__23816));
    Span4Mux_v I__3162 (
            .O(N__23820),
            .I(N__23813));
    InMux I__3161 (
            .O(N__23819),
            .I(N__23810));
    InMux I__3160 (
            .O(N__23816),
            .I(N__23807));
    Sp12to4 I__3159 (
            .O(N__23813),
            .I(N__23800));
    LocalMux I__3158 (
            .O(N__23810),
            .I(N__23800));
    LocalMux I__3157 (
            .O(N__23807),
            .I(N__23797));
    InMux I__3156 (
            .O(N__23806),
            .I(N__23792));
    InMux I__3155 (
            .O(N__23805),
            .I(N__23792));
    Odrv12 I__3154 (
            .O(N__23800),
            .I(buf_cfgRTD_2));
    Odrv4 I__3153 (
            .O(N__23797),
            .I(buf_cfgRTD_2));
    LocalMux I__3152 (
            .O(N__23792),
            .I(buf_cfgRTD_2));
    CascadeMux I__3151 (
            .O(N__23785),
            .I(N__23782));
    InMux I__3150 (
            .O(N__23782),
            .I(N__23779));
    LocalMux I__3149 (
            .O(N__23779),
            .I(N__23774));
    CascadeMux I__3148 (
            .O(N__23778),
            .I(N__23771));
    CascadeMux I__3147 (
            .O(N__23777),
            .I(N__23768));
    Span4Mux_h I__3146 (
            .O(N__23774),
            .I(N__23764));
    InMux I__3145 (
            .O(N__23771),
            .I(N__23760));
    InMux I__3144 (
            .O(N__23768),
            .I(N__23755));
    InMux I__3143 (
            .O(N__23767),
            .I(N__23755));
    Sp12to4 I__3142 (
            .O(N__23764),
            .I(N__23752));
    InMux I__3141 (
            .O(N__23763),
            .I(N__23749));
    LocalMux I__3140 (
            .O(N__23760),
            .I(N__23744));
    LocalMux I__3139 (
            .O(N__23755),
            .I(N__23744));
    Odrv12 I__3138 (
            .O(N__23752),
            .I(buf_cfgRTD_3));
    LocalMux I__3137 (
            .O(N__23749),
            .I(buf_cfgRTD_3));
    Odrv4 I__3136 (
            .O(N__23744),
            .I(buf_cfgRTD_3));
    CascadeMux I__3135 (
            .O(N__23737),
            .I(N__23734));
    InMux I__3134 (
            .O(N__23734),
            .I(N__23729));
    InMux I__3133 (
            .O(N__23733),
            .I(N__23724));
    InMux I__3132 (
            .O(N__23732),
            .I(N__23724));
    LocalMux I__3131 (
            .O(N__23729),
            .I(N__23719));
    LocalMux I__3130 (
            .O(N__23724),
            .I(N__23719));
    Span4Mux_v I__3129 (
            .O(N__23719),
            .I(N__23714));
    InMux I__3128 (
            .O(N__23718),
            .I(N__23711));
    InMux I__3127 (
            .O(N__23717),
            .I(N__23708));
    Odrv4 I__3126 (
            .O(N__23714),
            .I(buf_cfgRTD_0));
    LocalMux I__3125 (
            .O(N__23711),
            .I(buf_cfgRTD_0));
    LocalMux I__3124 (
            .O(N__23708),
            .I(buf_cfgRTD_0));
    CascadeMux I__3123 (
            .O(N__23701),
            .I(n14490_cascade_));
    CascadeMux I__3122 (
            .O(N__23698),
            .I(N__23694));
    InMux I__3121 (
            .O(N__23697),
            .I(N__23691));
    InMux I__3120 (
            .O(N__23694),
            .I(N__23688));
    LocalMux I__3119 (
            .O(N__23691),
            .I(N__23683));
    LocalMux I__3118 (
            .O(N__23688),
            .I(N__23683));
    Span4Mux_v I__3117 (
            .O(N__23683),
            .I(N__23677));
    InMux I__3116 (
            .O(N__23682),
            .I(N__23674));
    InMux I__3115 (
            .O(N__23681),
            .I(N__23671));
    InMux I__3114 (
            .O(N__23680),
            .I(N__23668));
    Odrv4 I__3113 (
            .O(N__23677),
            .I(buf_cfgRTD_1));
    LocalMux I__3112 (
            .O(N__23674),
            .I(buf_cfgRTD_1));
    LocalMux I__3111 (
            .O(N__23671),
            .I(buf_cfgRTD_1));
    LocalMux I__3110 (
            .O(N__23668),
            .I(buf_cfgRTD_1));
    CascadeMux I__3109 (
            .O(N__23659),
            .I(N__23656));
    InMux I__3108 (
            .O(N__23656),
            .I(N__23653));
    LocalMux I__3107 (
            .O(N__23653),
            .I(N__23650));
    Span4Mux_v I__3106 (
            .O(N__23650),
            .I(N__23647));
    Span4Mux_h I__3105 (
            .O(N__23647),
            .I(N__23643));
    InMux I__3104 (
            .O(N__23646),
            .I(N__23640));
    Odrv4 I__3103 (
            .O(N__23643),
            .I(buf_readRTD_9));
    LocalMux I__3102 (
            .O(N__23640),
            .I(buf_readRTD_9));
    InMux I__3101 (
            .O(N__23635),
            .I(N__23632));
    LocalMux I__3100 (
            .O(N__23632),
            .I(n22165));
    InMux I__3099 (
            .O(N__23629),
            .I(N__23624));
    InMux I__3098 (
            .O(N__23628),
            .I(N__23621));
    CascadeMux I__3097 (
            .O(N__23627),
            .I(N__23618));
    LocalMux I__3096 (
            .O(N__23624),
            .I(N__23615));
    LocalMux I__3095 (
            .O(N__23621),
            .I(N__23612));
    InMux I__3094 (
            .O(N__23618),
            .I(N__23609));
    Span4Mux_v I__3093 (
            .O(N__23615),
            .I(N__23606));
    Span12Mux_s9_h I__3092 (
            .O(N__23612),
            .I(N__23603));
    LocalMux I__3091 (
            .O(N__23609),
            .I(buf_adcdata_iac_1));
    Odrv4 I__3090 (
            .O(N__23606),
            .I(buf_adcdata_iac_1));
    Odrv12 I__3089 (
            .O(N__23603),
            .I(buf_adcdata_iac_1));
    InMux I__3088 (
            .O(N__23596),
            .I(N__23593));
    LocalMux I__3087 (
            .O(N__23593),
            .I(N__23590));
    Span4Mux_v I__3086 (
            .O(N__23590),
            .I(N__23587));
    Odrv4 I__3085 (
            .O(N__23587),
            .I(buf_data_iac_1));
    CascadeMux I__3084 (
            .O(N__23584),
            .I(n22_adj_1618_cascade_));
    InMux I__3083 (
            .O(N__23581),
            .I(N__23578));
    LocalMux I__3082 (
            .O(N__23578),
            .I(N__23574));
    CascadeMux I__3081 (
            .O(N__23577),
            .I(N__23571));
    Span4Mux_v I__3080 (
            .O(N__23574),
            .I(N__23568));
    InMux I__3079 (
            .O(N__23571),
            .I(N__23565));
    Odrv4 I__3078 (
            .O(N__23568),
            .I(buf_adcdata_vdc_15));
    LocalMux I__3077 (
            .O(N__23565),
            .I(buf_adcdata_vdc_15));
    InMux I__3076 (
            .O(N__23560),
            .I(N__23557));
    LocalMux I__3075 (
            .O(N__23557),
            .I(N__23554));
    Span4Mux_v I__3074 (
            .O(N__23554),
            .I(N__23550));
    InMux I__3073 (
            .O(N__23553),
            .I(N__23547));
    Odrv4 I__3072 (
            .O(N__23550),
            .I(buf_adcdata_vdc_14));
    LocalMux I__3071 (
            .O(N__23547),
            .I(buf_adcdata_vdc_14));
    CascadeMux I__3070 (
            .O(N__23542),
            .I(N__23538));
    CascadeMux I__3069 (
            .O(N__23541),
            .I(N__23535));
    InMux I__3068 (
            .O(N__23538),
            .I(N__23532));
    InMux I__3067 (
            .O(N__23535),
            .I(N__23529));
    LocalMux I__3066 (
            .O(N__23532),
            .I(buf_adcdata_vdc_22));
    LocalMux I__3065 (
            .O(N__23529),
            .I(buf_adcdata_vdc_22));
    CascadeMux I__3064 (
            .O(N__23524),
            .I(N__23520));
    CascadeMux I__3063 (
            .O(N__23523),
            .I(N__23517));
    InMux I__3062 (
            .O(N__23520),
            .I(N__23514));
    InMux I__3061 (
            .O(N__23517),
            .I(N__23511));
    LocalMux I__3060 (
            .O(N__23514),
            .I(N__23508));
    LocalMux I__3059 (
            .O(N__23511),
            .I(N__23505));
    Odrv4 I__3058 (
            .O(N__23508),
            .I(buf_adcdata_vdc_17));
    Odrv4 I__3057 (
            .O(N__23505),
            .I(buf_adcdata_vdc_17));
    InMux I__3056 (
            .O(N__23500),
            .I(N__23496));
    CascadeMux I__3055 (
            .O(N__23499),
            .I(N__23493));
    LocalMux I__3054 (
            .O(N__23496),
            .I(N__23490));
    InMux I__3053 (
            .O(N__23493),
            .I(N__23487));
    Odrv12 I__3052 (
            .O(N__23490),
            .I(buf_adcdata_vdc_0));
    LocalMux I__3051 (
            .O(N__23487),
            .I(buf_adcdata_vdc_0));
    InMux I__3050 (
            .O(N__23482),
            .I(N__23479));
    LocalMux I__3049 (
            .O(N__23479),
            .I(N__23474));
    InMux I__3048 (
            .O(N__23478),
            .I(N__23471));
    InMux I__3047 (
            .O(N__23477),
            .I(N__23468));
    Span4Mux_h I__3046 (
            .O(N__23474),
            .I(N__23463));
    LocalMux I__3045 (
            .O(N__23471),
            .I(N__23463));
    LocalMux I__3044 (
            .O(N__23468),
            .I(buf_adcdata_vac_0));
    Odrv4 I__3043 (
            .O(N__23463),
            .I(buf_adcdata_vac_0));
    InMux I__3042 (
            .O(N__23458),
            .I(N__23454));
    InMux I__3041 (
            .O(N__23457),
            .I(N__23451));
    LocalMux I__3040 (
            .O(N__23454),
            .I(N__23447));
    LocalMux I__3039 (
            .O(N__23451),
            .I(N__23444));
    InMux I__3038 (
            .O(N__23450),
            .I(N__23441));
    Span4Mux_v I__3037 (
            .O(N__23447),
            .I(N__23436));
    Span4Mux_v I__3036 (
            .O(N__23444),
            .I(N__23436));
    LocalMux I__3035 (
            .O(N__23441),
            .I(buf_adcdata_iac_0));
    Odrv4 I__3034 (
            .O(N__23436),
            .I(buf_adcdata_iac_0));
    CascadeMux I__3033 (
            .O(N__23431),
            .I(n19_adj_1477_cascade_));
    CascadeMux I__3032 (
            .O(N__23428),
            .I(N__23425));
    InMux I__3031 (
            .O(N__23425),
            .I(N__23422));
    LocalMux I__3030 (
            .O(N__23422),
            .I(N__23419));
    Span4Mux_h I__3029 (
            .O(N__23419),
            .I(N__23416));
    Span4Mux_h I__3028 (
            .O(N__23416),
            .I(N__23412));
    InMux I__3027 (
            .O(N__23415),
            .I(N__23409));
    Odrv4 I__3026 (
            .O(N__23412),
            .I(buf_readRTD_14));
    LocalMux I__3025 (
            .O(N__23409),
            .I(buf_readRTD_14));
    InMux I__3024 (
            .O(N__23404),
            .I(N__23401));
    LocalMux I__3023 (
            .O(N__23401),
            .I(n22141));
    InMux I__3022 (
            .O(N__23398),
            .I(N__23395));
    LocalMux I__3021 (
            .O(N__23395),
            .I(N__23392));
    Span4Mux_v I__3020 (
            .O(N__23392),
            .I(N__23388));
    CascadeMux I__3019 (
            .O(N__23391),
            .I(N__23385));
    Span4Mux_h I__3018 (
            .O(N__23388),
            .I(N__23382));
    InMux I__3017 (
            .O(N__23385),
            .I(N__23379));
    Odrv4 I__3016 (
            .O(N__23382),
            .I(buf_readRTD_10));
    LocalMux I__3015 (
            .O(N__23379),
            .I(buf_readRTD_10));
    CascadeMux I__3014 (
            .O(N__23374),
            .I(N__23371));
    InMux I__3013 (
            .O(N__23371),
            .I(N__23368));
    LocalMux I__3012 (
            .O(N__23368),
            .I(N__23364));
    CascadeMux I__3011 (
            .O(N__23367),
            .I(N__23361));
    Span4Mux_v I__3010 (
            .O(N__23364),
            .I(N__23358));
    InMux I__3009 (
            .O(N__23361),
            .I(N__23355));
    Odrv4 I__3008 (
            .O(N__23358),
            .I(buf_adcdata_vdc_21));
    LocalMux I__3007 (
            .O(N__23355),
            .I(buf_adcdata_vdc_21));
    InMux I__3006 (
            .O(N__23350),
            .I(N__23347));
    LocalMux I__3005 (
            .O(N__23347),
            .I(N__23344));
    Span4Mux_v I__3004 (
            .O(N__23344),
            .I(N__23340));
    CascadeMux I__3003 (
            .O(N__23343),
            .I(N__23337));
    Span4Mux_v I__3002 (
            .O(N__23340),
            .I(N__23334));
    InMux I__3001 (
            .O(N__23337),
            .I(N__23331));
    Odrv4 I__3000 (
            .O(N__23334),
            .I(buf_adcdata_vdc_13));
    LocalMux I__2999 (
            .O(N__23331),
            .I(buf_adcdata_vdc_13));
    InMux I__2998 (
            .O(N__23326),
            .I(N__23322));
    CascadeMux I__2997 (
            .O(N__23325),
            .I(N__23319));
    LocalMux I__2996 (
            .O(N__23322),
            .I(N__23316));
    InMux I__2995 (
            .O(N__23319),
            .I(N__23313));
    Odrv4 I__2994 (
            .O(N__23316),
            .I(buf_adcdata_vdc_16));
    LocalMux I__2993 (
            .O(N__23313),
            .I(buf_adcdata_vdc_16));
    InMux I__2992 (
            .O(N__23308),
            .I(N__23304));
    CascadeMux I__2991 (
            .O(N__23307),
            .I(N__23301));
    LocalMux I__2990 (
            .O(N__23304),
            .I(N__23298));
    InMux I__2989 (
            .O(N__23301),
            .I(N__23295));
    Odrv4 I__2988 (
            .O(N__23298),
            .I(buf_adcdata_vdc_2));
    LocalMux I__2987 (
            .O(N__23295),
            .I(buf_adcdata_vdc_2));
    InMux I__2986 (
            .O(N__23290),
            .I(N__23287));
    LocalMux I__2985 (
            .O(N__23287),
            .I(N__23283));
    CascadeMux I__2984 (
            .O(N__23286),
            .I(N__23280));
    Span4Mux_v I__2983 (
            .O(N__23283),
            .I(N__23277));
    InMux I__2982 (
            .O(N__23280),
            .I(N__23274));
    Odrv4 I__2981 (
            .O(N__23277),
            .I(buf_adcdata_vdc_19));
    LocalMux I__2980 (
            .O(N__23274),
            .I(buf_adcdata_vdc_19));
    CEMux I__2979 (
            .O(N__23269),
            .I(N__23266));
    LocalMux I__2978 (
            .O(N__23266),
            .I(N__23263));
    Odrv4 I__2977 (
            .O(N__23263),
            .I(\CLK_DDS.n9_adj_1386 ));
    InMux I__2976 (
            .O(N__23260),
            .I(\ADC_IAC.n19355 ));
    InMux I__2975 (
            .O(N__23257),
            .I(\ADC_IAC.n19356 ));
    CEMux I__2974 (
            .O(N__23254),
            .I(N__23251));
    LocalMux I__2973 (
            .O(N__23251),
            .I(N__23248));
    Span4Mux_v I__2972 (
            .O(N__23248),
            .I(N__23245));
    Span4Mux_h I__2971 (
            .O(N__23245),
            .I(N__23242));
    Odrv4 I__2970 (
            .O(N__23242),
            .I(\ADC_IAC.n12459 ));
    SRMux I__2969 (
            .O(N__23239),
            .I(N__23236));
    LocalMux I__2968 (
            .O(N__23236),
            .I(\ADC_IAC.n14791 ));
    InMux I__2967 (
            .O(N__23233),
            .I(N__23226));
    InMux I__2966 (
            .O(N__23232),
            .I(N__23219));
    InMux I__2965 (
            .O(N__23231),
            .I(N__23219));
    InMux I__2964 (
            .O(N__23230),
            .I(N__23219));
    InMux I__2963 (
            .O(N__23229),
            .I(N__23216));
    LocalMux I__2962 (
            .O(N__23226),
            .I(bit_cnt_0_adj_1449));
    LocalMux I__2961 (
            .O(N__23219),
            .I(bit_cnt_0_adj_1449));
    LocalMux I__2960 (
            .O(N__23216),
            .I(bit_cnt_0_adj_1449));
    CascadeMux I__2959 (
            .O(N__23209),
            .I(N__23206));
    InMux I__2958 (
            .O(N__23206),
            .I(N__23202));
    InMux I__2957 (
            .O(N__23205),
            .I(N__23199));
    LocalMux I__2956 (
            .O(N__23202),
            .I(N__23194));
    LocalMux I__2955 (
            .O(N__23199),
            .I(N__23194));
    Odrv4 I__2954 (
            .O(N__23194),
            .I(bit_cnt_3));
    InMux I__2953 (
            .O(N__23191),
            .I(N__23188));
    LocalMux I__2952 (
            .O(N__23188),
            .I(N__23185));
    Span4Mux_v I__2951 (
            .O(N__23185),
            .I(N__23182));
    Odrv4 I__2950 (
            .O(N__23182),
            .I(n21206));
    InMux I__2949 (
            .O(N__23179),
            .I(N__23176));
    LocalMux I__2948 (
            .O(N__23176),
            .I(N__23173));
    Span4Mux_v I__2947 (
            .O(N__23173),
            .I(N__23169));
    CascadeMux I__2946 (
            .O(N__23172),
            .I(N__23166));
    Span4Mux_v I__2945 (
            .O(N__23169),
            .I(N__23163));
    InMux I__2944 (
            .O(N__23166),
            .I(N__23160));
    Odrv4 I__2943 (
            .O(N__23163),
            .I(buf_adcdata_vdc_3));
    LocalMux I__2942 (
            .O(N__23160),
            .I(buf_adcdata_vdc_3));
    CascadeMux I__2941 (
            .O(N__23155),
            .I(\ADC_IAC.n12459_cascade_ ));
    InMux I__2940 (
            .O(N__23152),
            .I(bfn_7_19_0_));
    InMux I__2939 (
            .O(N__23149),
            .I(\ADC_IAC.n19350 ));
    InMux I__2938 (
            .O(N__23146),
            .I(\ADC_IAC.n19351 ));
    InMux I__2937 (
            .O(N__23143),
            .I(\ADC_IAC.n19352 ));
    InMux I__2936 (
            .O(N__23140),
            .I(\ADC_IAC.n19353 ));
    InMux I__2935 (
            .O(N__23137),
            .I(\ADC_IAC.n19354 ));
    InMux I__2934 (
            .O(N__23134),
            .I(N__23130));
    InMux I__2933 (
            .O(N__23133),
            .I(N__23127));
    LocalMux I__2932 (
            .O(N__23130),
            .I(\ADC_VAC.bit_cnt_2 ));
    LocalMux I__2931 (
            .O(N__23127),
            .I(\ADC_VAC.bit_cnt_2 ));
    InMux I__2930 (
            .O(N__23122),
            .I(\ADC_VAC.n19358 ));
    InMux I__2929 (
            .O(N__23119),
            .I(N__23115));
    InMux I__2928 (
            .O(N__23118),
            .I(N__23112));
    LocalMux I__2927 (
            .O(N__23115),
            .I(\ADC_VAC.bit_cnt_3 ));
    LocalMux I__2926 (
            .O(N__23112),
            .I(\ADC_VAC.bit_cnt_3 ));
    InMux I__2925 (
            .O(N__23107),
            .I(\ADC_VAC.n19359 ));
    InMux I__2924 (
            .O(N__23104),
            .I(N__23100));
    InMux I__2923 (
            .O(N__23103),
            .I(N__23097));
    LocalMux I__2922 (
            .O(N__23100),
            .I(N__23094));
    LocalMux I__2921 (
            .O(N__23097),
            .I(\ADC_VAC.bit_cnt_4 ));
    Odrv4 I__2920 (
            .O(N__23094),
            .I(\ADC_VAC.bit_cnt_4 ));
    InMux I__2919 (
            .O(N__23089),
            .I(\ADC_VAC.n19360 ));
    InMux I__2918 (
            .O(N__23086),
            .I(N__23082));
    InMux I__2917 (
            .O(N__23085),
            .I(N__23079));
    LocalMux I__2916 (
            .O(N__23082),
            .I(\ADC_VAC.bit_cnt_5 ));
    LocalMux I__2915 (
            .O(N__23079),
            .I(\ADC_VAC.bit_cnt_5 ));
    InMux I__2914 (
            .O(N__23074),
            .I(\ADC_VAC.n19361 ));
    InMux I__2913 (
            .O(N__23071),
            .I(N__23067));
    InMux I__2912 (
            .O(N__23070),
            .I(N__23064));
    LocalMux I__2911 (
            .O(N__23067),
            .I(\ADC_VAC.bit_cnt_6 ));
    LocalMux I__2910 (
            .O(N__23064),
            .I(\ADC_VAC.bit_cnt_6 ));
    InMux I__2909 (
            .O(N__23059),
            .I(\ADC_VAC.n19362 ));
    InMux I__2908 (
            .O(N__23056),
            .I(\ADC_VAC.n19363 ));
    InMux I__2907 (
            .O(N__23053),
            .I(N__23049));
    InMux I__2906 (
            .O(N__23052),
            .I(N__23046));
    LocalMux I__2905 (
            .O(N__23049),
            .I(\ADC_VAC.bit_cnt_7 ));
    LocalMux I__2904 (
            .O(N__23046),
            .I(\ADC_VAC.bit_cnt_7 ));
    CEMux I__2903 (
            .O(N__23041),
            .I(N__23038));
    LocalMux I__2902 (
            .O(N__23038),
            .I(N__23035));
    Span4Mux_v I__2901 (
            .O(N__23035),
            .I(N__23032));
    Odrv4 I__2900 (
            .O(N__23032),
            .I(\ADC_VAC.n12556 ));
    SRMux I__2899 (
            .O(N__23029),
            .I(N__23026));
    LocalMux I__2898 (
            .O(N__23026),
            .I(N__23023));
    Span4Mux_v I__2897 (
            .O(N__23023),
            .I(N__23020));
    Odrv4 I__2896 (
            .O(N__23020),
            .I(\ADC_VAC.n14829 ));
    CascadeMux I__2895 (
            .O(N__23017),
            .I(\ADC_VAC.n20747_cascade_ ));
    CascadeMux I__2894 (
            .O(N__23014),
            .I(\ADC_VAC.n20763_cascade_ ));
    CascadeMux I__2893 (
            .O(N__23011),
            .I(\ADC_VAC.n21031_cascade_ ));
    CEMux I__2892 (
            .O(N__23008),
            .I(N__23005));
    LocalMux I__2891 (
            .O(N__23005),
            .I(N__23002));
    Odrv4 I__2890 (
            .O(N__23002),
            .I(\ADC_VAC.n20668 ));
    CascadeMux I__2889 (
            .O(N__22999),
            .I(N__22995));
    InMux I__2888 (
            .O(N__22998),
            .I(N__22988));
    InMux I__2887 (
            .O(N__22995),
            .I(N__22988));
    InMux I__2886 (
            .O(N__22994),
            .I(N__22983));
    InMux I__2885 (
            .O(N__22993),
            .I(N__22983));
    LocalMux I__2884 (
            .O(N__22988),
            .I(N__22977));
    LocalMux I__2883 (
            .O(N__22983),
            .I(N__22977));
    InMux I__2882 (
            .O(N__22982),
            .I(N__22974));
    Span4Mux_v I__2881 (
            .O(N__22977),
            .I(N__22971));
    LocalMux I__2880 (
            .O(N__22974),
            .I(N__22968));
    Span4Mux_h I__2879 (
            .O(N__22971),
            .I(N__22965));
    Span4Mux_v I__2878 (
            .O(N__22968),
            .I(N__22962));
    Sp12to4 I__2877 (
            .O(N__22965),
            .I(N__22957));
    Sp12to4 I__2876 (
            .O(N__22962),
            .I(N__22957));
    Odrv12 I__2875 (
            .O(N__22957),
            .I(VAC_DRDY));
    CascadeMux I__2874 (
            .O(N__22954),
            .I(\ADC_VAC.n17_cascade_ ));
    CEMux I__2873 (
            .O(N__22951),
            .I(N__22948));
    LocalMux I__2872 (
            .O(N__22948),
            .I(N__22945));
    Odrv4 I__2871 (
            .O(N__22945),
            .I(\ADC_VAC.n12 ));
    InMux I__2870 (
            .O(N__22942),
            .I(N__22938));
    InMux I__2869 (
            .O(N__22941),
            .I(N__22935));
    LocalMux I__2868 (
            .O(N__22938),
            .I(\ADC_VAC.bit_cnt_0 ));
    LocalMux I__2867 (
            .O(N__22935),
            .I(\ADC_VAC.bit_cnt_0 ));
    InMux I__2866 (
            .O(N__22930),
            .I(bfn_7_17_0_));
    CascadeMux I__2865 (
            .O(N__22927),
            .I(N__22923));
    InMux I__2864 (
            .O(N__22926),
            .I(N__22920));
    InMux I__2863 (
            .O(N__22923),
            .I(N__22917));
    LocalMux I__2862 (
            .O(N__22920),
            .I(\ADC_VAC.bit_cnt_1 ));
    LocalMux I__2861 (
            .O(N__22917),
            .I(\ADC_VAC.bit_cnt_1 ));
    InMux I__2860 (
            .O(N__22912),
            .I(\ADC_VAC.n19357 ));
    CascadeMux I__2859 (
            .O(N__22909),
            .I(N__22906));
    InMux I__2858 (
            .O(N__22906),
            .I(N__22900));
    InMux I__2857 (
            .O(N__22905),
            .I(N__22900));
    LocalMux I__2856 (
            .O(N__22900),
            .I(cmd_rdadctmp_0_adj_1443));
    InMux I__2855 (
            .O(N__22897),
            .I(N__22891));
    InMux I__2854 (
            .O(N__22896),
            .I(N__22891));
    LocalMux I__2853 (
            .O(N__22891),
            .I(cmd_rdadctmp_1_adj_1442));
    InMux I__2852 (
            .O(N__22888),
            .I(N__22882));
    InMux I__2851 (
            .O(N__22887),
            .I(N__22882));
    LocalMux I__2850 (
            .O(N__22882),
            .I(cmd_rdadctmp_2_adj_1441));
    CascadeMux I__2849 (
            .O(N__22879),
            .I(N__22876));
    InMux I__2848 (
            .O(N__22876),
            .I(N__22872));
    InMux I__2847 (
            .O(N__22875),
            .I(N__22869));
    LocalMux I__2846 (
            .O(N__22872),
            .I(cmd_rdadctmp_3_adj_1440));
    LocalMux I__2845 (
            .O(N__22869),
            .I(cmd_rdadctmp_3_adj_1440));
    InMux I__2844 (
            .O(N__22864),
            .I(N__22861));
    LocalMux I__2843 (
            .O(N__22861),
            .I(N__22858));
    Odrv12 I__2842 (
            .O(N__22858),
            .I(n20573));
    CascadeMux I__2841 (
            .O(N__22855),
            .I(\ADC_VAC.n12556_cascade_ ));
    InMux I__2840 (
            .O(N__22852),
            .I(N__22849));
    LocalMux I__2839 (
            .O(N__22849),
            .I(\ADC_VAC.n20667 ));
    CascadeMux I__2838 (
            .O(N__22846),
            .I(N__22842));
    CascadeMux I__2837 (
            .O(N__22845),
            .I(N__22839));
    InMux I__2836 (
            .O(N__22842),
            .I(N__22835));
    InMux I__2835 (
            .O(N__22839),
            .I(N__22830));
    InMux I__2834 (
            .O(N__22838),
            .I(N__22830));
    LocalMux I__2833 (
            .O(N__22835),
            .I(cmd_rdadctmp_11_adj_1432));
    LocalMux I__2832 (
            .O(N__22830),
            .I(cmd_rdadctmp_11_adj_1432));
    InMux I__2831 (
            .O(N__22825),
            .I(N__22822));
    LocalMux I__2830 (
            .O(N__22822),
            .I(N__22819));
    Span4Mux_v I__2829 (
            .O(N__22819),
            .I(N__22815));
    InMux I__2828 (
            .O(N__22818),
            .I(N__22812));
    Odrv4 I__2827 (
            .O(N__22815),
            .I(cmd_rdadctmp_7_adj_1436));
    LocalMux I__2826 (
            .O(N__22812),
            .I(cmd_rdadctmp_7_adj_1436));
    CascadeMux I__2825 (
            .O(N__22807),
            .I(N__22804));
    InMux I__2824 (
            .O(N__22804),
            .I(N__22800));
    CascadeMux I__2823 (
            .O(N__22803),
            .I(N__22797));
    LocalMux I__2822 (
            .O(N__22800),
            .I(N__22793));
    InMux I__2821 (
            .O(N__22797),
            .I(N__22788));
    InMux I__2820 (
            .O(N__22796),
            .I(N__22788));
    Odrv4 I__2819 (
            .O(N__22793),
            .I(cmd_rdadctmp_8_adj_1435));
    LocalMux I__2818 (
            .O(N__22788),
            .I(cmd_rdadctmp_8_adj_1435));
    CascadeMux I__2817 (
            .O(N__22783),
            .I(N__22779));
    CascadeMux I__2816 (
            .O(N__22782),
            .I(N__22776));
    InMux I__2815 (
            .O(N__22779),
            .I(N__22768));
    InMux I__2814 (
            .O(N__22776),
            .I(N__22768));
    InMux I__2813 (
            .O(N__22775),
            .I(N__22768));
    LocalMux I__2812 (
            .O(N__22768),
            .I(cmd_rdadctmp_9_adj_1434));
    CascadeMux I__2811 (
            .O(N__22765),
            .I(N__22762));
    InMux I__2810 (
            .O(N__22762),
            .I(N__22759));
    LocalMux I__2809 (
            .O(N__22759),
            .I(N__22756));
    Span4Mux_h I__2808 (
            .O(N__22756),
            .I(N__22753));
    Sp12to4 I__2807 (
            .O(N__22753),
            .I(N__22750));
    Odrv12 I__2806 (
            .O(N__22750),
            .I(VAC_MISO));
    InMux I__2805 (
            .O(N__22747),
            .I(N__22744));
    LocalMux I__2804 (
            .O(N__22744),
            .I(n21973));
    InMux I__2803 (
            .O(N__22741),
            .I(N__22734));
    InMux I__2802 (
            .O(N__22740),
            .I(N__22734));
    InMux I__2801 (
            .O(N__22739),
            .I(N__22731));
    LocalMux I__2800 (
            .O(N__22734),
            .I(cmd_rdadctmp_17_adj_1426));
    LocalMux I__2799 (
            .O(N__22731),
            .I(cmd_rdadctmp_17_adj_1426));
    InMux I__2798 (
            .O(N__22726),
            .I(N__22721));
    InMux I__2797 (
            .O(N__22725),
            .I(N__22716));
    InMux I__2796 (
            .O(N__22724),
            .I(N__22716));
    LocalMux I__2795 (
            .O(N__22721),
            .I(cmd_rdadctmp_16_adj_1427));
    LocalMux I__2794 (
            .O(N__22716),
            .I(cmd_rdadctmp_16_adj_1427));
    InMux I__2793 (
            .O(N__22711),
            .I(N__22708));
    LocalMux I__2792 (
            .O(N__22708),
            .I(N__22705));
    Span4Mux_h I__2791 (
            .O(N__22705),
            .I(N__22700));
    InMux I__2790 (
            .O(N__22704),
            .I(N__22697));
    InMux I__2789 (
            .O(N__22703),
            .I(N__22694));
    Sp12to4 I__2788 (
            .O(N__22700),
            .I(N__22691));
    LocalMux I__2787 (
            .O(N__22697),
            .I(N__22688));
    LocalMux I__2786 (
            .O(N__22694),
            .I(buf_adcdata_vac_22));
    Odrv12 I__2785 (
            .O(N__22691),
            .I(buf_adcdata_vac_22));
    Odrv4 I__2784 (
            .O(N__22688),
            .I(buf_adcdata_vac_22));
    InMux I__2783 (
            .O(N__22681),
            .I(N__22678));
    LocalMux I__2782 (
            .O(N__22678),
            .I(N__22674));
    InMux I__2781 (
            .O(N__22677),
            .I(N__22670));
    Span4Mux_v I__2780 (
            .O(N__22674),
            .I(N__22667));
    InMux I__2779 (
            .O(N__22673),
            .I(N__22664));
    LocalMux I__2778 (
            .O(N__22670),
            .I(buf_adcdata_vac_14));
    Odrv4 I__2777 (
            .O(N__22667),
            .I(buf_adcdata_vac_14));
    LocalMux I__2776 (
            .O(N__22664),
            .I(buf_adcdata_vac_14));
    InMux I__2775 (
            .O(N__22657),
            .I(N__22653));
    CascadeMux I__2774 (
            .O(N__22656),
            .I(N__22649));
    LocalMux I__2773 (
            .O(N__22653),
            .I(N__22646));
    InMux I__2772 (
            .O(N__22652),
            .I(N__22643));
    InMux I__2771 (
            .O(N__22649),
            .I(N__22640));
    Span4Mux_h I__2770 (
            .O(N__22646),
            .I(N__22637));
    LocalMux I__2769 (
            .O(N__22643),
            .I(N__22634));
    LocalMux I__2768 (
            .O(N__22640),
            .I(buf_adcdata_vac_17));
    Odrv4 I__2767 (
            .O(N__22637),
            .I(buf_adcdata_vac_17));
    Odrv12 I__2766 (
            .O(N__22634),
            .I(buf_adcdata_vac_17));
    CascadeMux I__2765 (
            .O(N__22627),
            .I(N__22623));
    CascadeMux I__2764 (
            .O(N__22626),
            .I(N__22620));
    InMux I__2763 (
            .O(N__22623),
            .I(N__22614));
    InMux I__2762 (
            .O(N__22620),
            .I(N__22614));
    InMux I__2761 (
            .O(N__22619),
            .I(N__22611));
    LocalMux I__2760 (
            .O(N__22614),
            .I(cmd_rdadctmp_30_adj_1413));
    LocalMux I__2759 (
            .O(N__22611),
            .I(cmd_rdadctmp_30_adj_1413));
    InMux I__2758 (
            .O(N__22606),
            .I(N__22600));
    InMux I__2757 (
            .O(N__22605),
            .I(N__22600));
    LocalMux I__2756 (
            .O(N__22600),
            .I(cmd_rdadctmp_31_adj_1412));
    CascadeMux I__2755 (
            .O(N__22597),
            .I(N__22592));
    InMux I__2754 (
            .O(N__22596),
            .I(N__22589));
    InMux I__2753 (
            .O(N__22595),
            .I(N__22586));
    InMux I__2752 (
            .O(N__22592),
            .I(N__22583));
    LocalMux I__2751 (
            .O(N__22589),
            .I(N__22580));
    LocalMux I__2750 (
            .O(N__22586),
            .I(N__22577));
    LocalMux I__2749 (
            .O(N__22583),
            .I(buf_adcdata_vac_16));
    Odrv4 I__2748 (
            .O(N__22580),
            .I(buf_adcdata_vac_16));
    Odrv12 I__2747 (
            .O(N__22577),
            .I(buf_adcdata_vac_16));
    CascadeMux I__2746 (
            .O(N__22570),
            .I(N__22567));
    InMux I__2745 (
            .O(N__22567),
            .I(N__22563));
    CascadeMux I__2744 (
            .O(N__22566),
            .I(N__22560));
    LocalMux I__2743 (
            .O(N__22563),
            .I(N__22556));
    InMux I__2742 (
            .O(N__22560),
            .I(N__22553));
    InMux I__2741 (
            .O(N__22559),
            .I(N__22550));
    Odrv12 I__2740 (
            .O(N__22556),
            .I(cmd_rdadctmp_10_adj_1433));
    LocalMux I__2739 (
            .O(N__22553),
            .I(cmd_rdadctmp_10_adj_1433));
    LocalMux I__2738 (
            .O(N__22550),
            .I(cmd_rdadctmp_10_adj_1433));
    CascadeMux I__2737 (
            .O(N__22543),
            .I(n22183_cascade_));
    CascadeMux I__2736 (
            .O(N__22540),
            .I(N__22537));
    InMux I__2735 (
            .O(N__22537),
            .I(N__22534));
    LocalMux I__2734 (
            .O(N__22534),
            .I(N__22531));
    Span4Mux_v I__2733 (
            .O(N__22531),
            .I(N__22528));
    Odrv4 I__2732 (
            .O(N__22528),
            .I(buf_data_iac_2));
    CascadeMux I__2731 (
            .O(N__22525),
            .I(N__22522));
    InMux I__2730 (
            .O(N__22522),
            .I(N__22519));
    LocalMux I__2729 (
            .O(N__22519),
            .I(N__22515));
    CascadeMux I__2728 (
            .O(N__22518),
            .I(N__22512));
    Span4Mux_v I__2727 (
            .O(N__22515),
            .I(N__22509));
    InMux I__2726 (
            .O(N__22512),
            .I(N__22506));
    Odrv4 I__2725 (
            .O(N__22509),
            .I(buf_readRTD_13));
    LocalMux I__2724 (
            .O(N__22506),
            .I(buf_readRTD_13));
    InMux I__2723 (
            .O(N__22501),
            .I(N__22498));
    LocalMux I__2722 (
            .O(N__22498),
            .I(n22153));
    InMux I__2721 (
            .O(N__22495),
            .I(N__22492));
    LocalMux I__2720 (
            .O(N__22492),
            .I(N__22487));
    InMux I__2719 (
            .O(N__22491),
            .I(N__22484));
    InMux I__2718 (
            .O(N__22490),
            .I(N__22481));
    Span4Mux_v I__2717 (
            .O(N__22487),
            .I(N__22478));
    LocalMux I__2716 (
            .O(N__22484),
            .I(N__22475));
    LocalMux I__2715 (
            .O(N__22481),
            .I(buf_adcdata_iac_2));
    Odrv4 I__2714 (
            .O(N__22478),
            .I(buf_adcdata_iac_2));
    Odrv12 I__2713 (
            .O(N__22475),
            .I(buf_adcdata_iac_2));
    CascadeMux I__2712 (
            .O(N__22468),
            .I(n19_adj_1613_cascade_));
    InMux I__2711 (
            .O(N__22465),
            .I(N__22462));
    LocalMux I__2710 (
            .O(N__22462),
            .I(n22_adj_1614));
    CascadeMux I__2709 (
            .O(N__22459),
            .I(N__22456));
    InMux I__2708 (
            .O(N__22456),
            .I(N__22453));
    LocalMux I__2707 (
            .O(N__22453),
            .I(N__22449));
    CascadeMux I__2706 (
            .O(N__22452),
            .I(N__22446));
    Span4Mux_v I__2705 (
            .O(N__22449),
            .I(N__22443));
    InMux I__2704 (
            .O(N__22446),
            .I(N__22440));
    Odrv4 I__2703 (
            .O(N__22443),
            .I(buf_readRTD_15));
    LocalMux I__2702 (
            .O(N__22440),
            .I(buf_readRTD_15));
    InMux I__2701 (
            .O(N__22435),
            .I(N__22432));
    LocalMux I__2700 (
            .O(N__22432),
            .I(N__22429));
    Span4Mux_h I__2699 (
            .O(N__22429),
            .I(N__22426));
    Span4Mux_v I__2698 (
            .O(N__22426),
            .I(N__22421));
    InMux I__2697 (
            .O(N__22425),
            .I(N__22416));
    InMux I__2696 (
            .O(N__22424),
            .I(N__22416));
    Odrv4 I__2695 (
            .O(N__22421),
            .I(buf_adcdata_vac_2));
    LocalMux I__2694 (
            .O(N__22416),
            .I(buf_adcdata_vac_2));
    CascadeMux I__2693 (
            .O(N__22411),
            .I(N__22405));
    CascadeMux I__2692 (
            .O(N__22410),
            .I(N__22399));
    CascadeMux I__2691 (
            .O(N__22409),
            .I(N__22396));
    CascadeMux I__2690 (
            .O(N__22408),
            .I(N__22390));
    InMux I__2689 (
            .O(N__22405),
            .I(N__22384));
    InMux I__2688 (
            .O(N__22404),
            .I(N__22381));
    InMux I__2687 (
            .O(N__22403),
            .I(N__22378));
    CascadeMux I__2686 (
            .O(N__22402),
            .I(N__22375));
    InMux I__2685 (
            .O(N__22399),
            .I(N__22362));
    InMux I__2684 (
            .O(N__22396),
            .I(N__22362));
    InMux I__2683 (
            .O(N__22395),
            .I(N__22362));
    InMux I__2682 (
            .O(N__22394),
            .I(N__22362));
    InMux I__2681 (
            .O(N__22393),
            .I(N__22362));
    InMux I__2680 (
            .O(N__22390),
            .I(N__22362));
    CascadeMux I__2679 (
            .O(N__22389),
            .I(N__22356));
    InMux I__2678 (
            .O(N__22388),
            .I(N__22345));
    InMux I__2677 (
            .O(N__22387),
            .I(N__22345));
    LocalMux I__2676 (
            .O(N__22384),
            .I(N__22342));
    LocalMux I__2675 (
            .O(N__22381),
            .I(N__22337));
    LocalMux I__2674 (
            .O(N__22378),
            .I(N__22337));
    InMux I__2673 (
            .O(N__22375),
            .I(N__22334));
    LocalMux I__2672 (
            .O(N__22362),
            .I(N__22330));
    InMux I__2671 (
            .O(N__22361),
            .I(N__22325));
    InMux I__2670 (
            .O(N__22360),
            .I(N__22325));
    InMux I__2669 (
            .O(N__22359),
            .I(N__22316));
    InMux I__2668 (
            .O(N__22356),
            .I(N__22316));
    InMux I__2667 (
            .O(N__22355),
            .I(N__22316));
    InMux I__2666 (
            .O(N__22354),
            .I(N__22313));
    InMux I__2665 (
            .O(N__22353),
            .I(N__22310));
    InMux I__2664 (
            .O(N__22352),
            .I(N__22303));
    InMux I__2663 (
            .O(N__22351),
            .I(N__22303));
    InMux I__2662 (
            .O(N__22350),
            .I(N__22303));
    LocalMux I__2661 (
            .O(N__22345),
            .I(N__22294));
    Span4Mux_h I__2660 (
            .O(N__22342),
            .I(N__22294));
    Span4Mux_v I__2659 (
            .O(N__22337),
            .I(N__22294));
    LocalMux I__2658 (
            .O(N__22334),
            .I(N__22294));
    InMux I__2657 (
            .O(N__22333),
            .I(N__22291));
    Span4Mux_h I__2656 (
            .O(N__22330),
            .I(N__22286));
    LocalMux I__2655 (
            .O(N__22325),
            .I(N__22286));
    InMux I__2654 (
            .O(N__22324),
            .I(N__22281));
    InMux I__2653 (
            .O(N__22323),
            .I(N__22281));
    LocalMux I__2652 (
            .O(N__22316),
            .I(N__22278));
    LocalMux I__2651 (
            .O(N__22313),
            .I(\RTD.adc_state_3 ));
    LocalMux I__2650 (
            .O(N__22310),
            .I(\RTD.adc_state_3 ));
    LocalMux I__2649 (
            .O(N__22303),
            .I(\RTD.adc_state_3 ));
    Odrv4 I__2648 (
            .O(N__22294),
            .I(\RTD.adc_state_3 ));
    LocalMux I__2647 (
            .O(N__22291),
            .I(\RTD.adc_state_3 ));
    Odrv4 I__2646 (
            .O(N__22286),
            .I(\RTD.adc_state_3 ));
    LocalMux I__2645 (
            .O(N__22281),
            .I(\RTD.adc_state_3 ));
    Odrv4 I__2644 (
            .O(N__22278),
            .I(\RTD.adc_state_3 ));
    CascadeMux I__2643 (
            .O(N__22261),
            .I(N__22249));
    InMux I__2642 (
            .O(N__22260),
            .I(N__22243));
    InMux I__2641 (
            .O(N__22259),
            .I(N__22240));
    InMux I__2640 (
            .O(N__22258),
            .I(N__22237));
    InMux I__2639 (
            .O(N__22257),
            .I(N__22224));
    InMux I__2638 (
            .O(N__22256),
            .I(N__22224));
    InMux I__2637 (
            .O(N__22255),
            .I(N__22224));
    InMux I__2636 (
            .O(N__22254),
            .I(N__22224));
    InMux I__2635 (
            .O(N__22253),
            .I(N__22224));
    InMux I__2634 (
            .O(N__22252),
            .I(N__22224));
    InMux I__2633 (
            .O(N__22249),
            .I(N__22212));
    InMux I__2632 (
            .O(N__22248),
            .I(N__22212));
    InMux I__2631 (
            .O(N__22247),
            .I(N__22212));
    InMux I__2630 (
            .O(N__22246),
            .I(N__22209));
    LocalMux I__2629 (
            .O(N__22243),
            .I(N__22204));
    LocalMux I__2628 (
            .O(N__22240),
            .I(N__22204));
    LocalMux I__2627 (
            .O(N__22237),
            .I(N__22199));
    LocalMux I__2626 (
            .O(N__22224),
            .I(N__22199));
    InMux I__2625 (
            .O(N__22223),
            .I(N__22196));
    InMux I__2624 (
            .O(N__22222),
            .I(N__22187));
    InMux I__2623 (
            .O(N__22221),
            .I(N__22182));
    InMux I__2622 (
            .O(N__22220),
            .I(N__22182));
    InMux I__2621 (
            .O(N__22219),
            .I(N__22179));
    LocalMux I__2620 (
            .O(N__22212),
            .I(N__22176));
    LocalMux I__2619 (
            .O(N__22209),
            .I(N__22169));
    Span4Mux_v I__2618 (
            .O(N__22204),
            .I(N__22169));
    Span4Mux_v I__2617 (
            .O(N__22199),
            .I(N__22169));
    LocalMux I__2616 (
            .O(N__22196),
            .I(N__22166));
    InMux I__2615 (
            .O(N__22195),
            .I(N__22163));
    InMux I__2614 (
            .O(N__22194),
            .I(N__22158));
    InMux I__2613 (
            .O(N__22193),
            .I(N__22158));
    InMux I__2612 (
            .O(N__22192),
            .I(N__22151));
    InMux I__2611 (
            .O(N__22191),
            .I(N__22151));
    InMux I__2610 (
            .O(N__22190),
            .I(N__22151));
    LocalMux I__2609 (
            .O(N__22187),
            .I(\RTD.adc_state_1 ));
    LocalMux I__2608 (
            .O(N__22182),
            .I(\RTD.adc_state_1 ));
    LocalMux I__2607 (
            .O(N__22179),
            .I(\RTD.adc_state_1 ));
    Odrv4 I__2606 (
            .O(N__22176),
            .I(\RTD.adc_state_1 ));
    Odrv4 I__2605 (
            .O(N__22169),
            .I(\RTD.adc_state_1 ));
    Odrv4 I__2604 (
            .O(N__22166),
            .I(\RTD.adc_state_1 ));
    LocalMux I__2603 (
            .O(N__22163),
            .I(\RTD.adc_state_1 ));
    LocalMux I__2602 (
            .O(N__22158),
            .I(\RTD.adc_state_1 ));
    LocalMux I__2601 (
            .O(N__22151),
            .I(\RTD.adc_state_1 ));
    CascadeMux I__2600 (
            .O(N__22132),
            .I(N__22110));
    CascadeMux I__2599 (
            .O(N__22131),
            .I(N__22106));
    CascadeMux I__2598 (
            .O(N__22130),
            .I(N__22096));
    InMux I__2597 (
            .O(N__22129),
            .I(N__22088));
    InMux I__2596 (
            .O(N__22128),
            .I(N__22088));
    InMux I__2595 (
            .O(N__22127),
            .I(N__22085));
    InMux I__2594 (
            .O(N__22126),
            .I(N__22076));
    InMux I__2593 (
            .O(N__22125),
            .I(N__22076));
    InMux I__2592 (
            .O(N__22124),
            .I(N__22076));
    InMux I__2591 (
            .O(N__22123),
            .I(N__22076));
    InMux I__2590 (
            .O(N__22122),
            .I(N__22069));
    InMux I__2589 (
            .O(N__22121),
            .I(N__22069));
    InMux I__2588 (
            .O(N__22120),
            .I(N__22069));
    InMux I__2587 (
            .O(N__22119),
            .I(N__22064));
    InMux I__2586 (
            .O(N__22118),
            .I(N__22064));
    InMux I__2585 (
            .O(N__22117),
            .I(N__22057));
    InMux I__2584 (
            .O(N__22116),
            .I(N__22057));
    InMux I__2583 (
            .O(N__22115),
            .I(N__22057));
    InMux I__2582 (
            .O(N__22114),
            .I(N__22044));
    InMux I__2581 (
            .O(N__22113),
            .I(N__22044));
    InMux I__2580 (
            .O(N__22110),
            .I(N__22044));
    InMux I__2579 (
            .O(N__22109),
            .I(N__22044));
    InMux I__2578 (
            .O(N__22106),
            .I(N__22044));
    InMux I__2577 (
            .O(N__22105),
            .I(N__22044));
    InMux I__2576 (
            .O(N__22104),
            .I(N__22041));
    InMux I__2575 (
            .O(N__22103),
            .I(N__22038));
    InMux I__2574 (
            .O(N__22102),
            .I(N__22027));
    InMux I__2573 (
            .O(N__22101),
            .I(N__22018));
    InMux I__2572 (
            .O(N__22100),
            .I(N__22018));
    InMux I__2571 (
            .O(N__22099),
            .I(N__22018));
    InMux I__2570 (
            .O(N__22096),
            .I(N__22015));
    InMux I__2569 (
            .O(N__22095),
            .I(N__22008));
    InMux I__2568 (
            .O(N__22094),
            .I(N__22008));
    InMux I__2567 (
            .O(N__22093),
            .I(N__22008));
    LocalMux I__2566 (
            .O(N__22088),
            .I(N__21999));
    LocalMux I__2565 (
            .O(N__22085),
            .I(N__21999));
    LocalMux I__2564 (
            .O(N__22076),
            .I(N__21999));
    LocalMux I__2563 (
            .O(N__22069),
            .I(N__21999));
    LocalMux I__2562 (
            .O(N__22064),
            .I(N__21992));
    LocalMux I__2561 (
            .O(N__22057),
            .I(N__21992));
    LocalMux I__2560 (
            .O(N__22044),
            .I(N__21992));
    LocalMux I__2559 (
            .O(N__22041),
            .I(N__21984));
    LocalMux I__2558 (
            .O(N__22038),
            .I(N__21984));
    InMux I__2557 (
            .O(N__22037),
            .I(N__21968));
    InMux I__2556 (
            .O(N__22036),
            .I(N__21968));
    InMux I__2555 (
            .O(N__22035),
            .I(N__21968));
    InMux I__2554 (
            .O(N__22034),
            .I(N__21968));
    InMux I__2553 (
            .O(N__22033),
            .I(N__21968));
    InMux I__2552 (
            .O(N__22032),
            .I(N__21968));
    InMux I__2551 (
            .O(N__22031),
            .I(N__21968));
    InMux I__2550 (
            .O(N__22030),
            .I(N__21965));
    LocalMux I__2549 (
            .O(N__22027),
            .I(N__21962));
    InMux I__2548 (
            .O(N__22026),
            .I(N__21959));
    InMux I__2547 (
            .O(N__22025),
            .I(N__21956));
    LocalMux I__2546 (
            .O(N__22018),
            .I(N__21953));
    LocalMux I__2545 (
            .O(N__22015),
            .I(N__21944));
    LocalMux I__2544 (
            .O(N__22008),
            .I(N__21944));
    Span4Mux_v I__2543 (
            .O(N__21999),
            .I(N__21944));
    Span4Mux_v I__2542 (
            .O(N__21992),
            .I(N__21944));
    InMux I__2541 (
            .O(N__21991),
            .I(N__21937));
    InMux I__2540 (
            .O(N__21990),
            .I(N__21937));
    InMux I__2539 (
            .O(N__21989),
            .I(N__21937));
    Span4Mux_h I__2538 (
            .O(N__21984),
            .I(N__21934));
    InMux I__2537 (
            .O(N__21983),
            .I(N__21931));
    LocalMux I__2536 (
            .O(N__21968),
            .I(adc_state_2_adj_1474));
    LocalMux I__2535 (
            .O(N__21965),
            .I(adc_state_2_adj_1474));
    Odrv4 I__2534 (
            .O(N__21962),
            .I(adc_state_2_adj_1474));
    LocalMux I__2533 (
            .O(N__21959),
            .I(adc_state_2_adj_1474));
    LocalMux I__2532 (
            .O(N__21956),
            .I(adc_state_2_adj_1474));
    Odrv4 I__2531 (
            .O(N__21953),
            .I(adc_state_2_adj_1474));
    Odrv4 I__2530 (
            .O(N__21944),
            .I(adc_state_2_adj_1474));
    LocalMux I__2529 (
            .O(N__21937),
            .I(adc_state_2_adj_1474));
    Odrv4 I__2528 (
            .O(N__21934),
            .I(adc_state_2_adj_1474));
    LocalMux I__2527 (
            .O(N__21931),
            .I(adc_state_2_adj_1474));
    CascadeMux I__2526 (
            .O(N__21910),
            .I(N__21907));
    InMux I__2525 (
            .O(N__21907),
            .I(N__21904));
    LocalMux I__2524 (
            .O(N__21904),
            .I(N__21900));
    InMux I__2523 (
            .O(N__21903),
            .I(N__21897));
    Span12Mux_v I__2522 (
            .O(N__21900),
            .I(N__21892));
    LocalMux I__2521 (
            .O(N__21897),
            .I(N__21892));
    Odrv12 I__2520 (
            .O(N__21892),
            .I(\RTD.n20487 ));
    InMux I__2519 (
            .O(N__21889),
            .I(N__21886));
    LocalMux I__2518 (
            .O(N__21886),
            .I(N__21883));
    Span4Mux_h I__2517 (
            .O(N__21883),
            .I(N__21880));
    Span4Mux_v I__2516 (
            .O(N__21880),
            .I(N__21877));
    Odrv4 I__2515 (
            .O(N__21877),
            .I(buf_data_iac_22));
    IoInMux I__2514 (
            .O(N__21874),
            .I(N__21871));
    LocalMux I__2513 (
            .O(N__21871),
            .I(N__21868));
    Span12Mux_s6_v I__2512 (
            .O(N__21868),
            .I(N__21864));
    InMux I__2511 (
            .O(N__21867),
            .I(N__21861));
    Odrv12 I__2510 (
            .O(N__21864),
            .I(DDS_MOSI1));
    LocalMux I__2509 (
            .O(N__21861),
            .I(DDS_MOSI1));
    InMux I__2508 (
            .O(N__21856),
            .I(N__21853));
    LocalMux I__2507 (
            .O(N__21853),
            .I(N__21849));
    InMux I__2506 (
            .O(N__21852),
            .I(N__21846));
    Span4Mux_v I__2505 (
            .O(N__21849),
            .I(N__21843));
    LocalMux I__2504 (
            .O(N__21846),
            .I(N__21840));
    Span4Mux_v I__2503 (
            .O(N__21843),
            .I(N__21834));
    Span4Mux_h I__2502 (
            .O(N__21840),
            .I(N__21834));
    InMux I__2501 (
            .O(N__21839),
            .I(N__21831));
    Sp12to4 I__2500 (
            .O(N__21834),
            .I(N__21828));
    LocalMux I__2499 (
            .O(N__21831),
            .I(buf_adcdata_vac_21));
    Odrv12 I__2498 (
            .O(N__21828),
            .I(buf_adcdata_vac_21));
    CascadeMux I__2497 (
            .O(N__21823),
            .I(N__21820));
    InMux I__2496 (
            .O(N__21820),
            .I(N__21817));
    LocalMux I__2495 (
            .O(N__21817),
            .I(N__21814));
    Span4Mux_h I__2494 (
            .O(N__21814),
            .I(N__21810));
    InMux I__2493 (
            .O(N__21813),
            .I(N__21807));
    Odrv4 I__2492 (
            .O(N__21810),
            .I(buf_readRTD_8));
    LocalMux I__2491 (
            .O(N__21807),
            .I(buf_readRTD_8));
    CascadeMux I__2490 (
            .O(N__21802),
            .I(N__21798));
    CascadeMux I__2489 (
            .O(N__21801),
            .I(N__21795));
    InMux I__2488 (
            .O(N__21798),
            .I(N__21791));
    InMux I__2487 (
            .O(N__21795),
            .I(N__21786));
    InMux I__2486 (
            .O(N__21794),
            .I(N__21786));
    LocalMux I__2485 (
            .O(N__21791),
            .I(cmd_rdadctmp_20));
    LocalMux I__2484 (
            .O(N__21786),
            .I(cmd_rdadctmp_20));
    CascadeMux I__2483 (
            .O(N__21781),
            .I(N__21778));
    InMux I__2482 (
            .O(N__21778),
            .I(N__21773));
    InMux I__2481 (
            .O(N__21777),
            .I(N__21770));
    InMux I__2480 (
            .O(N__21776),
            .I(N__21767));
    LocalMux I__2479 (
            .O(N__21773),
            .I(cmd_rdadctmp_21));
    LocalMux I__2478 (
            .O(N__21770),
            .I(cmd_rdadctmp_21));
    LocalMux I__2477 (
            .O(N__21767),
            .I(cmd_rdadctmp_21));
    CascadeMux I__2476 (
            .O(N__21760),
            .I(N__21756));
    CascadeMux I__2475 (
            .O(N__21759),
            .I(N__21753));
    InMux I__2474 (
            .O(N__21756),
            .I(N__21749));
    InMux I__2473 (
            .O(N__21753),
            .I(N__21746));
    InMux I__2472 (
            .O(N__21752),
            .I(N__21743));
    LocalMux I__2471 (
            .O(N__21749),
            .I(cmd_rdadctmp_19));
    LocalMux I__2470 (
            .O(N__21746),
            .I(cmd_rdadctmp_19));
    LocalMux I__2469 (
            .O(N__21743),
            .I(cmd_rdadctmp_19));
    CascadeMux I__2468 (
            .O(N__21736),
            .I(N__21733));
    InMux I__2467 (
            .O(N__21733),
            .I(N__21729));
    CascadeMux I__2466 (
            .O(N__21732),
            .I(N__21726));
    LocalMux I__2465 (
            .O(N__21729),
            .I(N__21722));
    InMux I__2464 (
            .O(N__21726),
            .I(N__21719));
    InMux I__2463 (
            .O(N__21725),
            .I(N__21716));
    Odrv4 I__2462 (
            .O(N__21722),
            .I(cmd_rdadctmp_18));
    LocalMux I__2461 (
            .O(N__21719),
            .I(cmd_rdadctmp_18));
    LocalMux I__2460 (
            .O(N__21716),
            .I(cmd_rdadctmp_18));
    InMux I__2459 (
            .O(N__21709),
            .I(N__21706));
    LocalMux I__2458 (
            .O(N__21706),
            .I(N__21703));
    Odrv4 I__2457 (
            .O(N__21703),
            .I(buf_data_iac_11));
    CascadeMux I__2456 (
            .O(N__21700),
            .I(N__21697));
    InMux I__2455 (
            .O(N__21697),
            .I(N__21692));
    InMux I__2454 (
            .O(N__21696),
            .I(N__21687));
    InMux I__2453 (
            .O(N__21695),
            .I(N__21687));
    LocalMux I__2452 (
            .O(N__21692),
            .I(N__21684));
    LocalMux I__2451 (
            .O(N__21687),
            .I(N__21681));
    Odrv4 I__2450 (
            .O(N__21684),
            .I(cmd_rdadctmp_17));
    Odrv4 I__2449 (
            .O(N__21681),
            .I(cmd_rdadctmp_17));
    InMux I__2448 (
            .O(N__21676),
            .I(N__21673));
    LocalMux I__2447 (
            .O(N__21673),
            .I(N__21668));
    InMux I__2446 (
            .O(N__21672),
            .I(N__21665));
    InMux I__2445 (
            .O(N__21671),
            .I(N__21662));
    Span4Mux_h I__2444 (
            .O(N__21668),
            .I(N__21659));
    LocalMux I__2443 (
            .O(N__21665),
            .I(N__21656));
    LocalMux I__2442 (
            .O(N__21662),
            .I(buf_adcdata_iac_9));
    Odrv4 I__2441 (
            .O(N__21659),
            .I(buf_adcdata_iac_9));
    Odrv12 I__2440 (
            .O(N__21656),
            .I(buf_adcdata_iac_9));
    IoInMux I__2439 (
            .O(N__21649),
            .I(N__21646));
    LocalMux I__2438 (
            .O(N__21646),
            .I(N__21643));
    Span4Mux_s2_v I__2437 (
            .O(N__21643),
            .I(N__21640));
    Span4Mux_v I__2436 (
            .O(N__21640),
            .I(N__21637));
    Span4Mux_h I__2435 (
            .O(N__21637),
            .I(N__21634));
    Odrv4 I__2434 (
            .O(N__21634),
            .I(DDS_MCLK1));
    IoInMux I__2433 (
            .O(N__21631),
            .I(N__21628));
    LocalMux I__2432 (
            .O(N__21628),
            .I(N__21625));
    Span4Mux_s3_v I__2431 (
            .O(N__21625),
            .I(N__21622));
    Span4Mux_v I__2430 (
            .O(N__21622),
            .I(N__21619));
    Span4Mux_h I__2429 (
            .O(N__21619),
            .I(N__21616));
    Odrv4 I__2428 (
            .O(N__21616),
            .I(DDS_CS1));
    IoInMux I__2427 (
            .O(N__21613),
            .I(N__21610));
    LocalMux I__2426 (
            .O(N__21610),
            .I(N__21607));
    IoSpan4Mux I__2425 (
            .O(N__21607),
            .I(N__21604));
    Span4Mux_s2_v I__2424 (
            .O(N__21604),
            .I(N__21600));
    CascadeMux I__2423 (
            .O(N__21603),
            .I(N__21597));
    Sp12to4 I__2422 (
            .O(N__21600),
            .I(N__21594));
    InMux I__2421 (
            .O(N__21597),
            .I(N__21591));
    Odrv12 I__2420 (
            .O(N__21594),
            .I(DDS_SCK1));
    LocalMux I__2419 (
            .O(N__21591),
            .I(DDS_SCK1));
    CascadeMux I__2418 (
            .O(N__21586),
            .I(n23_adj_1512_cascade_));
    CascadeMux I__2417 (
            .O(N__21583),
            .I(N__21580));
    InMux I__2416 (
            .O(N__21580),
            .I(N__21576));
    InMux I__2415 (
            .O(N__21579),
            .I(N__21573));
    LocalMux I__2414 (
            .O(N__21576),
            .I(cmd_rdadctmp_6_adj_1437));
    LocalMux I__2413 (
            .O(N__21573),
            .I(cmd_rdadctmp_6_adj_1437));
    CascadeMux I__2412 (
            .O(N__21568),
            .I(N__21564));
    InMux I__2411 (
            .O(N__21567),
            .I(N__21561));
    InMux I__2410 (
            .O(N__21564),
            .I(N__21558));
    LocalMux I__2409 (
            .O(N__21561),
            .I(N__21554));
    LocalMux I__2408 (
            .O(N__21558),
            .I(N__21551));
    InMux I__2407 (
            .O(N__21557),
            .I(N__21548));
    Odrv12 I__2406 (
            .O(N__21554),
            .I(cmd_rdadctmp_21_adj_1422));
    Odrv4 I__2405 (
            .O(N__21551),
            .I(cmd_rdadctmp_21_adj_1422));
    LocalMux I__2404 (
            .O(N__21548),
            .I(cmd_rdadctmp_21_adj_1422));
    CascadeMux I__2403 (
            .O(N__21541),
            .I(N__21537));
    InMux I__2402 (
            .O(N__21540),
            .I(N__21534));
    InMux I__2401 (
            .O(N__21537),
            .I(N__21530));
    LocalMux I__2400 (
            .O(N__21534),
            .I(N__21527));
    InMux I__2399 (
            .O(N__21533),
            .I(N__21524));
    LocalMux I__2398 (
            .O(N__21530),
            .I(buf_adcdata_vac_13));
    Odrv4 I__2397 (
            .O(N__21527),
            .I(buf_adcdata_vac_13));
    LocalMux I__2396 (
            .O(N__21524),
            .I(buf_adcdata_vac_13));
    CascadeMux I__2395 (
            .O(N__21517),
            .I(N__21514));
    InMux I__2394 (
            .O(N__21514),
            .I(N__21510));
    InMux I__2393 (
            .O(N__21513),
            .I(N__21507));
    LocalMux I__2392 (
            .O(N__21510),
            .I(cmd_rdadctmp_4_adj_1439));
    LocalMux I__2391 (
            .O(N__21507),
            .I(cmd_rdadctmp_4_adj_1439));
    InMux I__2390 (
            .O(N__21502),
            .I(N__21496));
    InMux I__2389 (
            .O(N__21501),
            .I(N__21496));
    LocalMux I__2388 (
            .O(N__21496),
            .I(cmd_rdadctmp_5_adj_1438));
    InMux I__2387 (
            .O(N__21493),
            .I(N__21490));
    LocalMux I__2386 (
            .O(N__21490),
            .I(N__21487));
    Span4Mux_h I__2385 (
            .O(N__21487),
            .I(N__21484));
    Odrv4 I__2384 (
            .O(N__21484),
            .I(buf_data_iac_14));
    InMux I__2383 (
            .O(N__21481),
            .I(N__21478));
    LocalMux I__2382 (
            .O(N__21478),
            .I(N__21475));
    Span4Mux_h I__2381 (
            .O(N__21475),
            .I(N__21470));
    InMux I__2380 (
            .O(N__21474),
            .I(N__21467));
    InMux I__2379 (
            .O(N__21473),
            .I(N__21464));
    Span4Mux_v I__2378 (
            .O(N__21470),
            .I(N__21461));
    LocalMux I__2377 (
            .O(N__21467),
            .I(N__21458));
    LocalMux I__2376 (
            .O(N__21464),
            .I(buf_adcdata_vac_3));
    Odrv4 I__2375 (
            .O(N__21461),
            .I(buf_adcdata_vac_3));
    Odrv4 I__2374 (
            .O(N__21458),
            .I(buf_adcdata_vac_3));
    CascadeMux I__2373 (
            .O(N__21451),
            .I(N__21448));
    InMux I__2372 (
            .O(N__21448),
            .I(N__21443));
    CascadeMux I__2371 (
            .O(N__21447),
            .I(N__21440));
    CascadeMux I__2370 (
            .O(N__21446),
            .I(N__21437));
    LocalMux I__2369 (
            .O(N__21443),
            .I(N__21434));
    InMux I__2368 (
            .O(N__21440),
            .I(N__21431));
    InMux I__2367 (
            .O(N__21437),
            .I(N__21428));
    Odrv4 I__2366 (
            .O(N__21434),
            .I(cmd_rdadctmp_8));
    LocalMux I__2365 (
            .O(N__21431),
            .I(cmd_rdadctmp_8));
    LocalMux I__2364 (
            .O(N__21428),
            .I(cmd_rdadctmp_8));
    CascadeMux I__2363 (
            .O(N__21421),
            .I(N__21417));
    CascadeMux I__2362 (
            .O(N__21420),
            .I(N__21414));
    InMux I__2361 (
            .O(N__21417),
            .I(N__21406));
    InMux I__2360 (
            .O(N__21414),
            .I(N__21406));
    InMux I__2359 (
            .O(N__21413),
            .I(N__21406));
    LocalMux I__2358 (
            .O(N__21406),
            .I(cmd_rdadctmp_22_adj_1421));
    InMux I__2357 (
            .O(N__21403),
            .I(N__21400));
    LocalMux I__2356 (
            .O(N__21400),
            .I(n19_adj_1487));
    InMux I__2355 (
            .O(N__21397),
            .I(N__21394));
    LocalMux I__2354 (
            .O(N__21394),
            .I(N__21391));
    Span4Mux_h I__2353 (
            .O(N__21391),
            .I(N__21388));
    Span4Mux_v I__2352 (
            .O(N__21388),
            .I(N__21383));
    InMux I__2351 (
            .O(N__21387),
            .I(N__21378));
    InMux I__2350 (
            .O(N__21386),
            .I(N__21378));
    Odrv4 I__2349 (
            .O(N__21383),
            .I(buf_adcdata_vac_8));
    LocalMux I__2348 (
            .O(N__21378),
            .I(buf_adcdata_vac_8));
    InMux I__2347 (
            .O(N__21373),
            .I(N__21370));
    LocalMux I__2346 (
            .O(N__21370),
            .I(N__21367));
    Span4Mux_v I__2345 (
            .O(N__21367),
            .I(N__21363));
    CascadeMux I__2344 (
            .O(N__21366),
            .I(N__21360));
    Span4Mux_h I__2343 (
            .O(N__21363),
            .I(N__21357));
    InMux I__2342 (
            .O(N__21360),
            .I(N__21354));
    Odrv4 I__2341 (
            .O(N__21357),
            .I(buf_readRTD_0));
    LocalMux I__2340 (
            .O(N__21354),
            .I(buf_readRTD_0));
    CascadeMux I__2339 (
            .O(N__21349),
            .I(n19_adj_1479_cascade_));
    CascadeMux I__2338 (
            .O(N__21346),
            .I(N__21342));
    CascadeMux I__2337 (
            .O(N__21345),
            .I(N__21339));
    InMux I__2336 (
            .O(N__21342),
            .I(N__21335));
    InMux I__2335 (
            .O(N__21339),
            .I(N__21332));
    InMux I__2334 (
            .O(N__21338),
            .I(N__21329));
    LocalMux I__2333 (
            .O(N__21335),
            .I(cmd_rdadctmp_29_adj_1414));
    LocalMux I__2332 (
            .O(N__21332),
            .I(cmd_rdadctmp_29_adj_1414));
    LocalMux I__2331 (
            .O(N__21329),
            .I(cmd_rdadctmp_29_adj_1414));
    CascadeMux I__2330 (
            .O(N__21322),
            .I(N__21318));
    CascadeMux I__2329 (
            .O(N__21321),
            .I(N__21315));
    InMux I__2328 (
            .O(N__21318),
            .I(N__21311));
    InMux I__2327 (
            .O(N__21315),
            .I(N__21308));
    InMux I__2326 (
            .O(N__21314),
            .I(N__21305));
    LocalMux I__2325 (
            .O(N__21311),
            .I(cmd_rdadctmp_10));
    LocalMux I__2324 (
            .O(N__21308),
            .I(cmd_rdadctmp_10));
    LocalMux I__2323 (
            .O(N__21305),
            .I(cmd_rdadctmp_10));
    CascadeMux I__2322 (
            .O(N__21298),
            .I(N__21294));
    CascadeMux I__2321 (
            .O(N__21297),
            .I(N__21291));
    InMux I__2320 (
            .O(N__21294),
            .I(N__21287));
    InMux I__2319 (
            .O(N__21291),
            .I(N__21282));
    InMux I__2318 (
            .O(N__21290),
            .I(N__21282));
    LocalMux I__2317 (
            .O(N__21287),
            .I(cmd_rdadctmp_26_adj_1417));
    LocalMux I__2316 (
            .O(N__21282),
            .I(cmd_rdadctmp_26_adj_1417));
    CascadeMux I__2315 (
            .O(N__21277),
            .I(N__21273));
    CascadeMux I__2314 (
            .O(N__21276),
            .I(N__21270));
    InMux I__2313 (
            .O(N__21273),
            .I(N__21266));
    InMux I__2312 (
            .O(N__21270),
            .I(N__21263));
    InMux I__2311 (
            .O(N__21269),
            .I(N__21260));
    LocalMux I__2310 (
            .O(N__21266),
            .I(cmd_rdadctmp_27_adj_1416));
    LocalMux I__2309 (
            .O(N__21263),
            .I(cmd_rdadctmp_27_adj_1416));
    LocalMux I__2308 (
            .O(N__21260),
            .I(cmd_rdadctmp_27_adj_1416));
    InMux I__2307 (
            .O(N__21253),
            .I(N__21246));
    InMux I__2306 (
            .O(N__21252),
            .I(N__21246));
    InMux I__2305 (
            .O(N__21251),
            .I(N__21243));
    LocalMux I__2304 (
            .O(N__21246),
            .I(cmd_rdadctmp_9));
    LocalMux I__2303 (
            .O(N__21243),
            .I(cmd_rdadctmp_9));
    InMux I__2302 (
            .O(N__21238),
            .I(N__21234));
    CascadeMux I__2301 (
            .O(N__21237),
            .I(N__21231));
    LocalMux I__2300 (
            .O(N__21234),
            .I(N__21227));
    InMux I__2299 (
            .O(N__21231),
            .I(N__21224));
    InMux I__2298 (
            .O(N__21230),
            .I(N__21221));
    Odrv4 I__2297 (
            .O(N__21227),
            .I(cmd_rdadctmp_23_adj_1420));
    LocalMux I__2296 (
            .O(N__21224),
            .I(cmd_rdadctmp_23_adj_1420));
    LocalMux I__2295 (
            .O(N__21221),
            .I(cmd_rdadctmp_23_adj_1420));
    InMux I__2294 (
            .O(N__21214),
            .I(N__21210));
    InMux I__2293 (
            .O(N__21213),
            .I(N__21207));
    LocalMux I__2292 (
            .O(N__21210),
            .I(\RTD.cfg_buf_5 ));
    LocalMux I__2291 (
            .O(N__21207),
            .I(\RTD.cfg_buf_5 ));
    InMux I__2290 (
            .O(N__21202),
            .I(N__21199));
    LocalMux I__2289 (
            .O(N__21199),
            .I(\RTD.n11_adj_1396 ));
    InMux I__2288 (
            .O(N__21196),
            .I(N__21190));
    InMux I__2287 (
            .O(N__21195),
            .I(N__21190));
    LocalMux I__2286 (
            .O(N__21190),
            .I(\RTD.cfg_buf_3 ));
    InMux I__2285 (
            .O(N__21187),
            .I(N__21170));
    InMux I__2284 (
            .O(N__21186),
            .I(N__21170));
    InMux I__2283 (
            .O(N__21185),
            .I(N__21170));
    InMux I__2282 (
            .O(N__21184),
            .I(N__21170));
    InMux I__2281 (
            .O(N__21183),
            .I(N__21170));
    InMux I__2280 (
            .O(N__21182),
            .I(N__21165));
    InMux I__2279 (
            .O(N__21181),
            .I(N__21165));
    LocalMux I__2278 (
            .O(N__21170),
            .I(n18586));
    LocalMux I__2277 (
            .O(N__21165),
            .I(n18586));
    InMux I__2276 (
            .O(N__21160),
            .I(N__21149));
    InMux I__2275 (
            .O(N__21159),
            .I(N__21146));
    InMux I__2274 (
            .O(N__21158),
            .I(N__21141));
    InMux I__2273 (
            .O(N__21157),
            .I(N__21141));
    InMux I__2272 (
            .O(N__21156),
            .I(N__21134));
    InMux I__2271 (
            .O(N__21155),
            .I(N__21134));
    InMux I__2270 (
            .O(N__21154),
            .I(N__21134));
    InMux I__2269 (
            .O(N__21153),
            .I(N__21131));
    InMux I__2268 (
            .O(N__21152),
            .I(N__21128));
    LocalMux I__2267 (
            .O(N__21149),
            .I(n13162));
    LocalMux I__2266 (
            .O(N__21146),
            .I(n13162));
    LocalMux I__2265 (
            .O(N__21141),
            .I(n13162));
    LocalMux I__2264 (
            .O(N__21134),
            .I(n13162));
    LocalMux I__2263 (
            .O(N__21131),
            .I(n13162));
    LocalMux I__2262 (
            .O(N__21128),
            .I(n13162));
    InMux I__2261 (
            .O(N__21115),
            .I(N__21111));
    InMux I__2260 (
            .O(N__21114),
            .I(N__21108));
    LocalMux I__2259 (
            .O(N__21111),
            .I(\RTD.cfg_buf_6 ));
    LocalMux I__2258 (
            .O(N__21108),
            .I(\RTD.cfg_buf_6 ));
    CascadeMux I__2257 (
            .O(N__21103),
            .I(N__21100));
    InMux I__2256 (
            .O(N__21100),
            .I(N__21097));
    LocalMux I__2255 (
            .O(N__21097),
            .I(N__21093));
    CascadeMux I__2254 (
            .O(N__21096),
            .I(N__21090));
    Span4Mux_h I__2253 (
            .O(N__21093),
            .I(N__21087));
    InMux I__2252 (
            .O(N__21090),
            .I(N__21084));
    Odrv4 I__2251 (
            .O(N__21087),
            .I(buf_readRTD_11));
    LocalMux I__2250 (
            .O(N__21084),
            .I(buf_readRTD_11));
    CascadeMux I__2249 (
            .O(N__21079),
            .I(n22099_cascade_));
    CascadeMux I__2248 (
            .O(N__21076),
            .I(n22102_cascade_));
    InMux I__2247 (
            .O(N__21073),
            .I(N__21070));
    LocalMux I__2246 (
            .O(N__21070),
            .I(N__21066));
    InMux I__2245 (
            .O(N__21069),
            .I(N__21062));
    Span4Mux_h I__2244 (
            .O(N__21066),
            .I(N__21059));
    InMux I__2243 (
            .O(N__21065),
            .I(N__21056));
    LocalMux I__2242 (
            .O(N__21062),
            .I(buf_adcdata_vac_19));
    Odrv4 I__2241 (
            .O(N__21059),
            .I(buf_adcdata_vac_19));
    LocalMux I__2240 (
            .O(N__21056),
            .I(buf_adcdata_vac_19));
    CascadeMux I__2239 (
            .O(N__21049),
            .I(n19_adj_1610_cascade_));
    InMux I__2238 (
            .O(N__21046),
            .I(N__21043));
    LocalMux I__2237 (
            .O(N__21043),
            .I(N__21039));
    InMux I__2236 (
            .O(N__21042),
            .I(N__21035));
    Span4Mux_v I__2235 (
            .O(N__21039),
            .I(N__21032));
    InMux I__2234 (
            .O(N__21038),
            .I(N__21029));
    LocalMux I__2233 (
            .O(N__21035),
            .I(buf_adcdata_iac_3));
    Odrv4 I__2232 (
            .O(N__21032),
            .I(buf_adcdata_iac_3));
    LocalMux I__2231 (
            .O(N__21029),
            .I(buf_adcdata_iac_3));
    InMux I__2230 (
            .O(N__21022),
            .I(N__21019));
    LocalMux I__2229 (
            .O(N__21019),
            .I(n22_adj_1611));
    InMux I__2228 (
            .O(N__21016),
            .I(N__21013));
    LocalMux I__2227 (
            .O(N__21013),
            .I(\RTD.cfg_tmp_5 ));
    InMux I__2226 (
            .O(N__21010),
            .I(N__21007));
    LocalMux I__2225 (
            .O(N__21007),
            .I(\RTD.cfg_tmp_6 ));
    CascadeMux I__2224 (
            .O(N__21004),
            .I(N__21001));
    InMux I__2223 (
            .O(N__21001),
            .I(N__20998));
    LocalMux I__2222 (
            .O(N__20998),
            .I(N__20995));
    Span4Mux_h I__2221 (
            .O(N__20995),
            .I(N__20991));
    InMux I__2220 (
            .O(N__20994),
            .I(N__20988));
    Odrv4 I__2219 (
            .O(N__20991),
            .I(\RTD.cfg_tmp_7 ));
    LocalMux I__2218 (
            .O(N__20988),
            .I(\RTD.cfg_tmp_7 ));
    InMux I__2217 (
            .O(N__20983),
            .I(N__20980));
    LocalMux I__2216 (
            .O(N__20980),
            .I(\RTD.cfg_tmp_0 ));
    CascadeMux I__2215 (
            .O(N__20977),
            .I(N__20974));
    InMux I__2214 (
            .O(N__20974),
            .I(N__20971));
    LocalMux I__2213 (
            .O(N__20971),
            .I(N__20960));
    InMux I__2212 (
            .O(N__20970),
            .I(N__20949));
    InMux I__2211 (
            .O(N__20969),
            .I(N__20949));
    InMux I__2210 (
            .O(N__20968),
            .I(N__20949));
    InMux I__2209 (
            .O(N__20967),
            .I(N__20949));
    InMux I__2208 (
            .O(N__20966),
            .I(N__20949));
    InMux I__2207 (
            .O(N__20965),
            .I(N__20946));
    InMux I__2206 (
            .O(N__20964),
            .I(N__20929));
    InMux I__2205 (
            .O(N__20963),
            .I(N__20920));
    Span4Mux_v I__2204 (
            .O(N__20960),
            .I(N__20915));
    LocalMux I__2203 (
            .O(N__20949),
            .I(N__20915));
    LocalMux I__2202 (
            .O(N__20946),
            .I(N__20910));
    InMux I__2201 (
            .O(N__20945),
            .I(N__20907));
    InMux I__2200 (
            .O(N__20944),
            .I(N__20898));
    InMux I__2199 (
            .O(N__20943),
            .I(N__20898));
    InMux I__2198 (
            .O(N__20942),
            .I(N__20898));
    InMux I__2197 (
            .O(N__20941),
            .I(N__20898));
    InMux I__2196 (
            .O(N__20940),
            .I(N__20890));
    InMux I__2195 (
            .O(N__20939),
            .I(N__20873));
    InMux I__2194 (
            .O(N__20938),
            .I(N__20873));
    InMux I__2193 (
            .O(N__20937),
            .I(N__20873));
    InMux I__2192 (
            .O(N__20936),
            .I(N__20873));
    InMux I__2191 (
            .O(N__20935),
            .I(N__20873));
    InMux I__2190 (
            .O(N__20934),
            .I(N__20873));
    InMux I__2189 (
            .O(N__20933),
            .I(N__20873));
    InMux I__2188 (
            .O(N__20932),
            .I(N__20873));
    LocalMux I__2187 (
            .O(N__20929),
            .I(N__20870));
    InMux I__2186 (
            .O(N__20928),
            .I(N__20867));
    InMux I__2185 (
            .O(N__20927),
            .I(N__20856));
    InMux I__2184 (
            .O(N__20926),
            .I(N__20856));
    InMux I__2183 (
            .O(N__20925),
            .I(N__20856));
    InMux I__2182 (
            .O(N__20924),
            .I(N__20856));
    InMux I__2181 (
            .O(N__20923),
            .I(N__20856));
    LocalMux I__2180 (
            .O(N__20920),
            .I(N__20851));
    Span4Mux_v I__2179 (
            .O(N__20915),
            .I(N__20851));
    InMux I__2178 (
            .O(N__20914),
            .I(N__20846));
    InMux I__2177 (
            .O(N__20913),
            .I(N__20846));
    Span4Mux_h I__2176 (
            .O(N__20910),
            .I(N__20839));
    LocalMux I__2175 (
            .O(N__20907),
            .I(N__20839));
    LocalMux I__2174 (
            .O(N__20898),
            .I(N__20839));
    InMux I__2173 (
            .O(N__20897),
            .I(N__20828));
    InMux I__2172 (
            .O(N__20896),
            .I(N__20828));
    InMux I__2171 (
            .O(N__20895),
            .I(N__20828));
    InMux I__2170 (
            .O(N__20894),
            .I(N__20828));
    InMux I__2169 (
            .O(N__20893),
            .I(N__20828));
    LocalMux I__2168 (
            .O(N__20890),
            .I(\RTD.adc_state_0 ));
    LocalMux I__2167 (
            .O(N__20873),
            .I(\RTD.adc_state_0 ));
    Odrv12 I__2166 (
            .O(N__20870),
            .I(\RTD.adc_state_0 ));
    LocalMux I__2165 (
            .O(N__20867),
            .I(\RTD.adc_state_0 ));
    LocalMux I__2164 (
            .O(N__20856),
            .I(\RTD.adc_state_0 ));
    Odrv4 I__2163 (
            .O(N__20851),
            .I(\RTD.adc_state_0 ));
    LocalMux I__2162 (
            .O(N__20846),
            .I(\RTD.adc_state_0 ));
    Odrv4 I__2161 (
            .O(N__20839),
            .I(\RTD.adc_state_0 ));
    LocalMux I__2160 (
            .O(N__20828),
            .I(\RTD.adc_state_0 ));
    CascadeMux I__2159 (
            .O(N__20809),
            .I(n18586_cascade_));
    InMux I__2158 (
            .O(N__20806),
            .I(N__20800));
    InMux I__2157 (
            .O(N__20805),
            .I(N__20800));
    LocalMux I__2156 (
            .O(N__20800),
            .I(cfg_buf_0));
    InMux I__2155 (
            .O(N__20797),
            .I(N__20794));
    LocalMux I__2154 (
            .O(N__20794),
            .I(\RTD.n9 ));
    InMux I__2153 (
            .O(N__20791),
            .I(N__20787));
    InMux I__2152 (
            .O(N__20790),
            .I(N__20784));
    LocalMux I__2151 (
            .O(N__20787),
            .I(\RTD.n11 ));
    LocalMux I__2150 (
            .O(N__20784),
            .I(\RTD.n11 ));
    InMux I__2149 (
            .O(N__20779),
            .I(N__20776));
    LocalMux I__2148 (
            .O(N__20776),
            .I(N__20773));
    Odrv4 I__2147 (
            .O(N__20773),
            .I(\RTD.n14 ));
    CascadeMux I__2146 (
            .O(N__20770),
            .I(\RTD.n20722_cascade_ ));
    CEMux I__2145 (
            .O(N__20767),
            .I(N__20764));
    LocalMux I__2144 (
            .O(N__20764),
            .I(N__20761));
    Span4Mux_h I__2143 (
            .O(N__20761),
            .I(N__20758));
    Odrv4 I__2142 (
            .O(N__20758),
            .I(\RTD.n13198 ));
    CascadeMux I__2141 (
            .O(N__20755),
            .I(\RTD.n13198_cascade_ ));
    SRMux I__2140 (
            .O(N__20752),
            .I(N__20749));
    LocalMux I__2139 (
            .O(N__20749),
            .I(N__20746));
    Span4Mux_h I__2138 (
            .O(N__20746),
            .I(N__20743));
    Odrv4 I__2137 (
            .O(N__20743),
            .I(\RTD.n14984 ));
    SRMux I__2136 (
            .O(N__20740),
            .I(N__20737));
    LocalMux I__2135 (
            .O(N__20737),
            .I(N__20734));
    Odrv4 I__2134 (
            .O(N__20734),
            .I(\CLK_DDS.n16711 ));
    InMux I__2133 (
            .O(N__20731),
            .I(N__20727));
    InMux I__2132 (
            .O(N__20730),
            .I(N__20724));
    LocalMux I__2131 (
            .O(N__20727),
            .I(\RTD.n7285 ));
    LocalMux I__2130 (
            .O(N__20724),
            .I(\RTD.n7285 ));
    CascadeMux I__2129 (
            .O(N__20719),
            .I(N__20716));
    InMux I__2128 (
            .O(N__20716),
            .I(N__20713));
    LocalMux I__2127 (
            .O(N__20713),
            .I(\RTD.n11_adj_1394 ));
    InMux I__2126 (
            .O(N__20710),
            .I(N__20707));
    LocalMux I__2125 (
            .O(N__20707),
            .I(\RTD.n21091 ));
    CascadeMux I__2124 (
            .O(N__20704),
            .I(N__20701));
    InMux I__2123 (
            .O(N__20701),
            .I(N__20698));
    LocalMux I__2122 (
            .O(N__20698),
            .I(\RTD.n33 ));
    InMux I__2121 (
            .O(N__20695),
            .I(N__20692));
    LocalMux I__2120 (
            .O(N__20692),
            .I(\RTD.n17676 ));
    InMux I__2119 (
            .O(N__20689),
            .I(N__20686));
    LocalMux I__2118 (
            .O(N__20686),
            .I(\RTD.n7_adj_1395 ));
    CEMux I__2117 (
            .O(N__20683),
            .I(N__20680));
    LocalMux I__2116 (
            .O(N__20680),
            .I(N__20676));
    CEMux I__2115 (
            .O(N__20679),
            .I(N__20673));
    Odrv12 I__2114 (
            .O(N__20676),
            .I(\RTD.n11712 ));
    LocalMux I__2113 (
            .O(N__20673),
            .I(\RTD.n11712 ));
    CascadeMux I__2112 (
            .O(N__20668),
            .I(N__20665));
    InMux I__2111 (
            .O(N__20665),
            .I(N__20662));
    LocalMux I__2110 (
            .O(N__20662),
            .I(\RTD.cfg_tmp_1 ));
    InMux I__2109 (
            .O(N__20659),
            .I(N__20656));
    LocalMux I__2108 (
            .O(N__20656),
            .I(\RTD.cfg_tmp_2 ));
    InMux I__2107 (
            .O(N__20653),
            .I(N__20650));
    LocalMux I__2106 (
            .O(N__20650),
            .I(\RTD.cfg_tmp_3 ));
    InMux I__2105 (
            .O(N__20647),
            .I(N__20644));
    LocalMux I__2104 (
            .O(N__20644),
            .I(\RTD.cfg_tmp_4 ));
    CEMux I__2103 (
            .O(N__20641),
            .I(N__20637));
    CEMux I__2102 (
            .O(N__20640),
            .I(N__20634));
    LocalMux I__2101 (
            .O(N__20637),
            .I(N__20631));
    LocalMux I__2100 (
            .O(N__20634),
            .I(N__20628));
    Span4Mux_h I__2099 (
            .O(N__20631),
            .I(N__20625));
    Odrv12 I__2098 (
            .O(N__20628),
            .I(\CLK_DDS.n9 ));
    Odrv4 I__2097 (
            .O(N__20625),
            .I(\CLK_DDS.n9 ));
    InMux I__2096 (
            .O(N__20620),
            .I(N__20617));
    LocalMux I__2095 (
            .O(N__20617),
            .I(N__20611));
    InMux I__2094 (
            .O(N__20616),
            .I(N__20606));
    InMux I__2093 (
            .O(N__20615),
            .I(N__20606));
    InMux I__2092 (
            .O(N__20614),
            .I(N__20603));
    Odrv4 I__2091 (
            .O(N__20611),
            .I(\RTD.bit_cnt_1 ));
    LocalMux I__2090 (
            .O(N__20606),
            .I(\RTD.bit_cnt_1 ));
    LocalMux I__2089 (
            .O(N__20603),
            .I(\RTD.bit_cnt_1 ));
    InMux I__2088 (
            .O(N__20596),
            .I(N__20592));
    CascadeMux I__2087 (
            .O(N__20595),
            .I(N__20589));
    LocalMux I__2086 (
            .O(N__20592),
            .I(N__20583));
    InMux I__2085 (
            .O(N__20589),
            .I(N__20576));
    InMux I__2084 (
            .O(N__20588),
            .I(N__20576));
    InMux I__2083 (
            .O(N__20587),
            .I(N__20576));
    InMux I__2082 (
            .O(N__20586),
            .I(N__20573));
    Odrv4 I__2081 (
            .O(N__20583),
            .I(\RTD.bit_cnt_0 ));
    LocalMux I__2080 (
            .O(N__20576),
            .I(\RTD.bit_cnt_0 ));
    LocalMux I__2079 (
            .O(N__20573),
            .I(\RTD.bit_cnt_0 ));
    InMux I__2078 (
            .O(N__20566),
            .I(N__20563));
    LocalMux I__2077 (
            .O(N__20563),
            .I(N__20558));
    InMux I__2076 (
            .O(N__20562),
            .I(N__20555));
    InMux I__2075 (
            .O(N__20561),
            .I(N__20552));
    Odrv4 I__2074 (
            .O(N__20558),
            .I(\RTD.bit_cnt_2 ));
    LocalMux I__2073 (
            .O(N__20555),
            .I(\RTD.bit_cnt_2 ));
    LocalMux I__2072 (
            .O(N__20552),
            .I(\RTD.bit_cnt_2 ));
    InMux I__2071 (
            .O(N__20545),
            .I(N__20541));
    InMux I__2070 (
            .O(N__20544),
            .I(N__20537));
    LocalMux I__2069 (
            .O(N__20541),
            .I(N__20534));
    InMux I__2068 (
            .O(N__20540),
            .I(N__20531));
    LocalMux I__2067 (
            .O(N__20537),
            .I(\RTD.n17638 ));
    Odrv4 I__2066 (
            .O(N__20534),
            .I(\RTD.n17638 ));
    LocalMux I__2065 (
            .O(N__20531),
            .I(\RTD.n17638 ));
    CascadeMux I__2064 (
            .O(N__20524),
            .I(N__20521));
    InMux I__2063 (
            .O(N__20521),
            .I(N__20514));
    InMux I__2062 (
            .O(N__20520),
            .I(N__20511));
    InMux I__2061 (
            .O(N__20519),
            .I(N__20508));
    InMux I__2060 (
            .O(N__20518),
            .I(N__20505));
    CascadeMux I__2059 (
            .O(N__20517),
            .I(N__20502));
    LocalMux I__2058 (
            .O(N__20514),
            .I(N__20493));
    LocalMux I__2057 (
            .O(N__20511),
            .I(N__20493));
    LocalMux I__2056 (
            .O(N__20508),
            .I(N__20493));
    LocalMux I__2055 (
            .O(N__20505),
            .I(N__20493));
    InMux I__2054 (
            .O(N__20502),
            .I(N__20490));
    Span4Mux_v I__2053 (
            .O(N__20493),
            .I(N__20487));
    LocalMux I__2052 (
            .O(N__20490),
            .I(\RTD.bit_cnt_3 ));
    Odrv4 I__2051 (
            .O(N__20487),
            .I(\RTD.bit_cnt_3 ));
    CascadeMux I__2050 (
            .O(N__20482),
            .I(\RTD.n17638_cascade_ ));
    InMux I__2049 (
            .O(N__20479),
            .I(N__20476));
    LocalMux I__2048 (
            .O(N__20476),
            .I(N__20472));
    InMux I__2047 (
            .O(N__20475),
            .I(N__20469));
    Span4Mux_h I__2046 (
            .O(N__20472),
            .I(N__20466));
    LocalMux I__2045 (
            .O(N__20469),
            .I(\RTD.n1_adj_1392 ));
    Odrv4 I__2044 (
            .O(N__20466),
            .I(\RTD.n1_adj_1392 ));
    CascadeMux I__2043 (
            .O(N__20461),
            .I(\RTD.n21063_cascade_ ));
    CascadeMux I__2042 (
            .O(N__20458),
            .I(N__20454));
    CascadeMux I__2041 (
            .O(N__20457),
            .I(N__20450));
    InMux I__2040 (
            .O(N__20454),
            .I(N__20446));
    InMux I__2039 (
            .O(N__20453),
            .I(N__20439));
    InMux I__2038 (
            .O(N__20450),
            .I(N__20439));
    InMux I__2037 (
            .O(N__20449),
            .I(N__20439));
    LocalMux I__2036 (
            .O(N__20446),
            .I(N__20436));
    LocalMux I__2035 (
            .O(N__20439),
            .I(bit_cnt_1));
    Odrv4 I__2034 (
            .O(N__20436),
            .I(bit_cnt_1));
    InMux I__2033 (
            .O(N__20431),
            .I(N__20426));
    InMux I__2032 (
            .O(N__20430),
            .I(N__20421));
    InMux I__2031 (
            .O(N__20429),
            .I(N__20421));
    LocalMux I__2030 (
            .O(N__20426),
            .I(N__20418));
    LocalMux I__2029 (
            .O(N__20421),
            .I(bit_cnt_2));
    Odrv4 I__2028 (
            .O(N__20418),
            .I(bit_cnt_2));
    InMux I__2027 (
            .O(N__20413),
            .I(N__20410));
    LocalMux I__2026 (
            .O(N__20410),
            .I(n8_adj_1409));
    InMux I__2025 (
            .O(N__20407),
            .I(N__20404));
    LocalMux I__2024 (
            .O(N__20404),
            .I(N__20401));
    Odrv4 I__2023 (
            .O(N__20401),
            .I(buf_data_iac_8));
    CascadeMux I__2022 (
            .O(N__20398),
            .I(N__20395));
    CascadeBuf I__2021 (
            .O(N__20395),
            .I(N__20392));
    CascadeMux I__2020 (
            .O(N__20392),
            .I(N__20389));
    CascadeBuf I__2019 (
            .O(N__20389),
            .I(N__20386));
    CascadeMux I__2018 (
            .O(N__20386),
            .I(N__20383));
    CascadeBuf I__2017 (
            .O(N__20383),
            .I(N__20380));
    CascadeMux I__2016 (
            .O(N__20380),
            .I(N__20377));
    CascadeBuf I__2015 (
            .O(N__20377),
            .I(N__20374));
    CascadeMux I__2014 (
            .O(N__20374),
            .I(N__20371));
    CascadeBuf I__2013 (
            .O(N__20371),
            .I(N__20368));
    CascadeMux I__2012 (
            .O(N__20368),
            .I(N__20364));
    CascadeMux I__2011 (
            .O(N__20367),
            .I(N__20361));
    CascadeBuf I__2010 (
            .O(N__20364),
            .I(N__20358));
    CascadeBuf I__2009 (
            .O(N__20361),
            .I(N__20355));
    CascadeMux I__2008 (
            .O(N__20358),
            .I(N__20352));
    CascadeMux I__2007 (
            .O(N__20355),
            .I(N__20349));
    CascadeBuf I__2006 (
            .O(N__20352),
            .I(N__20346));
    InMux I__2005 (
            .O(N__20349),
            .I(N__20343));
    CascadeMux I__2004 (
            .O(N__20346),
            .I(N__20340));
    LocalMux I__2003 (
            .O(N__20343),
            .I(N__20337));
    CascadeBuf I__2002 (
            .O(N__20340),
            .I(N__20334));
    Span4Mux_v I__2001 (
            .O(N__20337),
            .I(N__20331));
    CascadeMux I__2000 (
            .O(N__20334),
            .I(N__20328));
    Span4Mux_v I__1999 (
            .O(N__20331),
            .I(N__20325));
    CascadeBuf I__1998 (
            .O(N__20328),
            .I(N__20322));
    Span4Mux_h I__1997 (
            .O(N__20325),
            .I(N__20319));
    CascadeMux I__1996 (
            .O(N__20322),
            .I(N__20316));
    Sp12to4 I__1995 (
            .O(N__20319),
            .I(N__20313));
    InMux I__1994 (
            .O(N__20316),
            .I(N__20310));
    Odrv12 I__1993 (
            .O(N__20313),
            .I(data_index_9_N_212_7));
    LocalMux I__1992 (
            .O(N__20310),
            .I(data_index_9_N_212_7));
    CascadeMux I__1991 (
            .O(N__20305),
            .I(N__20301));
    InMux I__1990 (
            .O(N__20304),
            .I(N__20293));
    InMux I__1989 (
            .O(N__20301),
            .I(N__20293));
    InMux I__1988 (
            .O(N__20300),
            .I(N__20293));
    LocalMux I__1987 (
            .O(N__20293),
            .I(cmd_rdadctmp_28_adj_1415));
    CascadeMux I__1986 (
            .O(N__20290),
            .I(N__20287));
    InMux I__1985 (
            .O(N__20287),
            .I(N__20284));
    LocalMux I__1984 (
            .O(N__20284),
            .I(N__20281));
    Span4Mux_v I__1983 (
            .O(N__20281),
            .I(N__20277));
    CascadeMux I__1982 (
            .O(N__20280),
            .I(N__20274));
    Span4Mux_v I__1981 (
            .O(N__20277),
            .I(N__20271));
    InMux I__1980 (
            .O(N__20274),
            .I(N__20268));
    Odrv4 I__1979 (
            .O(N__20271),
            .I(buf_readRTD_5));
    LocalMux I__1978 (
            .O(N__20268),
            .I(buf_readRTD_5));
    InMux I__1977 (
            .O(N__20263),
            .I(N__20260));
    LocalMux I__1976 (
            .O(N__20260),
            .I(n14_adj_1577));
    CascadeMux I__1975 (
            .O(N__20257),
            .I(n20573_cascade_));
    IoInMux I__1974 (
            .O(N__20254),
            .I(N__20251));
    LocalMux I__1973 (
            .O(N__20251),
            .I(N__20248));
    Span4Mux_s2_h I__1972 (
            .O(N__20248),
            .I(N__20245));
    Span4Mux_h I__1971 (
            .O(N__20245),
            .I(N__20241));
    CascadeMux I__1970 (
            .O(N__20244),
            .I(N__20238));
    Span4Mux_v I__1969 (
            .O(N__20241),
            .I(N__20235));
    InMux I__1968 (
            .O(N__20238),
            .I(N__20232));
    Odrv4 I__1967 (
            .O(N__20235),
            .I(VAC_CS));
    LocalMux I__1966 (
            .O(N__20232),
            .I(VAC_CS));
    IoInMux I__1965 (
            .O(N__20227),
            .I(N__20224));
    LocalMux I__1964 (
            .O(N__20224),
            .I(N__20221));
    IoSpan4Mux I__1963 (
            .O(N__20221),
            .I(N__20218));
    Span4Mux_s2_h I__1962 (
            .O(N__20218),
            .I(N__20214));
    CascadeMux I__1961 (
            .O(N__20217),
            .I(N__20211));
    Span4Mux_h I__1960 (
            .O(N__20214),
            .I(N__20208));
    InMux I__1959 (
            .O(N__20211),
            .I(N__20205));
    Odrv4 I__1958 (
            .O(N__20208),
            .I(VAC_SCLK));
    LocalMux I__1957 (
            .O(N__20205),
            .I(VAC_SCLK));
    CascadeMux I__1956 (
            .O(N__20200),
            .I(n19_adj_1622_cascade_));
    InMux I__1955 (
            .O(N__20197),
            .I(N__20194));
    LocalMux I__1954 (
            .O(N__20194),
            .I(N__20191));
    Span4Mux_v I__1953 (
            .O(N__20191),
            .I(N__20186));
    InMux I__1952 (
            .O(N__20190),
            .I(N__20181));
    InMux I__1951 (
            .O(N__20189),
            .I(N__20181));
    Odrv4 I__1950 (
            .O(N__20186),
            .I(buf_adcdata_vac_15));
    LocalMux I__1949 (
            .O(N__20181),
            .I(buf_adcdata_vac_15));
    InMux I__1948 (
            .O(N__20176),
            .I(N__20173));
    LocalMux I__1947 (
            .O(N__20173),
            .I(N__20170));
    Span4Mux_v I__1946 (
            .O(N__20170),
            .I(N__20167));
    Odrv4 I__1945 (
            .O(N__20167),
            .I(buf_data_iac_3));
    InMux I__1944 (
            .O(N__20164),
            .I(N__20161));
    LocalMux I__1943 (
            .O(N__20161),
            .I(N__20158));
    Span4Mux_v I__1942 (
            .O(N__20158),
            .I(N__20155));
    Span4Mux_v I__1941 (
            .O(N__20155),
            .I(N__20152));
    Odrv4 I__1940 (
            .O(N__20152),
            .I(buf_data_iac_21));
    CascadeMux I__1939 (
            .O(N__20149),
            .I(N__20146));
    InMux I__1938 (
            .O(N__20146),
            .I(N__20139));
    InMux I__1937 (
            .O(N__20145),
            .I(N__20136));
    InMux I__1936 (
            .O(N__20144),
            .I(N__20133));
    InMux I__1935 (
            .O(N__20143),
            .I(N__20130));
    InMux I__1934 (
            .O(N__20142),
            .I(N__20127));
    LocalMux I__1933 (
            .O(N__20139),
            .I(N__20120));
    LocalMux I__1932 (
            .O(N__20136),
            .I(N__20120));
    LocalMux I__1931 (
            .O(N__20133),
            .I(N__20120));
    LocalMux I__1930 (
            .O(N__20130),
            .I(\RTD.adress_7_N_1331_7 ));
    LocalMux I__1929 (
            .O(N__20127),
            .I(\RTD.adress_7_N_1331_7 ));
    Odrv4 I__1928 (
            .O(N__20120),
            .I(\RTD.adress_7_N_1331_7 ));
    InMux I__1927 (
            .O(N__20113),
            .I(N__20110));
    LocalMux I__1926 (
            .O(N__20110),
            .I(N__20107));
    Odrv4 I__1925 (
            .O(N__20107),
            .I(\RTD.n16 ));
    CascadeMux I__1924 (
            .O(N__20104),
            .I(N__20099));
    InMux I__1923 (
            .O(N__20103),
            .I(N__20093));
    InMux I__1922 (
            .O(N__20102),
            .I(N__20093));
    InMux I__1921 (
            .O(N__20099),
            .I(N__20088));
    InMux I__1920 (
            .O(N__20098),
            .I(N__20088));
    LocalMux I__1919 (
            .O(N__20093),
            .I(N__20085));
    LocalMux I__1918 (
            .O(N__20088),
            .I(N__20082));
    Odrv12 I__1917 (
            .O(N__20085),
            .I(\RTD.mode ));
    Odrv4 I__1916 (
            .O(N__20082),
            .I(\RTD.mode ));
    InMux I__1915 (
            .O(N__20077),
            .I(N__20074));
    LocalMux I__1914 (
            .O(N__20074),
            .I(\RTD.n10 ));
    InMux I__1913 (
            .O(N__20071),
            .I(N__20065));
    InMux I__1912 (
            .O(N__20070),
            .I(N__20065));
    LocalMux I__1911 (
            .O(N__20065),
            .I(\RTD.cfg_buf_2 ));
    InMux I__1910 (
            .O(N__20062),
            .I(N__20056));
    InMux I__1909 (
            .O(N__20061),
            .I(N__20056));
    LocalMux I__1908 (
            .O(N__20056),
            .I(\RTD.cfg_buf_4 ));
    InMux I__1907 (
            .O(N__20053),
            .I(N__20047));
    InMux I__1906 (
            .O(N__20052),
            .I(N__20047));
    LocalMux I__1905 (
            .O(N__20047),
            .I(\RTD.cfg_buf_7 ));
    CascadeMux I__1904 (
            .O(N__20044),
            .I(N__20041));
    InMux I__1903 (
            .O(N__20041),
            .I(N__20038));
    LocalMux I__1902 (
            .O(N__20038),
            .I(\RTD.n12 ));
    InMux I__1901 (
            .O(N__20035),
            .I(N__20029));
    InMux I__1900 (
            .O(N__20034),
            .I(N__20029));
    LocalMux I__1899 (
            .O(N__20029),
            .I(cfg_buf_1));
    InMux I__1898 (
            .O(N__20026),
            .I(N__20023));
    LocalMux I__1897 (
            .O(N__20023),
            .I(N__20019));
    CascadeMux I__1896 (
            .O(N__20022),
            .I(N__20016));
    Span4Mux_v I__1895 (
            .O(N__20019),
            .I(N__20013));
    InMux I__1894 (
            .O(N__20016),
            .I(N__20010));
    Odrv4 I__1893 (
            .O(N__20013),
            .I(buf_readRTD_7));
    LocalMux I__1892 (
            .O(N__20010),
            .I(buf_readRTD_7));
    InMux I__1891 (
            .O(N__20005),
            .I(N__20002));
    LocalMux I__1890 (
            .O(N__20002),
            .I(\RTD.n32 ));
    InMux I__1889 (
            .O(N__19999),
            .I(N__19996));
    LocalMux I__1888 (
            .O(N__19996),
            .I(N__19993));
    Span4Mux_h I__1887 (
            .O(N__19993),
            .I(N__19989));
    InMux I__1886 (
            .O(N__19992),
            .I(N__19986));
    Odrv4 I__1885 (
            .O(N__19989),
            .I(adress_6));
    LocalMux I__1884 (
            .O(N__19986),
            .I(adress_6));
    InMux I__1883 (
            .O(N__19981),
            .I(N__19977));
    InMux I__1882 (
            .O(N__19980),
            .I(N__19974));
    LocalMux I__1881 (
            .O(N__19977),
            .I(N__19971));
    LocalMux I__1880 (
            .O(N__19974),
            .I(\RTD.adress_7 ));
    Odrv12 I__1879 (
            .O(N__19971),
            .I(\RTD.adress_7 ));
    InMux I__1878 (
            .O(N__19966),
            .I(N__19963));
    LocalMux I__1877 (
            .O(N__19963),
            .I(N__19960));
    Odrv12 I__1876 (
            .O(N__19960),
            .I(adress_0));
    SRMux I__1875 (
            .O(N__19957),
            .I(N__19954));
    LocalMux I__1874 (
            .O(N__19954),
            .I(N__19950));
    SRMux I__1873 (
            .O(N__19953),
            .I(N__19947));
    Span4Mux_v I__1872 (
            .O(N__19950),
            .I(N__19942));
    LocalMux I__1871 (
            .O(N__19947),
            .I(N__19942));
    Span4Mux_v I__1870 (
            .O(N__19942),
            .I(N__19939));
    Odrv4 I__1869 (
            .O(N__19939),
            .I(\RTD.n19855 ));
    CascadeMux I__1868 (
            .O(N__19936),
            .I(\RTD.adress_7_N_1331_7_cascade_ ));
    InMux I__1867 (
            .O(N__19933),
            .I(N__19930));
    LocalMux I__1866 (
            .O(N__19930),
            .I(N__19925));
    InMux I__1865 (
            .O(N__19929),
            .I(N__19922));
    InMux I__1864 (
            .O(N__19928),
            .I(N__19919));
    Span4Mux_v I__1863 (
            .O(N__19925),
            .I(N__19912));
    LocalMux I__1862 (
            .O(N__19922),
            .I(N__19912));
    LocalMux I__1861 (
            .O(N__19919),
            .I(N__19912));
    Span4Mux_v I__1860 (
            .O(N__19912),
            .I(N__19909));
    Span4Mux_v I__1859 (
            .O(N__19909),
            .I(N__19906));
    Sp12to4 I__1858 (
            .O(N__19906),
            .I(N__19903));
    Odrv12 I__1857 (
            .O(N__19903),
            .I(RTD_DRDY));
    CascadeMux I__1856 (
            .O(N__19900),
            .I(\RTD.n11_cascade_ ));
    CascadeMux I__1855 (
            .O(N__19897),
            .I(\RTD.n19_cascade_ ));
    CEMux I__1854 (
            .O(N__19894),
            .I(N__19885));
    InMux I__1853 (
            .O(N__19893),
            .I(N__19872));
    InMux I__1852 (
            .O(N__19892),
            .I(N__19872));
    InMux I__1851 (
            .O(N__19891),
            .I(N__19872));
    InMux I__1850 (
            .O(N__19890),
            .I(N__19872));
    InMux I__1849 (
            .O(N__19889),
            .I(N__19872));
    InMux I__1848 (
            .O(N__19888),
            .I(N__19872));
    LocalMux I__1847 (
            .O(N__19885),
            .I(N__19867));
    LocalMux I__1846 (
            .O(N__19872),
            .I(N__19867));
    Odrv4 I__1845 (
            .O(N__19867),
            .I(n13151));
    CascadeMux I__1844 (
            .O(N__19864),
            .I(N__19860));
    InMux I__1843 (
            .O(N__19863),
            .I(N__19854));
    InMux I__1842 (
            .O(N__19860),
            .I(N__19854));
    InMux I__1841 (
            .O(N__19859),
            .I(N__19851));
    LocalMux I__1840 (
            .O(N__19854),
            .I(N__19848));
    LocalMux I__1839 (
            .O(N__19851),
            .I(\RTD.n1_adj_1393 ));
    Odrv4 I__1838 (
            .O(N__19848),
            .I(\RTD.n1_adj_1393 ));
    InMux I__1837 (
            .O(N__19843),
            .I(N__19840));
    LocalMux I__1836 (
            .O(N__19840),
            .I(\RTD.n19482 ));
    CascadeMux I__1835 (
            .O(N__19837),
            .I(\RTD.n19482_cascade_ ));
    CascadeMux I__1834 (
            .O(N__19834),
            .I(\RTD.n7285_cascade_ ));
    CascadeMux I__1833 (
            .O(N__19831),
            .I(\RTD.n21_cascade_ ));
    InMux I__1832 (
            .O(N__19828),
            .I(N__19825));
    LocalMux I__1831 (
            .O(N__19825),
            .I(N__19822));
    Odrv12 I__1830 (
            .O(N__19822),
            .I(\RTD.n4 ));
    CascadeMux I__1829 (
            .O(N__19819),
            .I(\RTD.n20969_cascade_ ));
    SRMux I__1828 (
            .O(N__19816),
            .I(N__19813));
    LocalMux I__1827 (
            .O(N__19813),
            .I(N__19809));
    SRMux I__1826 (
            .O(N__19812),
            .I(N__19806));
    Span4Mux_h I__1825 (
            .O(N__19809),
            .I(N__19801));
    LocalMux I__1824 (
            .O(N__19806),
            .I(N__19801));
    Odrv4 I__1823 (
            .O(N__19801),
            .I(\RTD.n15050 ));
    IoInMux I__1822 (
            .O(N__19798),
            .I(N__19795));
    LocalMux I__1821 (
            .O(N__19795),
            .I(N__19792));
    IoSpan4Mux I__1820 (
            .O(N__19792),
            .I(N__19789));
    Span4Mux_s3_h I__1819 (
            .O(N__19789),
            .I(N__19786));
    Span4Mux_v I__1818 (
            .O(N__19786),
            .I(N__19783));
    Sp12to4 I__1817 (
            .O(N__19783),
            .I(N__19780));
    Odrv12 I__1816 (
            .O(N__19780),
            .I(RTD_SDI));
    CEMux I__1815 (
            .O(N__19777),
            .I(N__19774));
    LocalMux I__1814 (
            .O(N__19774),
            .I(N__19771));
    Span4Mux_v I__1813 (
            .O(N__19771),
            .I(N__19768));
    Span4Mux_h I__1812 (
            .O(N__19768),
            .I(N__19765));
    Odrv4 I__1811 (
            .O(N__19765),
            .I(\RTD.n11704 ));
    CascadeMux I__1810 (
            .O(N__19762),
            .I(\RTD.n33_cascade_ ));
    CascadeMux I__1809 (
            .O(N__19759),
            .I(N__19752));
    CascadeMux I__1808 (
            .O(N__19758),
            .I(N__19746));
    CascadeMux I__1807 (
            .O(N__19757),
            .I(N__19741));
    CascadeMux I__1806 (
            .O(N__19756),
            .I(N__19738));
    InMux I__1805 (
            .O(N__19755),
            .I(N__19729));
    InMux I__1804 (
            .O(N__19752),
            .I(N__19726));
    InMux I__1803 (
            .O(N__19751),
            .I(N__19723));
    InMux I__1802 (
            .O(N__19750),
            .I(N__19720));
    InMux I__1801 (
            .O(N__19749),
            .I(N__19717));
    InMux I__1800 (
            .O(N__19746),
            .I(N__19712));
    InMux I__1799 (
            .O(N__19745),
            .I(N__19712));
    InMux I__1798 (
            .O(N__19744),
            .I(N__19703));
    InMux I__1797 (
            .O(N__19741),
            .I(N__19703));
    InMux I__1796 (
            .O(N__19738),
            .I(N__19703));
    InMux I__1795 (
            .O(N__19737),
            .I(N__19703));
    InMux I__1794 (
            .O(N__19736),
            .I(N__19692));
    InMux I__1793 (
            .O(N__19735),
            .I(N__19692));
    InMux I__1792 (
            .O(N__19734),
            .I(N__19692));
    InMux I__1791 (
            .O(N__19733),
            .I(N__19692));
    InMux I__1790 (
            .O(N__19732),
            .I(N__19692));
    LocalMux I__1789 (
            .O(N__19729),
            .I(N__19689));
    LocalMux I__1788 (
            .O(N__19726),
            .I(N__19674));
    LocalMux I__1787 (
            .O(N__19723),
            .I(N__19674));
    LocalMux I__1786 (
            .O(N__19720),
            .I(N__19674));
    LocalMux I__1785 (
            .O(N__19717),
            .I(N__19674));
    LocalMux I__1784 (
            .O(N__19712),
            .I(N__19674));
    LocalMux I__1783 (
            .O(N__19703),
            .I(N__19674));
    LocalMux I__1782 (
            .O(N__19692),
            .I(N__19674));
    Span4Mux_v I__1781 (
            .O(N__19689),
            .I(N__19669));
    Span4Mux_v I__1780 (
            .O(N__19674),
            .I(N__19669));
    Odrv4 I__1779 (
            .O(N__19669),
            .I(n1_adj_1575));
    InMux I__1778 (
            .O(N__19666),
            .I(N__19663));
    LocalMux I__1777 (
            .O(N__19663),
            .I(N__19660));
    Odrv12 I__1776 (
            .O(N__19660),
            .I(\RTD.n16614 ));
    CascadeMux I__1775 (
            .O(N__19657),
            .I(\RTD.n16614_cascade_ ));
    CascadeMux I__1774 (
            .O(N__19654),
            .I(N__19648));
    CascadeMux I__1773 (
            .O(N__19653),
            .I(N__19645));
    CascadeMux I__1772 (
            .O(N__19652),
            .I(N__19642));
    CascadeMux I__1771 (
            .O(N__19651),
            .I(N__19637));
    InMux I__1770 (
            .O(N__19648),
            .I(N__19626));
    InMux I__1769 (
            .O(N__19645),
            .I(N__19626));
    InMux I__1768 (
            .O(N__19642),
            .I(N__19626));
    InMux I__1767 (
            .O(N__19641),
            .I(N__19626));
    InMux I__1766 (
            .O(N__19640),
            .I(N__19626));
    InMux I__1765 (
            .O(N__19637),
            .I(N__19623));
    LocalMux I__1764 (
            .O(N__19626),
            .I(n14465));
    LocalMux I__1763 (
            .O(N__19623),
            .I(n14465));
    InMux I__1762 (
            .O(N__19618),
            .I(N__19613));
    InMux I__1761 (
            .O(N__19617),
            .I(N__19610));
    InMux I__1760 (
            .O(N__19616),
            .I(N__19607));
    LocalMux I__1759 (
            .O(N__19613),
            .I(read_buf_8));
    LocalMux I__1758 (
            .O(N__19610),
            .I(read_buf_8));
    LocalMux I__1757 (
            .O(N__19607),
            .I(read_buf_8));
    CascadeMux I__1756 (
            .O(N__19600),
            .I(N__19597));
    InMux I__1755 (
            .O(N__19597),
            .I(N__19592));
    InMux I__1754 (
            .O(N__19596),
            .I(N__19589));
    InMux I__1753 (
            .O(N__19595),
            .I(N__19586));
    LocalMux I__1752 (
            .O(N__19592),
            .I(read_buf_4));
    LocalMux I__1751 (
            .O(N__19589),
            .I(read_buf_4));
    LocalMux I__1750 (
            .O(N__19586),
            .I(read_buf_4));
    InMux I__1749 (
            .O(N__19579),
            .I(N__19569));
    InMux I__1748 (
            .O(N__19578),
            .I(N__19569));
    InMux I__1747 (
            .O(N__19577),
            .I(N__19563));
    InMux I__1746 (
            .O(N__19576),
            .I(N__19563));
    InMux I__1745 (
            .O(N__19575),
            .I(N__19553));
    InMux I__1744 (
            .O(N__19574),
            .I(N__19553));
    LocalMux I__1743 (
            .O(N__19569),
            .I(N__19547));
    InMux I__1742 (
            .O(N__19568),
            .I(N__19544));
    LocalMux I__1741 (
            .O(N__19563),
            .I(N__19541));
    InMux I__1740 (
            .O(N__19562),
            .I(N__19530));
    InMux I__1739 (
            .O(N__19561),
            .I(N__19530));
    InMux I__1738 (
            .O(N__19560),
            .I(N__19530));
    InMux I__1737 (
            .O(N__19559),
            .I(N__19530));
    InMux I__1736 (
            .O(N__19558),
            .I(N__19530));
    LocalMux I__1735 (
            .O(N__19553),
            .I(N__19527));
    InMux I__1734 (
            .O(N__19552),
            .I(N__19520));
    InMux I__1733 (
            .O(N__19551),
            .I(N__19520));
    InMux I__1732 (
            .O(N__19550),
            .I(N__19520));
    Odrv4 I__1731 (
            .O(N__19547),
            .I(n13279));
    LocalMux I__1730 (
            .O(N__19544),
            .I(n13279));
    Odrv4 I__1729 (
            .O(N__19541),
            .I(n13279));
    LocalMux I__1728 (
            .O(N__19530),
            .I(n13279));
    Odrv4 I__1727 (
            .O(N__19527),
            .I(n13279));
    LocalMux I__1726 (
            .O(N__19520),
            .I(n13279));
    InMux I__1725 (
            .O(N__19507),
            .I(N__19500));
    InMux I__1724 (
            .O(N__19506),
            .I(N__19500));
    InMux I__1723 (
            .O(N__19505),
            .I(N__19497));
    LocalMux I__1722 (
            .O(N__19500),
            .I(read_buf_2));
    LocalMux I__1721 (
            .O(N__19497),
            .I(read_buf_2));
    CascadeMux I__1720 (
            .O(N__19492),
            .I(N__19488));
    InMux I__1719 (
            .O(N__19491),
            .I(N__19484));
    InMux I__1718 (
            .O(N__19488),
            .I(N__19479));
    InMux I__1717 (
            .O(N__19487),
            .I(N__19479));
    LocalMux I__1716 (
            .O(N__19484),
            .I(read_buf_3));
    LocalMux I__1715 (
            .O(N__19479),
            .I(read_buf_3));
    CascadeMux I__1714 (
            .O(N__19474),
            .I(N__19469));
    InMux I__1713 (
            .O(N__19473),
            .I(N__19461));
    InMux I__1712 (
            .O(N__19472),
            .I(N__19461));
    InMux I__1711 (
            .O(N__19469),
            .I(N__19448));
    InMux I__1710 (
            .O(N__19468),
            .I(N__19448));
    InMux I__1709 (
            .O(N__19467),
            .I(N__19448));
    InMux I__1708 (
            .O(N__19466),
            .I(N__19448));
    LocalMux I__1707 (
            .O(N__19461),
            .I(N__19444));
    InMux I__1706 (
            .O(N__19460),
            .I(N__19437));
    InMux I__1705 (
            .O(N__19459),
            .I(N__19437));
    InMux I__1704 (
            .O(N__19458),
            .I(N__19437));
    InMux I__1703 (
            .O(N__19457),
            .I(N__19434));
    LocalMux I__1702 (
            .O(N__19448),
            .I(N__19427));
    InMux I__1701 (
            .O(N__19447),
            .I(N__19424));
    Span4Mux_v I__1700 (
            .O(N__19444),
            .I(N__19417));
    LocalMux I__1699 (
            .O(N__19437),
            .I(N__19417));
    LocalMux I__1698 (
            .O(N__19434),
            .I(N__19417));
    InMux I__1697 (
            .O(N__19433),
            .I(N__19410));
    InMux I__1696 (
            .O(N__19432),
            .I(N__19410));
    InMux I__1695 (
            .O(N__19431),
            .I(N__19410));
    InMux I__1694 (
            .O(N__19430),
            .I(N__19407));
    Odrv12 I__1693 (
            .O(N__19427),
            .I(n11700));
    LocalMux I__1692 (
            .O(N__19424),
            .I(n11700));
    Odrv4 I__1691 (
            .O(N__19417),
            .I(n11700));
    LocalMux I__1690 (
            .O(N__19410),
            .I(n11700));
    LocalMux I__1689 (
            .O(N__19407),
            .I(n11700));
    CEMux I__1688 (
            .O(N__19396),
            .I(N__19393));
    LocalMux I__1687 (
            .O(N__19393),
            .I(N__19390));
    Span4Mux_h I__1686 (
            .O(N__19390),
            .I(N__19386));
    CEMux I__1685 (
            .O(N__19389),
            .I(N__19383));
    Odrv4 I__1684 (
            .O(N__19386),
            .I(\RTD.n11726 ));
    LocalMux I__1683 (
            .O(N__19383),
            .I(\RTD.n11726 ));
    InMux I__1682 (
            .O(N__19378),
            .I(N__19373));
    InMux I__1681 (
            .O(N__19377),
            .I(N__19370));
    InMux I__1680 (
            .O(N__19376),
            .I(N__19367));
    LocalMux I__1679 (
            .O(N__19373),
            .I(read_buf_13));
    LocalMux I__1678 (
            .O(N__19370),
            .I(read_buf_13));
    LocalMux I__1677 (
            .O(N__19367),
            .I(read_buf_13));
    CascadeMux I__1676 (
            .O(N__19360),
            .I(N__19356));
    InMux I__1675 (
            .O(N__19359),
            .I(N__19348));
    InMux I__1674 (
            .O(N__19356),
            .I(N__19348));
    InMux I__1673 (
            .O(N__19355),
            .I(N__19348));
    LocalMux I__1672 (
            .O(N__19348),
            .I(read_buf_9));
    InMux I__1671 (
            .O(N__19345),
            .I(N__19339));
    InMux I__1670 (
            .O(N__19344),
            .I(N__19339));
    LocalMux I__1669 (
            .O(N__19339),
            .I(adress_1));
    InMux I__1668 (
            .O(N__19336),
            .I(N__19330));
    InMux I__1667 (
            .O(N__19335),
            .I(N__19330));
    LocalMux I__1666 (
            .O(N__19330),
            .I(adress_2));
    CascadeMux I__1665 (
            .O(N__19327),
            .I(N__19323));
    InMux I__1664 (
            .O(N__19326),
            .I(N__19318));
    InMux I__1663 (
            .O(N__19323),
            .I(N__19318));
    LocalMux I__1662 (
            .O(N__19318),
            .I(adress_3));
    InMux I__1661 (
            .O(N__19315),
            .I(N__19309));
    InMux I__1660 (
            .O(N__19314),
            .I(N__19309));
    LocalMux I__1659 (
            .O(N__19309),
            .I(N__19306));
    Odrv4 I__1658 (
            .O(N__19306),
            .I(adress_4));
    CascadeMux I__1657 (
            .O(N__19303),
            .I(N__19299));
    InMux I__1656 (
            .O(N__19302),
            .I(N__19294));
    InMux I__1655 (
            .O(N__19299),
            .I(N__19294));
    LocalMux I__1654 (
            .O(N__19294),
            .I(adress_5));
    CascadeMux I__1653 (
            .O(N__19291),
            .I(N__19287));
    InMux I__1652 (
            .O(N__19290),
            .I(N__19283));
    InMux I__1651 (
            .O(N__19287),
            .I(N__19280));
    InMux I__1650 (
            .O(N__19286),
            .I(N__19277));
    LocalMux I__1649 (
            .O(N__19283),
            .I(read_buf_10));
    LocalMux I__1648 (
            .O(N__19280),
            .I(read_buf_10));
    LocalMux I__1647 (
            .O(N__19277),
            .I(read_buf_10));
    InMux I__1646 (
            .O(N__19270),
            .I(N__19265));
    CascadeMux I__1645 (
            .O(N__19269),
            .I(N__19262));
    CascadeMux I__1644 (
            .O(N__19268),
            .I(N__19259));
    LocalMux I__1643 (
            .O(N__19265),
            .I(N__19256));
    InMux I__1642 (
            .O(N__19262),
            .I(N__19251));
    InMux I__1641 (
            .O(N__19259),
            .I(N__19251));
    Odrv4 I__1640 (
            .O(N__19256),
            .I(read_buf_11));
    LocalMux I__1639 (
            .O(N__19251),
            .I(read_buf_11));
    CascadeMux I__1638 (
            .O(N__19246),
            .I(n11700_cascade_));
    CascadeMux I__1637 (
            .O(N__19243),
            .I(N__19240));
    InMux I__1636 (
            .O(N__19240),
            .I(N__19233));
    InMux I__1635 (
            .O(N__19239),
            .I(N__19233));
    InMux I__1634 (
            .O(N__19238),
            .I(N__19230));
    LocalMux I__1633 (
            .O(N__19233),
            .I(read_buf_14));
    LocalMux I__1632 (
            .O(N__19230),
            .I(read_buf_14));
    InMux I__1631 (
            .O(N__19225),
            .I(N__19219));
    InMux I__1630 (
            .O(N__19224),
            .I(N__19219));
    LocalMux I__1629 (
            .O(N__19219),
            .I(read_buf_15));
    CascadeMux I__1628 (
            .O(N__19216),
            .I(N__19213));
    InMux I__1627 (
            .O(N__19213),
            .I(N__19210));
    LocalMux I__1626 (
            .O(N__19210),
            .I(N__19205));
    InMux I__1625 (
            .O(N__19209),
            .I(N__19202));
    InMux I__1624 (
            .O(N__19208),
            .I(N__19199));
    Odrv12 I__1623 (
            .O(N__19205),
            .I(read_buf_1));
    LocalMux I__1622 (
            .O(N__19202),
            .I(read_buf_1));
    LocalMux I__1621 (
            .O(N__19199),
            .I(read_buf_1));
    InMux I__1620 (
            .O(N__19192),
            .I(N__19187));
    InMux I__1619 (
            .O(N__19191),
            .I(N__19182));
    InMux I__1618 (
            .O(N__19190),
            .I(N__19182));
    LocalMux I__1617 (
            .O(N__19187),
            .I(read_buf_0));
    LocalMux I__1616 (
            .O(N__19182),
            .I(read_buf_0));
    InMux I__1615 (
            .O(N__19177),
            .I(N__19172));
    InMux I__1614 (
            .O(N__19176),
            .I(N__19167));
    InMux I__1613 (
            .O(N__19175),
            .I(N__19167));
    LocalMux I__1612 (
            .O(N__19172),
            .I(read_buf_5));
    LocalMux I__1611 (
            .O(N__19167),
            .I(read_buf_5));
    CascadeMux I__1610 (
            .O(N__19162),
            .I(N__19158));
    InMux I__1609 (
            .O(N__19161),
            .I(N__19154));
    InMux I__1608 (
            .O(N__19158),
            .I(N__19149));
    InMux I__1607 (
            .O(N__19157),
            .I(N__19149));
    LocalMux I__1606 (
            .O(N__19154),
            .I(read_buf_12));
    LocalMux I__1605 (
            .O(N__19149),
            .I(read_buf_12));
    CascadeMux I__1604 (
            .O(N__19144),
            .I(N__19141));
    InMux I__1603 (
            .O(N__19141),
            .I(N__19135));
    InMux I__1602 (
            .O(N__19140),
            .I(N__19135));
    LocalMux I__1601 (
            .O(N__19135),
            .I(N__19131));
    InMux I__1600 (
            .O(N__19134),
            .I(N__19128));
    Odrv4 I__1599 (
            .O(N__19131),
            .I(read_buf_6));
    LocalMux I__1598 (
            .O(N__19128),
            .I(read_buf_6));
    InMux I__1597 (
            .O(N__19123),
            .I(N__19119));
    CascadeMux I__1596 (
            .O(N__19122),
            .I(N__19116));
    LocalMux I__1595 (
            .O(N__19119),
            .I(N__19112));
    InMux I__1594 (
            .O(N__19116),
            .I(N__19109));
    InMux I__1593 (
            .O(N__19115),
            .I(N__19106));
    Odrv4 I__1592 (
            .O(N__19112),
            .I(read_buf_7));
    LocalMux I__1591 (
            .O(N__19109),
            .I(read_buf_7));
    LocalMux I__1590 (
            .O(N__19106),
            .I(read_buf_7));
    IoInMux I__1589 (
            .O(N__19099),
            .I(N__19096));
    LocalMux I__1588 (
            .O(N__19096),
            .I(N__19093));
    IoSpan4Mux I__1587 (
            .O(N__19093),
            .I(N__19090));
    Span4Mux_s3_h I__1586 (
            .O(N__19090),
            .I(N__19087));
    Span4Mux_v I__1585 (
            .O(N__19087),
            .I(N__19084));
    Span4Mux_v I__1584 (
            .O(N__19084),
            .I(N__19081));
    Odrv4 I__1583 (
            .O(N__19081),
            .I(RTD_CS));
    CEMux I__1582 (
            .O(N__19078),
            .I(N__19075));
    LocalMux I__1581 (
            .O(N__19075),
            .I(N__19072));
    Odrv12 I__1580 (
            .O(N__19072),
            .I(\RTD.n11673 ));
    CascadeMux I__1579 (
            .O(N__19069),
            .I(n13279_cascade_));
    CascadeMux I__1578 (
            .O(N__19066),
            .I(N__19063));
    InMux I__1577 (
            .O(N__19063),
            .I(N__19060));
    LocalMux I__1576 (
            .O(N__19060),
            .I(N__19057));
    Span4Mux_h I__1575 (
            .O(N__19057),
            .I(N__19054));
    Sp12to4 I__1574 (
            .O(N__19054),
            .I(N__19051));
    Span12Mux_v I__1573 (
            .O(N__19051),
            .I(N__19048));
    Odrv12 I__1572 (
            .O(N__19048),
            .I(RTD_SDO));
    IoInMux I__1571 (
            .O(N__19045),
            .I(N__19042));
    LocalMux I__1570 (
            .O(N__19042),
            .I(N__19039));
    IoSpan4Mux I__1569 (
            .O(N__19039),
            .I(N__19036));
    Span4Mux_s3_h I__1568 (
            .O(N__19036),
            .I(N__19033));
    Span4Mux_v I__1567 (
            .O(N__19033),
            .I(N__19030));
    Odrv4 I__1566 (
            .O(N__19030),
            .I(RTD_SCLK));
    CEMux I__1565 (
            .O(N__19027),
            .I(N__19024));
    LocalMux I__1564 (
            .O(N__19024),
            .I(N__19021));
    Odrv4 I__1563 (
            .O(N__19021),
            .I(\RTD.n8 ));
    IoInMux I__1562 (
            .O(N__19018),
            .I(N__19015));
    LocalMux I__1561 (
            .O(N__19015),
            .I(N__19012));
    IoSpan4Mux I__1560 (
            .O(N__19012),
            .I(N__19009));
    IoSpan4Mux I__1559 (
            .O(N__19009),
            .I(N__19006));
    Odrv4 I__1558 (
            .O(N__19006),
            .I(ICE_SYSCLK));
    IoInMux I__1557 (
            .O(N__19003),
            .I(N__19000));
    LocalMux I__1556 (
            .O(N__19000),
            .I(N__18997));
    IoSpan4Mux I__1555 (
            .O(N__18997),
            .I(N__18994));
    Span4Mux_s3_v I__1554 (
            .O(N__18994),
            .I(N__18991));
    Sp12to4 I__1553 (
            .O(N__18991),
            .I(N__18988));
    Span12Mux_h I__1552 (
            .O(N__18988),
            .I(N__18985));
    Odrv12 I__1551 (
            .O(N__18985),
            .I(ICE_GPMO_2));
    INV INVdds0_mclkcnt_i7_3772__i0C (
            .O(INVdds0_mclkcnt_i7_3772__i0C_net),
            .I(N__56030));
    INV INVdds0_mclk_294C (
            .O(INVdds0_mclk_294C_net),
            .I(N__56029));
    INV INVdata_cntvec_i0_i8C (
            .O(INVdata_cntvec_i0_i8C_net),
            .I(N__55186));
    INV INVdata_cntvec_i0_i0C (
            .O(INVdata_cntvec_i0_i0C_net),
            .I(N__55172));
    INV \INVcomm_spi.data_valid_85C  (
            .O(\INVcomm_spi.data_valid_85C_net ),
            .I(N__55130));
    INV \INVcomm_spi.MISO_48_12187_12188_resetC  (
            .O(\INVcomm_spi.MISO_48_12187_12188_resetC_net ),
            .I(N__55090));
    INV \INVcomm_spi.imiso_83_12193_12194_resetC  (
            .O(\INVcomm_spi.imiso_83_12193_12194_resetC_net ),
            .I(N__52368));
    INV INVdata_count_i0_i8C (
            .O(INVdata_count_i0_i8C_net),
            .I(N__55211));
    INV INVdata_count_i0_i0C (
            .O(INVdata_count_i0_i0C_net),
            .I(N__55198));
    INV \INVcomm_spi.MISO_48_12187_12188_setC  (
            .O(\INVcomm_spi.MISO_48_12187_12188_setC_net ),
            .I(N__55078));
    INV \INVADC_VDC.genclk.t0on_i8C  (
            .O(\INVADC_VDC.genclk.t0on_i8C_net ),
            .I(N__56022));
    INV \INVADC_VDC.genclk.t0on_i0C  (
            .O(\INVADC_VDC.genclk.t0on_i0C_net ),
            .I(N__56018));
    INV \INVADC_VDC.genclk.div_state_i1C  (
            .O(\INVADC_VDC.genclk.div_state_i1C_net ),
            .I(N__56023));
    INV INVacadc_skipcnt_i0_i9C (
            .O(INVacadc_skipcnt_i0_i9C_net),
            .I(N__55182));
    INV INVacadc_skipcnt_i0_i1C (
            .O(INVacadc_skipcnt_i0_i1C_net),
            .I(N__55167));
    INV INVacadc_skipcnt_i0_i0C (
            .O(INVacadc_skipcnt_i0_i0C_net),
            .I(N__55152));
    INV \INVcomm_spi.bit_cnt_3767__i1C  (
            .O(\INVcomm_spi.bit_cnt_3767__i1C_net ),
            .I(N__52414));
    INV \INVcomm_spi.imiso_83_12193_12194_setC  (
            .O(\INVcomm_spi.imiso_83_12193_12194_setC_net ),
            .I(N__52413));
    INV \INVADC_VDC.genclk.t_clk_24C  (
            .O(\INVADC_VDC.genclk.t_clk_24C_net ),
            .I(N__56016));
    INV INVacadc_trig_300C (
            .O(INVacadc_trig_300C_net),
            .I(N__55181));
    INV INVeis_state_i0C (
            .O(INVeis_state_i0C_net),
            .I(N__55117));
    INV \INVADC_VDC.genclk.t0off_i8C  (
            .O(\INVADC_VDC.genclk.t0off_i8C_net ),
            .I(N__56017));
    INV \INVADC_VDC.genclk.t0off_i0C  (
            .O(\INVADC_VDC.genclk.t0off_i0C_net ),
            .I(N__56015));
    INV INViac_raw_buf_vac_raw_buf_merged2WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged2WCLKN_net),
            .I(N__55159));
    INV INViac_raw_buf_vac_raw_buf_merged7WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged7WCLKN_net),
            .I(N__55246));
    INV INViac_raw_buf_vac_raw_buf_merged1WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged1WCLKN_net),
            .I(N__55092));
    INV INViac_raw_buf_vac_raw_buf_merged6WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged6WCLKN_net),
            .I(N__55243));
    INV INViac_raw_buf_vac_raw_buf_merged0WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged0WCLKN_net),
            .I(N__55080));
    INV INViac_raw_buf_vac_raw_buf_merged5WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged5WCLKN_net),
            .I(N__55236));
    INV INViac_raw_buf_vac_raw_buf_merged9WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged9WCLKN_net),
            .I(N__55226));
    INV INViac_raw_buf_vac_raw_buf_merged4WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged4WCLKN_net),
            .I(N__55215));
    INV INViac_raw_buf_vac_raw_buf_merged8WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged8WCLKN_net),
            .I(N__55203));
    INV INViac_raw_buf_vac_raw_buf_merged10WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged10WCLKN_net),
            .I(N__55111));
    INV INViac_raw_buf_vac_raw_buf_merged3WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged3WCLKN_net),
            .I(N__55189));
    INV INViac_raw_buf_vac_raw_buf_merged11WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged11WCLKN_net),
            .I(N__55132));
    defparam IN_MUX_bfv_17_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_17_9_0_));
    defparam IN_MUX_bfv_17_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_10_0_ (
            .carryinitin(n19454),
            .carryinitout(bfn_17_10_0_));
    defparam IN_MUX_bfv_17_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_17_11_0_ (
            .carryinitin(n19462),
            .carryinitout(bfn_17_11_0_));
    defparam IN_MUX_bfv_22_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_22_11_0_));
    defparam IN_MUX_bfv_13_16_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_16_0_));
    defparam IN_MUX_bfv_13_17_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_17_0_ (
            .carryinitin(n19311_THRU_CRY_6_THRU_CO),
            .carryinitout(bfn_13_17_0_));
    defparam IN_MUX_bfv_13_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_18_0_ (
            .carryinitin(n19319),
            .carryinitout(bfn_13_18_0_));
    defparam IN_MUX_bfv_18_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_12_0_));
    defparam IN_MUX_bfv_18_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_13_0_ (
            .carryinitin(n19303),
            .carryinitout(bfn_18_13_0_));
    defparam IN_MUX_bfv_15_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_17_0_));
    defparam IN_MUX_bfv_15_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_18_0_ (
            .carryinitin(n19294),
            .carryinitout(bfn_15_18_0_));
    defparam IN_MUX_bfv_12_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_12_0_));
    defparam IN_MUX_bfv_12_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_13_0_ (
            .carryinitin(n19342),
            .carryinitout(bfn_12_13_0_));
    defparam IN_MUX_bfv_16_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_16_15_0_));
    defparam IN_MUX_bfv_16_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_16_16_0_ (
            .carryinitin(n19333),
            .carryinitout(bfn_16_16_0_));
    defparam IN_MUX_bfv_11_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_3_0_));
    defparam IN_MUX_bfv_11_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_4_0_ (
            .carryinitin(\ADC_VDC.genclk.n19417 ),
            .carryinitout(bfn_11_4_0_));
    defparam IN_MUX_bfv_15_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_3_0_));
    defparam IN_MUX_bfv_15_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_4_0_ (
            .carryinitin(\ADC_VDC.genclk.n19432 ),
            .carryinitout(bfn_15_4_0_));
    defparam IN_MUX_bfv_13_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_6_0_));
    defparam IN_MUX_bfv_11_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_7_0_));
    defparam IN_MUX_bfv_11_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_8_0_ (
            .carryinitin(\ADC_VDC.n19406 ),
            .carryinitout(bfn_11_8_0_));
    defparam IN_MUX_bfv_9_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_5_0_));
    defparam IN_MUX_bfv_9_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_6_0_ (
            .carryinitin(\ADC_VDC.n19371 ),
            .carryinitout(bfn_9_6_0_));
    defparam IN_MUX_bfv_9_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_7_0_ (
            .carryinitin(\ADC_VDC.n19379 ),
            .carryinitout(bfn_9_7_0_));
    defparam IN_MUX_bfv_9_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_8_0_ (
            .carryinitin(\ADC_VDC.n19387 ),
            .carryinitout(bfn_9_8_0_));
    defparam IN_MUX_bfv_9_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_9_0_ (
            .carryinitin(\ADC_VDC.n19395 ),
            .carryinitout(bfn_9_9_0_));
    defparam IN_MUX_bfv_7_17_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_17_0_));
    defparam IN_MUX_bfv_7_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_19_0_));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \RTD.SCLK_51_LC_2_5_0 .C_ON=1'b0;
    defparam \RTD.SCLK_51_LC_2_5_0 .SEQ_MODE=4'b1000;
    defparam \RTD.SCLK_51_LC_2_5_0 .LUT_INIT=16'b0010110000110110;
    LogicCell40 \RTD.SCLK_51_LC_2_5_0  (
            .in0(N__22257),
            .in1(N__22114),
            .in2(N__22410),
            .in3(N__20970),
            .lcout(RTD_SCLK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41081),
            .ce(N__19027),
            .sr(_gnd_net_));
    defparam \RTD.i19108_4_lut_4_lut_LC_2_5_1 .C_ON=1'b0;
    defparam \RTD.i19108_4_lut_4_lut_LC_2_5_1 .SEQ_MODE=4'b0000;
    defparam \RTD.i19108_4_lut_4_lut_LC_2_5_1 .LUT_INIT=16'b1111011110111111;
    LogicCell40 \RTD.i19108_4_lut_4_lut_LC_2_5_1  (
            .in0(N__20969),
            .in1(N__22393),
            .in2(N__22132),
            .in3(N__22255),
            .lcout(\RTD.n8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i27_4_lut_4_lut_LC_2_5_2 .C_ON=1'b0;
    defparam \RTD.i27_4_lut_4_lut_LC_2_5_2 .SEQ_MODE=4'b0000;
    defparam \RTD.i27_4_lut_4_lut_LC_2_5_2 .LUT_INIT=16'b1100110010000110;
    LogicCell40 \RTD.i27_4_lut_4_lut_LC_2_5_2  (
            .in0(N__22254),
            .in1(N__22109),
            .in2(N__22409),
            .in3(N__20968),
            .lcout(\RTD.n11704 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i19151_4_lut_4_lut_LC_2_5_3 .C_ON=1'b0;
    defparam \RTD.i19151_4_lut_4_lut_LC_2_5_3 .SEQ_MODE=4'b0000;
    defparam \RTD.i19151_4_lut_4_lut_LC_2_5_3 .LUT_INIT=16'b1101001110101100;
    LogicCell40 \RTD.i19151_4_lut_4_lut_LC_2_5_3  (
            .in0(N__20966),
            .in1(N__22394),
            .in2(N__22131),
            .in3(N__22253),
            .lcout(\RTD.n11726 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_3_lut_4_lut_adj_25_LC_2_5_4 .C_ON=1'b0;
    defparam \RTD.i1_3_lut_4_lut_adj_25_LC_2_5_4 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_3_lut_4_lut_adj_25_LC_2_5_4 .LUT_INIT=16'b1100010010010010;
    LogicCell40 \RTD.i1_3_lut_4_lut_adj_25_LC_2_5_4  (
            .in0(N__22252),
            .in1(N__22105),
            .in2(N__22408),
            .in3(N__20967),
            .lcout(\RTD.n15050 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i19070_3_lut_3_lut_LC_2_5_7 .C_ON=1'b0;
    defparam \RTD.i19070_3_lut_3_lut_LC_2_5_7 .SEQ_MODE=4'b0000;
    defparam \RTD.i19070_3_lut_3_lut_LC_2_5_7 .LUT_INIT=16'b1000100010011001;
    LogicCell40 \RTD.i19070_3_lut_3_lut_LC_2_5_7  (
            .in0(N__22113),
            .in1(N__22395),
            .in2(_gnd_net_),
            .in3(N__22256),
            .lcout(\RTD.n11673 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.CS_52_LC_2_7_5 .C_ON=1'b0;
    defparam \RTD.CS_52_LC_2_7_5 .SEQ_MODE=4'b1000;
    defparam \RTD.CS_52_LC_2_7_5 .LUT_INIT=16'b0000011101010111;
    LogicCell40 \RTD.CS_52_LC_2_7_5  (
            .in0(N__20964),
            .in1(N__19666),
            .in2(N__22411),
            .in3(N__22258),
            .lcout(RTD_CS),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41131),
            .ce(N__19078),
            .sr(_gnd_net_));
    defparam \RTD.i1_4_lut_4_lut_adj_21_LC_2_8_0 .C_ON=1'b0;
    defparam \RTD.i1_4_lut_4_lut_adj_21_LC_2_8_0 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_4_lut_4_lut_adj_21_LC_2_8_0 .LUT_INIT=16'b1101100100000001;
    LogicCell40 \RTD.i1_4_lut_4_lut_adj_21_LC_2_8_0  (
            .in0(N__22259),
            .in1(N__22118),
            .in2(N__20977),
            .in3(N__22403),
            .lcout(n13279),
            .ltout(n13279_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i14_LC_2_8_1 .C_ON=1'b0;
    defparam \RTD.read_buf_i14_LC_2_8_1 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i14_LC_2_8_1 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \RTD.read_buf_i14_LC_2_8_1  (
            .in0(N__19377),
            .in1(N__19238),
            .in2(N__19069),
            .in3(N__19744),
            .lcout(read_buf_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41143),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i7_LC_2_8_3 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i7_LC_2_8_3 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i7_LC_2_8_3 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \RTD.READ_DATA_i7_LC_2_8_3  (
            .in0(N__22119),
            .in1(N__19447),
            .in2(N__20022),
            .in3(N__19123),
            .lcout(buf_readRTD_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41143),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i1_LC_2_8_4 .C_ON=1'b0;
    defparam \RTD.read_buf_i1_LC_2_8_4 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i1_LC_2_8_4 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \RTD.read_buf_i1_LC_2_8_4  (
            .in0(N__19551),
            .in1(N__19191),
            .in2(N__19756),
            .in3(N__19208),
            .lcout(read_buf_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41143),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i6_LC_2_8_6 .C_ON=1'b0;
    defparam \RTD.read_buf_i6_LC_2_8_6 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i6_LC_2_8_6 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \RTD.read_buf_i6_LC_2_8_6  (
            .in0(N__19552),
            .in1(N__19177),
            .in2(N__19757),
            .in3(N__19134),
            .lcout(read_buf_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41143),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i0_LC_2_8_7 .C_ON=1'b0;
    defparam \RTD.read_buf_i0_LC_2_8_7 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i0_LC_2_8_7 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \RTD.read_buf_i0_LC_2_8_7  (
            .in0(N__19190),
            .in1(N__19737),
            .in2(N__19066),
            .in3(N__19550),
            .lcout(read_buf_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41143),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i11_LC_2_9_0 .C_ON=1'b0;
    defparam \RTD.read_buf_i11_LC_2_9_0 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i11_LC_2_9_0 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \RTD.read_buf_i11_LC_2_9_0  (
            .in0(N__19733),
            .in1(N__19286),
            .in2(N__19268),
            .in3(N__19558),
            .lcout(read_buf_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41080),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i13_LC_2_9_1 .C_ON=1'b0;
    defparam \RTD.read_buf_i13_LC_2_9_1 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i13_LC_2_9_1 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \RTD.read_buf_i13_LC_2_9_1  (
            .in0(N__19560),
            .in1(N__19376),
            .in2(N__19162),
            .in3(N__19736),
            .lcout(read_buf_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41080),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i5_LC_2_9_2 .C_ON=1'b0;
    defparam \RTD.read_buf_i5_LC_2_9_2 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i5_LC_2_9_2 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \RTD.read_buf_i5_LC_2_9_2  (
            .in0(N__19735),
            .in1(N__19175),
            .in2(N__19600),
            .in3(N__19561),
            .lcout(read_buf_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41080),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i8_LC_2_9_3 .C_ON=1'b0;
    defparam \RTD.read_buf_i8_LC_2_9_3 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i8_LC_2_9_3 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \RTD.read_buf_i8_LC_2_9_3  (
            .in0(N__19562),
            .in1(N__19616),
            .in2(N__19122),
            .in3(N__19732),
            .lcout(read_buf_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41080),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i12_LC_2_9_4 .C_ON=1'b0;
    defparam \RTD.read_buf_i12_LC_2_9_4 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i12_LC_2_9_4 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \RTD.read_buf_i12_LC_2_9_4  (
            .in0(N__19734),
            .in1(N__19157),
            .in2(N__19269),
            .in3(N__19559),
            .lcout(read_buf_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41080),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i0_LC_2_9_5 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i0_LC_2_9_5 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i0_LC_2_9_5 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \RTD.READ_DATA_i0_LC_2_9_5  (
            .in0(N__22120),
            .in1(N__19192),
            .in2(N__21366),
            .in3(N__19458),
            .lcout(buf_readRTD_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41080),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i5_LC_2_9_6 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i5_LC_2_9_6 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i5_LC_2_9_6 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \RTD.READ_DATA_i5_LC_2_9_6  (
            .in0(N__19460),
            .in1(N__19176),
            .in2(N__20280),
            .in3(N__22122),
            .lcout(buf_readRTD_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41080),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i12_LC_2_9_7 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i12_LC_2_9_7 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i12_LC_2_9_7 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \RTD.READ_DATA_i12_LC_2_9_7  (
            .in0(N__22121),
            .in1(N__19161),
            .in2(N__25746),
            .in3(N__19459),
            .lcout(buf_readRTD_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41080),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i6_LC_2_10_0 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i6_LC_2_10_0 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i6_LC_2_10_0 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \RTD.READ_DATA_i6_LC_2_10_0  (
            .in0(N__19140),
            .in1(N__19473),
            .in2(N__29607),
            .in3(N__22129),
            .lcout(buf_readRTD_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41130),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i7_LC_2_10_2 .C_ON=1'b0;
    defparam \RTD.read_buf_i7_LC_2_10_2 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i7_LC_2_10_2 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \RTD.read_buf_i7_LC_2_10_2  (
            .in0(N__19577),
            .in1(N__19115),
            .in2(N__19144),
            .in3(N__19755),
            .lcout(read_buf_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41130),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i2_LC_2_10_3 .C_ON=1'b0;
    defparam \RTD.read_buf_i2_LC_2_10_3 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i2_LC_2_10_3 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \RTD.read_buf_i2_LC_2_10_3  (
            .in0(N__19505),
            .in1(N__19576),
            .in2(N__19216),
            .in3(N__19751),
            .lcout(read_buf_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41130),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i11_LC_2_10_4 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i11_LC_2_10_4 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i11_LC_2_10_4 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \RTD.READ_DATA_i11_LC_2_10_4  (
            .in0(N__19270),
            .in1(N__19472),
            .in2(N__21096),
            .in3(N__22128),
            .lcout(buf_readRTD_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41130),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.bit_cnt_3771__i3_LC_3_5_3 .C_ON=1'b0;
    defparam \RTD.bit_cnt_3771__i3_LC_3_5_3 .SEQ_MODE=4'b1000;
    defparam \RTD.bit_cnt_3771__i3_LC_3_5_3 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \RTD.bit_cnt_3771__i3_LC_3_5_3  (
            .in0(N__20596),
            .in1(N__20566),
            .in2(N__20517),
            .in3(N__20620),
            .lcout(\RTD.bit_cnt_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41132),
            .ce(N__19389),
            .sr(N__19812));
    defparam \RTD.i1_4_lut_4_lut_adj_22_LC_3_7_0 .C_ON=1'b0;
    defparam \RTD.i1_4_lut_4_lut_adj_22_LC_3_7_0 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_4_lut_4_lut_adj_22_LC_3_7_0 .LUT_INIT=16'b1110000010000000;
    LogicCell40 \RTD.i1_4_lut_4_lut_adj_22_LC_3_7_0  (
            .in0(N__22246),
            .in1(N__22115),
            .in2(N__22402),
            .in3(N__20963),
            .lcout(n11700),
            .ltout(n11700_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i14_LC_3_7_1 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i14_LC_3_7_1 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i14_LC_3_7_1 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \RTD.READ_DATA_i14_LC_3_7_1  (
            .in0(N__22116),
            .in1(N__23415),
            .in2(N__19246),
            .in3(N__19239),
            .lcout(buf_readRTD_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41115),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i15_LC_3_7_3 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i15_LC_3_7_3 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i15_LC_3_7_3 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \RTD.READ_DATA_i15_LC_3_7_3  (
            .in0(N__22117),
            .in1(N__19225),
            .in2(N__22452),
            .in3(N__19430),
            .lcout(buf_readRTD_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41115),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i15_LC_3_7_4 .C_ON=1'b0;
    defparam \RTD.read_buf_i15_LC_3_7_4 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i15_LC_3_7_4 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \RTD.read_buf_i15_LC_3_7_4  (
            .in0(N__19224),
            .in1(N__19749),
            .in2(N__19243),
            .in3(N__19568),
            .lcout(read_buf_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41115),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i1_LC_3_8_1 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i1_LC_3_8_1 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i1_LC_3_8_1 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \RTD.READ_DATA_i1_LC_3_8_1  (
            .in0(N__22093),
            .in1(N__19432),
            .in2(N__35325),
            .in3(N__19209),
            .lcout(buf_readRTD_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41141),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i9_LC_3_8_2 .C_ON=1'b0;
    defparam \RTD.read_buf_i9_LC_3_8_2 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i9_LC_3_8_2 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \RTD.read_buf_i9_LC_3_8_2  (
            .in0(N__19575),
            .in1(N__19618),
            .in2(N__19758),
            .in3(N__19355),
            .lcout(read_buf_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41141),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i10_LC_3_8_3 .C_ON=1'b0;
    defparam \RTD.read_buf_i10_LC_3_8_3 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i10_LC_3_8_3 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \RTD.read_buf_i10_LC_3_8_3  (
            .in0(N__19359),
            .in1(N__19745),
            .in2(N__19291),
            .in3(N__19574),
            .lcout(read_buf_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41141),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i13_LC_3_8_4 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i13_LC_3_8_4 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i13_LC_3_8_4 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \RTD.READ_DATA_i13_LC_3_8_4  (
            .in0(N__19431),
            .in1(N__19378),
            .in2(N__22518),
            .in3(N__22095),
            .lcout(buf_readRTD_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41141),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i9_LC_3_8_5 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i9_LC_3_8_5 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i9_LC_3_8_5 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \RTD.READ_DATA_i9_LC_3_8_5  (
            .in0(N__22094),
            .in1(N__19433),
            .in2(N__19360),
            .in3(N__23646),
            .lcout(buf_readRTD_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41141),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adress_i1_LC_3_9_0 .C_ON=1'b0;
    defparam \RTD.adress_i1_LC_3_9_0 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i1_LC_3_9_0 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \RTD.adress_i1_LC_3_9_0  (
            .in0(N__19344),
            .in1(N__19966),
            .in2(N__19651),
            .in3(N__19888),
            .lcout(adress_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41133),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adress_i2_LC_3_9_1 .C_ON=1'b0;
    defparam \RTD.adress_i2_LC_3_9_1 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i2_LC_3_9_1 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \RTD.adress_i2_LC_3_9_1  (
            .in0(N__19889),
            .in1(N__19345),
            .in2(N__19652),
            .in3(N__19335),
            .lcout(adress_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41133),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adress_i3_LC_3_9_2 .C_ON=1'b0;
    defparam \RTD.adress_i3_LC_3_9_2 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i3_LC_3_9_2 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \RTD.adress_i3_LC_3_9_2  (
            .in0(N__19336),
            .in1(N__19640),
            .in2(N__19327),
            .in3(N__19890),
            .lcout(adress_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41133),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adress_i4_LC_3_9_3 .C_ON=1'b0;
    defparam \RTD.adress_i4_LC_3_9_3 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i4_LC_3_9_3 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \RTD.adress_i4_LC_3_9_3  (
            .in0(N__19891),
            .in1(N__19314),
            .in2(N__19653),
            .in3(N__19326),
            .lcout(adress_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41133),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adress_i5_LC_3_9_4 .C_ON=1'b0;
    defparam \RTD.adress_i5_LC_3_9_4 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i5_LC_3_9_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \RTD.adress_i5_LC_3_9_4  (
            .in0(N__19315),
            .in1(N__19641),
            .in2(N__19303),
            .in3(N__19892),
            .lcout(adress_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41133),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adress_i6_LC_3_9_5 .C_ON=1'b0;
    defparam \RTD.adress_i6_LC_3_9_5 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i6_LC_3_9_5 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \RTD.adress_i6_LC_3_9_5  (
            .in0(N__19893),
            .in1(N__19992),
            .in2(N__19654),
            .in3(N__19302),
            .lcout(adress_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41133),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i10_LC_3_9_6 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i10_LC_3_9_6 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i10_LC_3_9_6 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \RTD.READ_DATA_i10_LC_3_9_6  (
            .in0(N__19290),
            .in1(N__19457),
            .in2(N__23391),
            .in3(N__22127),
            .lcout(buf_readRTD_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41133),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i12069_2_lut_LC_3_9_7 .C_ON=1'b0;
    defparam \RTD.i12069_2_lut_LC_3_9_7 .SEQ_MODE=4'b0000;
    defparam \RTD.i12069_2_lut_LC_3_9_7 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \RTD.i12069_2_lut_LC_3_9_7  (
            .in0(N__22260),
            .in1(N__22404),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n14465),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i8_LC_3_10_0 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i8_LC_3_10_0 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i8_LC_3_10_0 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \RTD.READ_DATA_i8_LC_3_10_0  (
            .in0(N__22123),
            .in1(N__21813),
            .in2(N__19474),
            .in3(N__19617),
            .lcout(buf_readRTD_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41129),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i2_LC_3_10_1 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i2_LC_3_10_1 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i2_LC_3_10_1 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \RTD.READ_DATA_i2_LC_3_10_1  (
            .in0(N__19506),
            .in1(N__19466),
            .in2(N__33261),
            .in3(N__22124),
            .lcout(buf_readRTD_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41129),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i4_LC_3_10_4 .C_ON=1'b0;
    defparam \RTD.read_buf_i4_LC_3_10_4 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i4_LC_3_10_4 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \RTD.read_buf_i4_LC_3_10_4  (
            .in0(N__19595),
            .in1(N__19579),
            .in2(N__19492),
            .in3(N__19750),
            .lcout(read_buf_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41129),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i4_LC_3_10_5 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i4_LC_3_10_5 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i4_LC_3_10_5 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \RTD.READ_DATA_i4_LC_3_10_5  (
            .in0(N__19596),
            .in1(N__19468),
            .in2(N__33207),
            .in3(N__22126),
            .lcout(buf_readRTD_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41129),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i3_LC_3_10_6 .C_ON=1'b0;
    defparam \RTD.read_buf_i3_LC_3_10_6 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i3_LC_3_10_6 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \RTD.read_buf_i3_LC_3_10_6  (
            .in0(N__19487),
            .in1(N__19578),
            .in2(N__19759),
            .in3(N__19507),
            .lcout(read_buf_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41129),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i3_LC_3_10_7 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i3_LC_3_10_7 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i3_LC_3_10_7 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \RTD.READ_DATA_i3_LC_3_10_7  (
            .in0(N__19491),
            .in1(N__19467),
            .in2(N__33558),
            .in3(N__22125),
            .lcout(buf_readRTD_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41129),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.bit_cnt_3771__i1_LC_5_5_1 .C_ON=1'b0;
    defparam \RTD.bit_cnt_3771__i1_LC_5_5_1 .SEQ_MODE=4'b1000;
    defparam \RTD.bit_cnt_3771__i1_LC_5_5_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \RTD.bit_cnt_3771__i1_LC_5_5_1  (
            .in0(_gnd_net_),
            .in1(N__20588),
            .in2(_gnd_net_),
            .in3(N__20615),
            .lcout(\RTD.bit_cnt_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41083),
            .ce(N__19396),
            .sr(N__19816));
    defparam \RTD.bit_cnt_3771__i0_LC_5_5_3 .C_ON=1'b0;
    defparam \RTD.bit_cnt_3771__i0_LC_5_5_3 .SEQ_MODE=4'b1000;
    defparam \RTD.bit_cnt_3771__i0_LC_5_5_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \RTD.bit_cnt_3771__i0_LC_5_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20587),
            .lcout(\RTD.bit_cnt_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41083),
            .ce(N__19396),
            .sr(N__19816));
    defparam \RTD.bit_cnt_3771__i2_LC_5_5_6 .C_ON=1'b0;
    defparam \RTD.bit_cnt_3771__i2_LC_5_5_6 .SEQ_MODE=4'b1000;
    defparam \RTD.bit_cnt_3771__i2_LC_5_5_6 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \RTD.bit_cnt_3771__i2_LC_5_5_6  (
            .in0(N__20616),
            .in1(_gnd_net_),
            .in2(N__20595),
            .in3(N__20562),
            .lcout(\RTD.bit_cnt_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41083),
            .ce(N__19396),
            .sr(N__19816));
    defparam \RTD.MOSI_59_LC_5_6_0 .C_ON=1'b0;
    defparam \RTD.MOSI_59_LC_5_6_0 .SEQ_MODE=4'b1000;
    defparam \RTD.MOSI_59_LC_5_6_0 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \RTD.MOSI_59_LC_5_6_0  (
            .in0(N__20927),
            .in1(N__19981),
            .in2(N__21004),
            .in3(N__22101),
            .lcout(RTD_SDI),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41142),
            .ce(N__19777),
            .sr(N__19953));
    defparam \RTD.i1_3_lut_4_lut_LC_5_6_3 .C_ON=1'b0;
    defparam \RTD.i1_3_lut_4_lut_LC_5_6_3 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_3_lut_4_lut_LC_5_6_3 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \RTD.i1_3_lut_4_lut_LC_5_6_3  (
            .in0(N__22220),
            .in1(N__20544),
            .in2(N__20524),
            .in3(N__20925),
            .lcout(\RTD.n33 ),
            .ltout(\RTD.n33_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i24_3_lut_4_lut_LC_5_6_4 .C_ON=1'b0;
    defparam \RTD.i24_3_lut_4_lut_LC_5_6_4 .SEQ_MODE=4'b0000;
    defparam \RTD.i24_3_lut_4_lut_LC_5_6_4 .LUT_INIT=16'b1111000001000100;
    LogicCell40 \RTD.i24_3_lut_4_lut_LC_5_6_4  (
            .in0(N__20926),
            .in1(N__22221),
            .in2(N__19762),
            .in3(N__22100),
            .lcout(\RTD.n11_adj_1394 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i2_3_lut_LC_5_6_6 .C_ON=1'b0;
    defparam \RTD.i2_3_lut_LC_5_6_6 .SEQ_MODE=4'b0000;
    defparam \RTD.i2_3_lut_LC_5_6_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \RTD.i2_3_lut_LC_5_6_6  (
            .in0(N__20923),
            .in1(N__22353),
            .in2(_gnd_net_),
            .in3(N__22099),
            .lcout(n1_adj_1575),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_2_lut_adj_20_LC_5_6_7 .C_ON=1'b0;
    defparam \RTD.i1_2_lut_adj_20_LC_5_6_7 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_2_lut_adj_20_LC_5_6_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \RTD.i1_2_lut_adj_20_LC_5_6_7  (
            .in0(_gnd_net_),
            .in1(N__22219),
            .in2(_gnd_net_),
            .in3(N__20924),
            .lcout(\RTD.n4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i31_3_lut_4_lut_3_lut_LC_5_7_0 .C_ON=1'b0;
    defparam \RTD.i31_3_lut_4_lut_3_lut_LC_5_7_0 .SEQ_MODE=4'b0000;
    defparam \RTD.i31_3_lut_4_lut_3_lut_LC_5_7_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \RTD.i31_3_lut_4_lut_3_lut_LC_5_7_0  (
            .in0(N__20894),
            .in1(N__22323),
            .in2(_gnd_net_),
            .in3(N__22191),
            .lcout(\RTD.n14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_2_lut_adj_24_LC_5_7_1 .C_ON=1'b0;
    defparam \RTD.i1_2_lut_adj_24_LC_5_7_1 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_2_lut_adj_24_LC_5_7_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \RTD.i1_2_lut_adj_24_LC_5_7_1  (
            .in0(_gnd_net_),
            .in1(N__19928),
            .in2(_gnd_net_),
            .in3(N__20144),
            .lcout(\RTD.n16614 ),
            .ltout(\RTD.n16614_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i2_3_lut_adj_19_LC_5_7_2 .C_ON=1'b0;
    defparam \RTD.i2_3_lut_adj_19_LC_5_7_2 .SEQ_MODE=4'b0000;
    defparam \RTD.i2_3_lut_adj_19_LC_5_7_2 .LUT_INIT=16'b1111111111110101;
    LogicCell40 \RTD.i2_3_lut_adj_19_LC_5_7_2  (
            .in0(N__20895),
            .in1(_gnd_net_),
            .in2(N__19657),
            .in3(N__21903),
            .lcout(\RTD.n11712 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_2_lut_adj_26_LC_5_7_3 .C_ON=1'b0;
    defparam \RTD.i1_2_lut_adj_26_LC_5_7_3 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_2_lut_adj_26_LC_5_7_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \RTD.i1_2_lut_adj_26_LC_5_7_3  (
            .in0(N__22324),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19859),
            .lcout(\RTD.n19855 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i19027_3_lut_LC_5_7_4 .C_ON=1'b0;
    defparam \RTD.i19027_3_lut_LC_5_7_4 .SEQ_MODE=4'b0000;
    defparam \RTD.i19027_3_lut_LC_5_7_4 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \RTD.i19027_3_lut_LC_5_7_4  (
            .in0(N__20896),
            .in1(N__20102),
            .in2(_gnd_net_),
            .in3(N__19843),
            .lcout(\RTD.n21091 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i16891_3_lut_LC_5_7_5 .C_ON=1'b0;
    defparam \RTD.i16891_3_lut_LC_5_7_5 .SEQ_MODE=4'b0000;
    defparam \RTD.i16891_3_lut_LC_5_7_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \RTD.i16891_3_lut_LC_5_7_5  (
            .in0(N__22192),
            .in1(N__20518),
            .in2(_gnd_net_),
            .in3(N__20540),
            .lcout(\RTD.n19482 ),
            .ltout(\RTD.n19482_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adc_state_3__I_0_66_Mux_0_i7_4_lut_LC_5_7_6 .C_ON=1'b0;
    defparam \RTD.adc_state_3__I_0_66_Mux_0_i7_4_lut_LC_5_7_6 .SEQ_MODE=4'b0000;
    defparam \RTD.adc_state_3__I_0_66_Mux_0_i7_4_lut_LC_5_7_6 .LUT_INIT=16'b0000010111010101;
    LogicCell40 \RTD.adc_state_3__I_0_66_Mux_0_i7_4_lut_LC_5_7_6  (
            .in0(N__20897),
            .in1(N__20103),
            .in2(N__19837),
            .in3(N__22030),
            .lcout(\RTD.n7_adj_1395 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_2_lut_3_lut_LC_5_7_7 .C_ON=1'b0;
    defparam \RTD.i1_2_lut_3_lut_LC_5_7_7 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_2_lut_3_lut_LC_5_7_7 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \RTD.i1_2_lut_3_lut_LC_5_7_7  (
            .in0(N__22190),
            .in1(N__21983),
            .in2(_gnd_net_),
            .in3(N__20893),
            .lcout(\RTD.n1_adj_1393 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i18129_2_lut_LC_5_8_0 .C_ON=1'b0;
    defparam \RTD.i18129_2_lut_LC_5_8_0 .SEQ_MODE=4'b0000;
    defparam \RTD.i18129_2_lut_LC_5_8_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \RTD.i18129_2_lut_LC_5_8_0  (
            .in0(_gnd_net_),
            .in1(N__22193),
            .in2(_gnd_net_),
            .in3(N__21989),
            .lcout(\RTD.n7285 ),
            .ltout(\RTD.n7285_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_4_lut_adj_13_LC_5_8_1 .C_ON=1'b0;
    defparam \RTD.i1_4_lut_adj_13_LC_5_8_1 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_4_lut_adj_13_LC_5_8_1 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \RTD.i1_4_lut_adj_13_LC_5_8_1  (
            .in0(N__20914),
            .in1(N__19929),
            .in2(N__19834),
            .in3(N__20142),
            .lcout(),
            .ltout(\RTD.n21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_4_lut_adj_14_LC_5_8_2 .C_ON=1'b0;
    defparam \RTD.i1_4_lut_adj_14_LC_5_8_2 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_4_lut_adj_14_LC_5_8_2 .LUT_INIT=16'b0100000011001000;
    LogicCell40 \RTD.i1_4_lut_adj_14_LC_5_8_2  (
            .in0(N__22350),
            .in1(N__20098),
            .in2(N__19831),
            .in3(N__21990),
            .lcout(\RTD.n16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i18734_4_lut_LC_5_8_3 .C_ON=1'b0;
    defparam \RTD.i18734_4_lut_LC_5_8_3 .SEQ_MODE=4'b0000;
    defparam \RTD.i18734_4_lut_LC_5_8_3 .LUT_INIT=16'b1010101010101000;
    LogicCell40 \RTD.i18734_4_lut_LC_5_8_3  (
            .in0(N__19828),
            .in1(N__22351),
            .in2(N__20104),
            .in3(N__20005),
            .lcout(),
            .ltout(\RTD.n20969_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adc_state_i2_LC_5_8_4 .C_ON=1'b0;
    defparam \RTD.adc_state_i2_LC_5_8_4 .SEQ_MODE=4'b1000;
    defparam \RTD.adc_state_i2_LC_5_8_4 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \RTD.adc_state_i2_LC_5_8_4  (
            .in0(N__22352),
            .in1(N__20475),
            .in2(N__19819),
            .in3(N__21991),
            .lcout(adc_state_2_adj_1474),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41134),
            .ce(N__20683),
            .sr(_gnd_net_));
    defparam \RTD.i1_2_lut_LC_5_8_5 .C_ON=1'b0;
    defparam \RTD.i1_2_lut_LC_5_8_5 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_2_lut_LC_5_8_5 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \RTD.i1_2_lut_LC_5_8_5  (
            .in0(N__20519),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20545),
            .lcout(\RTD.n32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i4916_2_lut_LC_5_8_6 .C_ON=1'b0;
    defparam \RTD.i4916_2_lut_LC_5_8_6 .SEQ_MODE=4'b0000;
    defparam \RTD.i4916_2_lut_LC_5_8_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \RTD.i4916_2_lut_LC_5_8_6  (
            .in0(_gnd_net_),
            .in1(N__22194),
            .in2(_gnd_net_),
            .in3(N__20913),
            .lcout(\RTD.n1_adj_1392 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adress_i7_LC_5_9_0 .C_ON=1'b0;
    defparam \RTD.adress_i7_LC_5_9_0 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i7_LC_5_9_0 .LUT_INIT=16'b1100101011000000;
    LogicCell40 \RTD.adress_i7_LC_5_9_0  (
            .in0(N__20143),
            .in1(N__19999),
            .in2(N__22261),
            .in3(N__20944),
            .lcout(\RTD.adress_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41082),
            .ce(N__19894),
            .sr(N__19957));
    defparam \RTD.adress_i0_LC_5_9_1 .C_ON=1'b0;
    defparam \RTD.adress_i0_LC_5_9_1 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i0_LC_5_9_1 .LUT_INIT=16'b1100110001011111;
    LogicCell40 \RTD.adress_i0_LC_5_9_1  (
            .in0(N__20943),
            .in1(N__19980),
            .in2(N__20149),
            .in3(N__22248),
            .lcout(adress_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41082),
            .ce(N__19894),
            .sr(N__19957));
    defparam \RTD.i7_4_lut_LC_5_9_2 .C_ON=1'b0;
    defparam \RTD.i7_4_lut_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \RTD.i7_4_lut_LC_5_9_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \RTD.i7_4_lut_LC_5_9_2  (
            .in0(N__20077),
            .in1(N__21202),
            .in2(N__20044),
            .in3(N__20797),
            .lcout(\RTD.adress_7_N_1331_7 ),
            .ltout(\RTD.adress_7_N_1331_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_2_lut_adj_16_LC_5_9_3 .C_ON=1'b0;
    defparam \RTD.i1_2_lut_adj_16_LC_5_9_3 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_2_lut_adj_16_LC_5_9_3 .LUT_INIT=16'b1111010111110101;
    LogicCell40 \RTD.i1_2_lut_adj_16_LC_5_9_3  (
            .in0(N__20941),
            .in1(_gnd_net_),
            .in2(N__19936),
            .in3(_gnd_net_),
            .lcout(\RTD.n11 ),
            .ltout(\RTD.n11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i34_4_lut_LC_5_9_4 .C_ON=1'b0;
    defparam \RTD.i34_4_lut_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \RTD.i34_4_lut_LC_5_9_4 .LUT_INIT=16'b1111101101010001;
    LogicCell40 \RTD.i34_4_lut_LC_5_9_4  (
            .in0(N__22247),
            .in1(N__19933),
            .in2(N__19900),
            .in3(N__20942),
            .lcout(),
            .ltout(\RTD.n19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i35_4_lut_LC_5_9_5 .C_ON=1'b0;
    defparam \RTD.i35_4_lut_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \RTD.i35_4_lut_LC_5_9_5 .LUT_INIT=16'b1000100011011000;
    LogicCell40 \RTD.i35_4_lut_LC_5_9_5  (
            .in0(N__22361),
            .in1(N__19863),
            .in2(N__19897),
            .in3(N__22026),
            .lcout(n13151),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i22_4_lut_LC_5_9_6 .C_ON=1'b0;
    defparam \RTD.i22_4_lut_LC_5_9_6 .SEQ_MODE=4'b0000;
    defparam \RTD.i22_4_lut_LC_5_9_6 .LUT_INIT=16'b1101000111000000;
    LogicCell40 \RTD.i22_4_lut_LC_5_9_6  (
            .in0(N__20730),
            .in1(N__22360),
            .in2(N__19864),
            .in3(N__20790),
            .lcout(n13162),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.mode_53_LC_5_10_0 .C_ON=1'b0;
    defparam \RTD.mode_53_LC_5_10_0 .SEQ_MODE=4'b1000;
    defparam \RTD.mode_53_LC_5_10_0 .LUT_INIT=16'b1111111100001000;
    LogicCell40 \RTD.mode_53_LC_5_10_0  (
            .in0(N__20965),
            .in1(N__20145),
            .in2(N__21910),
            .in3(N__20113),
            .lcout(\RTD.mode ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41116),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i2_4_lut_LC_5_10_1 .C_ON=1'b0;
    defparam \RTD.i2_4_lut_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \RTD.i2_4_lut_LC_5_10_1 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \RTD.i2_4_lut_LC_5_10_1  (
            .in0(N__23819),
            .in1(N__20061),
            .in2(N__42075),
            .in3(N__20070),
            .lcout(\RTD.n10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i2_LC_5_10_2 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i2_LC_5_10_2 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i2_LC_5_10_2 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \RTD.cfg_buf_i2_LC_5_10_2  (
            .in0(N__20071),
            .in1(N__21155),
            .in2(N__23823),
            .in3(N__21184),
            .lcout(\RTD.cfg_buf_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41116),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i4_LC_5_10_3 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i4_LC_5_10_3 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i4_LC_5_10_3 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \RTD.cfg_buf_i4_LC_5_10_3  (
            .in0(N__21185),
            .in1(N__20062),
            .in2(N__42074),
            .in3(N__21157),
            .lcout(\RTD.cfg_buf_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41116),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i7_LC_5_10_4 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i7_LC_5_10_4 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i7_LC_5_10_4 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \RTD.cfg_buf_i7_LC_5_10_4  (
            .in0(N__20053),
            .in1(N__21156),
            .in2(N__24194),
            .in3(N__21187),
            .lcout(\RTD.cfg_buf_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41116),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i4_4_lut_LC_5_10_5 .C_ON=1'b0;
    defparam \RTD.i4_4_lut_LC_5_10_5 .SEQ_MODE=4'b0000;
    defparam \RTD.i4_4_lut_LC_5_10_5 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \RTD.i4_4_lut_LC_5_10_5  (
            .in0(N__23697),
            .in1(N__20052),
            .in2(N__24195),
            .in3(N__20034),
            .lcout(\RTD.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i1_LC_5_10_6 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i1_LC_5_10_6 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i1_LC_5_10_6 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \RTD.cfg_buf_i1_LC_5_10_6  (
            .in0(N__20035),
            .in1(N__21154),
            .in2(N__23698),
            .in3(N__21183),
            .lcout(cfg_buf_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41116),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i5_LC_5_10_7 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i5_LC_5_10_7 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i5_LC_5_10_7 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \RTD.cfg_buf_i5_LC_5_10_7  (
            .in0(N__21186),
            .in1(N__21214),
            .in2(N__41436),
            .in3(N__21158),
            .lcout(\RTD.cfg_buf_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41116),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_7_i19_3_lut_LC_5_11_0.C_ON=1'b0;
    defparam mux_129_Mux_7_i19_3_lut_LC_5_11_0.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_7_i19_3_lut_LC_5_11_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_129_Mux_7_i19_3_lut_LC_5_11_0 (
            .in0(N__23581),
            .in1(N__20189),
            .in2(_gnd_net_),
            .in3(N__56901),
            .lcout(),
            .ltout(n19_adj_1622_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19365_LC_5_11_1.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19365_LC_5_11_1.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19365_LC_5_11_1.LUT_INIT=16'b1011100011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_19365_LC_5_11_1 (
            .in0(N__20026),
            .in1(N__57503),
            .in2(N__20200),
            .in3(N__47737),
            .lcout(n21961),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i15_LC_5_11_2 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i15_LC_5_11_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i15_LC_5_11_2 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \ADC_VAC.ADC_DATA_i15_LC_5_11_2  (
            .in0(N__48315),
            .in1(N__20190),
            .in2(N__48533),
            .in3(N__21238),
            .lcout(buf_adcdata_vac_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55174),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_3_i30_3_lut_LC_5_11_3.C_ON=1'b0;
    defparam mux_130_Mux_3_i30_3_lut_LC_5_11_3.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_3_i30_3_lut_LC_5_11_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_130_Mux_3_i30_3_lut_LC_5_11_3 (
            .in0(N__20176),
            .in1(N__21022),
            .in2(_gnd_net_),
            .in3(N__56347),
            .lcout(n30_adj_1612),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i3_LC_5_11_5 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i3_LC_5_11_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i3_LC_5_11_5 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i3_LC_5_11_5  (
            .in0(N__50908),
            .in1(N__48999),
            .in2(N__49041),
            .in3(N__21042),
            .lcout(buf_adcdata_iac_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55174),
            .ce(),
            .sr(_gnd_net_));
    defparam i18784_2_lut_LC_5_11_6.C_ON=1'b0;
    defparam i18784_2_lut_LC_5_11_6.SEQ_MODE=4'b0000;
    defparam i18784_2_lut_LC_5_11_6.LUT_INIT=16'b0000000011001100;
    LogicCell40 i18784_2_lut_LC_5_11_6 (
            .in0(_gnd_net_),
            .in1(N__20164),
            .in2(_gnd_net_),
            .in3(N__56902),
            .lcout(n20937),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i2_LC_5_11_7 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i2_LC_5_11_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i2_LC_5_11_7 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i2_LC_5_11_7  (
            .in0(N__50907),
            .in1(N__48998),
            .in2(N__21322),
            .in3(N__22490),
            .lcout(buf_adcdata_iac_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55174),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i18_LC_5_12_0 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i18_LC_5_12_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i18_LC_5_12_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i18_LC_5_12_0  (
            .in0(N__48505),
            .in1(N__48321),
            .in2(N__21298),
            .in3(N__23852),
            .lcout(buf_adcdata_vac_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55190),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i21_LC_5_12_2 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i21_LC_5_12_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i21_LC_5_12_2 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i21_LC_5_12_2  (
            .in0(N__48506),
            .in1(N__48322),
            .in2(N__21346),
            .in3(N__21839),
            .lcout(buf_adcdata_vac_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55190),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i9_LC_5_12_3 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i9_LC_5_12_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i9_LC_5_12_3 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i9_LC_5_12_3  (
            .in0(N__21251),
            .in1(N__50935),
            .in2(N__21447),
            .in3(N__50516),
            .lcout(cmd_rdadctmp_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55190),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i11_LC_5_12_5 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i11_LC_5_12_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i11_LC_5_12_5 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i11_LC_5_12_5  (
            .in0(N__49025),
            .in1(N__50934),
            .in2(N__21321),
            .in3(N__50515),
            .lcout(cmd_rdadctmp_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55190),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19423_LC_5_13_0.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19423_LC_5_13_0.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19423_LC_5_13_0.LUT_INIT=16'b1101101010001010;
    LogicCell40 comm_cmd_0__bdd_4_lut_19423_LC_5_13_0 (
            .in0(N__56904),
            .in1(N__24690),
            .in2(N__57538),
            .in3(N__27873),
            .lcout(n22039),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i29_LC_5_13_1 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i29_LC_5_13_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i29_LC_5_13_1 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i29_LC_5_13_1  (
            .in0(N__37878),
            .in1(N__21338),
            .in2(N__20305),
            .in3(N__48286),
            .lcout(cmd_rdadctmp_29_adj_1414),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55204),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i28_LC_5_13_4 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i28_LC_5_13_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i28_LC_5_13_4 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i28_LC_5_13_4  (
            .in0(N__48285),
            .in1(N__20300),
            .in2(N__21276),
            .in3(N__37877),
            .lcout(cmd_rdadctmp_28_adj_1415),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55204),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i20_LC_5_13_6 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i20_LC_5_13_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i20_LC_5_13_6 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC.ADC_DATA_i20_LC_5_13_6  (
            .in0(N__48284),
            .in1(N__48492),
            .in2(N__25706),
            .in3(N__20304),
            .lcout(buf_adcdata_vac_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55204),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i7_LC_5_14_0 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i7_LC_5_14_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i7_LC_5_14_0 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i7_LC_5_14_0  (
            .in0(N__22818),
            .in1(N__48287),
            .in2(N__21583),
            .in3(N__37872),
            .lcout(cmd_rdadctmp_7_adj_1436),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55216),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19516_LC_5_14_5.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19516_LC_5_14_5.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19516_LC_5_14_5.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_19516_LC_5_14_5 (
            .in0(N__21403),
            .in1(N__57446),
            .in2(N__20290),
            .in3(N__47823),
            .lcout(n22117),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_199_LC_5_15_1.C_ON=1'b0;
    defparam i1_4_lut_adj_199_LC_5_15_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_199_LC_5_15_1.LUT_INIT=16'b0000111100000110;
    LogicCell40 i1_4_lut_adj_199_LC_5_15_1 (
            .in0(N__48203),
            .in1(N__29855),
            .in2(N__20244),
            .in3(N__29782),
            .lcout(n14_adj_1577),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_104_LC_5_15_5.C_ON=1'b0;
    defparam i1_2_lut_adj_104_LC_5_15_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_104_LC_5_15_5.LUT_INIT=16'b0011001100000000;
    LogicCell40 i1_2_lut_adj_104_LC_5_15_5 (
            .in0(_gnd_net_),
            .in1(N__29854),
            .in2(_gnd_net_),
            .in3(N__29781),
            .lcout(n20573),
            .ltout(n20573_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.CS_37_LC_5_15_6 .C_ON=1'b0;
    defparam \ADC_VAC.CS_37_LC_5_15_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.CS_37_LC_5_15_6 .LUT_INIT=16'b0011001100100011;
    LogicCell40 \ADC_VAC.CS_37_LC_5_15_6  (
            .in0(N__22982),
            .in1(N__20263),
            .in2(N__20257),
            .in3(N__48205),
            .lcout(VAC_CS),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55227),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.SCLK_35_LC_5_15_7 .C_ON=1'b0;
    defparam \ADC_VAC.SCLK_35_LC_5_15_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.SCLK_35_LC_5_15_7 .LUT_INIT=16'b1101000011100100;
    LogicCell40 \ADC_VAC.SCLK_35_LC_5_15_7  (
            .in0(N__48204),
            .in1(N__29856),
            .in2(N__20217),
            .in3(N__29783),
            .lcout(VAC_SCLK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55227),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i12_LC_5_16_1 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i12_LC_5_16_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i12_LC_5_16_1 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i12_LC_5_16_1  (
            .in0(N__48961),
            .in1(N__50954),
            .in2(N__21801),
            .in3(N__33462),
            .lcout(buf_adcdata_iac_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55237),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i22_LC_5_16_4 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i22_LC_5_16_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i22_LC_5_16_4 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i22_LC_5_16_4  (
            .in0(N__50493),
            .in1(N__21777),
            .in2(N__50965),
            .in3(N__24446),
            .lcout(cmd_rdadctmp_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55237),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i20_LC_5_16_5 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i20_LC_5_16_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i20_LC_5_16_5 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i20_LC_5_16_5  (
            .in0(N__21794),
            .in1(N__50956),
            .in2(N__21759),
            .in3(N__50494),
            .lcout(cmd_rdadctmp_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55237),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i14_LC_5_16_7 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i14_LC_5_16_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i14_LC_5_16_7 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i14_LC_5_16_7  (
            .in0(N__48962),
            .in1(N__50955),
            .in2(N__24453),
            .in3(N__29576),
            .lcout(buf_adcdata_iac_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55237),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i13_LC_5_17_2 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i13_LC_5_17_2 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i13_LC_5_17_2 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i13_LC_5_17_2  (
            .in0(N__50880),
            .in1(N__48967),
            .in2(N__21781),
            .in3(N__25808),
            .lcout(buf_adcdata_iac_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55240),
            .ce(),
            .sr(_gnd_net_));
    defparam i18773_2_lut_LC_5_17_5.C_ON=1'b0;
    defparam i18773_2_lut_LC_5_17_5.SEQ_MODE=4'b0000;
    defparam i18773_2_lut_LC_5_17_5.LUT_INIT=16'b0101010100000000;
    LogicCell40 i18773_2_lut_LC_5_17_5 (
            .in0(N__56911),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20407),
            .lcout(n21001),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i11_LC_5_17_7 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i11_LC_5_17_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i11_LC_5_17_7 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i11_LC_5_17_7  (
            .in0(N__48966),
            .in1(N__50881),
            .in2(N__21760),
            .in3(N__33534),
            .lcout(buf_adcdata_iac_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55240),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_354_Mux_7_i15_4_lut_LC_5_19_5.C_ON=1'b0;
    defparam comm_state_3__I_0_354_Mux_7_i15_4_lut_LC_5_19_5.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_354_Mux_7_i15_4_lut_LC_5_19_5.LUT_INIT=16'b0101110100001000;
    LogicCell40 comm_state_3__I_0_354_Mux_7_i15_4_lut_LC_5_19_5 (
            .in0(N__54723),
            .in1(N__30079),
            .in2(N__52192),
            .in3(N__42435),
            .lcout(data_index_9_N_212_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.bit_cnt_i3_LC_6_4_0 .C_ON=1'b0;
    defparam \CLK_DDS.bit_cnt_i3_LC_6_4_0 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.bit_cnt_i3_LC_6_4_0 .LUT_INIT=16'b0111100011110000;
    LogicCell40 \CLK_DDS.bit_cnt_i3_LC_6_4_0  (
            .in0(N__20430),
            .in1(N__23232),
            .in2(N__23209),
            .in3(N__20453),
            .lcout(bit_cnt_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55082),
            .ce(N__28907),
            .sr(N__20740));
    defparam \CLK_DDS.bit_cnt_i2_LC_6_4_1 .C_ON=1'b0;
    defparam \CLK_DDS.bit_cnt_i2_LC_6_4_1 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.bit_cnt_i2_LC_6_4_1 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \CLK_DDS.bit_cnt_i2_LC_6_4_1  (
            .in0(N__23231),
            .in1(_gnd_net_),
            .in2(N__20457),
            .in3(N__20429),
            .lcout(bit_cnt_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55082),
            .ce(N__28907),
            .sr(N__20740));
    defparam \CLK_DDS.bit_cnt_i1_LC_6_4_2 .C_ON=1'b0;
    defparam \CLK_DDS.bit_cnt_i1_LC_6_4_2 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.bit_cnt_i1_LC_6_4_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \CLK_DDS.bit_cnt_i1_LC_6_4_2  (
            .in0(_gnd_net_),
            .in1(N__20449),
            .in2(_gnd_net_),
            .in3(N__23230),
            .lcout(bit_cnt_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55082),
            .ce(N__28907),
            .sr(N__20740));
    defparam \CLK_DDS.dds_state_i0_LC_6_5_0 .C_ON=1'b0;
    defparam \CLK_DDS.dds_state_i0_LC_6_5_0 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.dds_state_i0_LC_6_5_0 .LUT_INIT=16'b1100010100000101;
    LogicCell40 \CLK_DDS.dds_state_i0_LC_6_5_0  (
            .in0(N__28612),
            .in1(N__20413),
            .in2(N__28908),
            .in3(N__23191),
            .lcout(dds_state_0_adj_1447),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55087),
            .ce(N__20640),
            .sr(_gnd_net_));
    defparam \CLK_DDS.i19109_4_lut_LC_6_6_0 .C_ON=1'b0;
    defparam \CLK_DDS.i19109_4_lut_LC_6_6_0 .SEQ_MODE=4'b0000;
    defparam \CLK_DDS.i19109_4_lut_LC_6_6_0 .LUT_INIT=16'b1111111111011110;
    LogicCell40 \CLK_DDS.i19109_4_lut_LC_6_6_0  (
            .in0(N__28593),
            .in1(N__28865),
            .in2(N__28678),
            .in3(N__28746),
            .lcout(\CLK_DDS.n9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.dds_state_i1_LC_6_6_1 .C_ON=1'b0;
    defparam \CLK_DDS.dds_state_i1_LC_6_6_1 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.dds_state_i1_LC_6_6_1 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \CLK_DDS.dds_state_i1_LC_6_6_1  (
            .in0(N__28749),
            .in1(N__28594),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(dds_state_1_adj_1446),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55095),
            .ce(N__20641),
            .sr(N__28973));
    defparam \RTD.i2_3_lut_adj_18_LC_6_6_2 .C_ON=1'b0;
    defparam \RTD.i2_3_lut_adj_18_LC_6_6_2 .SEQ_MODE=4'b0000;
    defparam \RTD.i2_3_lut_adj_18_LC_6_6_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \RTD.i2_3_lut_adj_18_LC_6_6_2  (
            .in0(N__20614),
            .in1(N__20586),
            .in2(_gnd_net_),
            .in3(N__20561),
            .lcout(\RTD.n17638 ),
            .ltout(\RTD.n17638_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i19033_3_lut_LC_6_6_3 .C_ON=1'b0;
    defparam \RTD.i19033_3_lut_LC_6_6_3 .SEQ_MODE=4'b0000;
    defparam \RTD.i19033_3_lut_LC_6_6_3 .LUT_INIT=16'b1111111100111111;
    LogicCell40 \RTD.i19033_3_lut_LC_6_6_3  (
            .in0(_gnd_net_),
            .in1(N__20520),
            .in2(N__20482),
            .in3(N__22222),
            .lcout(),
            .ltout(\RTD.n21063_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adc_state_3__I_0_66_Mux_0_i14_4_lut_LC_6_6_4 .C_ON=1'b0;
    defparam \RTD.adc_state_3__I_0_66_Mux_0_i14_4_lut_LC_6_6_4 .SEQ_MODE=4'b0000;
    defparam \RTD.adc_state_3__I_0_66_Mux_0_i14_4_lut_LC_6_6_4 .LUT_INIT=16'b1011100010001000;
    LogicCell40 \RTD.adc_state_3__I_0_66_Mux_0_i14_4_lut_LC_6_6_4  (
            .in0(N__20479),
            .in1(N__22102),
            .in2(N__20461),
            .in3(N__20928),
            .lcout(\RTD.n17676 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.i3_3_lut_4_lut_LC_6_6_5 .C_ON=1'b0;
    defparam \CLK_DDS.i3_3_lut_4_lut_LC_6_6_5 .SEQ_MODE=4'b0000;
    defparam \CLK_DDS.i3_3_lut_4_lut_LC_6_6_5 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \CLK_DDS.i3_3_lut_4_lut_LC_6_6_5  (
            .in0(N__28748),
            .in1(N__28591),
            .in2(N__20458),
            .in3(N__20431),
            .lcout(n8_adj_1409),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.i1_3_lut_LC_6_6_6 .C_ON=1'b0;
    defparam \CLK_DDS.i1_3_lut_LC_6_6_6 .SEQ_MODE=4'b0000;
    defparam \CLK_DDS.i1_3_lut_LC_6_6_6 .LUT_INIT=16'b1100110001000100;
    LogicCell40 \CLK_DDS.i1_3_lut_LC_6_6_6  (
            .in0(N__28592),
            .in1(N__28866),
            .in2(_gnd_net_),
            .in3(N__28747),
            .lcout(\CLK_DDS.n16711 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adc_state_i1_LC_6_7_3 .C_ON=1'b0;
    defparam \RTD.adc_state_i1_LC_6_7_3 .SEQ_MODE=4'b1000;
    defparam \RTD.adc_state_i1_LC_6_7_3 .LUT_INIT=16'b0111001101010000;
    LogicCell40 \RTD.adc_state_i1_LC_6_7_3  (
            .in0(N__22387),
            .in1(N__20731),
            .in2(N__20719),
            .in3(N__20940),
            .lcout(\RTD.adc_state_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41099),
            .ce(N__20679),
            .sr(_gnd_net_));
    defparam \RTD.adc_state_i3_LC_6_7_4 .C_ON=1'b0;
    defparam \RTD.adc_state_i3_LC_6_7_4 .SEQ_MODE=4'b1000;
    defparam \RTD.adc_state_i3_LC_6_7_4 .LUT_INIT=16'b0000010110111011;
    LogicCell40 \RTD.adc_state_i3_LC_6_7_4  (
            .in0(N__22354),
            .in1(N__20710),
            .in2(N__20704),
            .in3(N__22104),
            .lcout(\RTD.adc_state_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41099),
            .ce(N__20679),
            .sr(_gnd_net_));
    defparam \RTD.adc_state_i0_LC_6_7_5 .C_ON=1'b0;
    defparam \RTD.adc_state_i0_LC_6_7_5 .SEQ_MODE=4'b1000;
    defparam \RTD.adc_state_i0_LC_6_7_5 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \RTD.adc_state_i0_LC_6_7_5  (
            .in0(N__22388),
            .in1(N__20695),
            .in2(_gnd_net_),
            .in3(N__20689),
            .lcout(\RTD.adc_state_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41099),
            .ce(N__20679),
            .sr(_gnd_net_));
    defparam \RTD.cfg_tmp_i1_LC_6_8_0 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i1_LC_6_8_0 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i1_LC_6_8_0 .LUT_INIT=16'b1100101011000000;
    LogicCell40 \RTD.cfg_tmp_i1_LC_6_8_0  (
            .in0(N__20932),
            .in1(N__20983),
            .in2(N__22130),
            .in3(N__23682),
            .lcout(\RTD.cfg_tmp_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41098),
            .ce(N__20767),
            .sr(N__20752));
    defparam \RTD.cfg_tmp_i2_LC_6_8_1 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i2_LC_6_8_1 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i2_LC_6_8_1 .LUT_INIT=16'b1110010010100000;
    LogicCell40 \RTD.cfg_tmp_i2_LC_6_8_1  (
            .in0(N__22032),
            .in1(N__23827),
            .in2(N__20668),
            .in3(N__20937),
            .lcout(\RTD.cfg_tmp_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41098),
            .ce(N__20767),
            .sr(N__20752));
    defparam \RTD.cfg_tmp_i3_LC_6_8_2 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i3_LC_6_8_2 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i3_LC_6_8_2 .LUT_INIT=16'b1100110010100000;
    LogicCell40 \RTD.cfg_tmp_i3_LC_6_8_2  (
            .in0(N__20933),
            .in1(N__20659),
            .in2(N__23785),
            .in3(N__22036),
            .lcout(\RTD.cfg_tmp_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41098),
            .ce(N__20767),
            .sr(N__20752));
    defparam \RTD.cfg_tmp_i4_LC_6_8_3 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i4_LC_6_8_3 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i4_LC_6_8_3 .LUT_INIT=16'b1101100010001000;
    LogicCell40 \RTD.cfg_tmp_i4_LC_6_8_3  (
            .in0(N__22033),
            .in1(N__20653),
            .in2(N__42076),
            .in3(N__20938),
            .lcout(\RTD.cfg_tmp_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41098),
            .ce(N__20767),
            .sr(N__20752));
    defparam \RTD.cfg_tmp_i5_LC_6_8_4 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i5_LC_6_8_4 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i5_LC_6_8_4 .LUT_INIT=16'b1110110000100000;
    LogicCell40 \RTD.cfg_tmp_i5_LC_6_8_4  (
            .in0(N__20934),
            .in1(N__22035),
            .in2(N__41437),
            .in3(N__20647),
            .lcout(\RTD.cfg_tmp_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41098),
            .ce(N__20767),
            .sr(N__20752));
    defparam \RTD.cfg_tmp_i6_LC_6_8_5 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i6_LC_6_8_5 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i6_LC_6_8_5 .LUT_INIT=16'b1101100010001000;
    LogicCell40 \RTD.cfg_tmp_i6_LC_6_8_5  (
            .in0(N__22034),
            .in1(N__21016),
            .in2(N__29329),
            .in3(N__20939),
            .lcout(\RTD.cfg_tmp_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41098),
            .ce(N__20767),
            .sr(N__20752));
    defparam \RTD.cfg_tmp_i7_LC_6_8_6 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i7_LC_6_8_6 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i7_LC_6_8_6 .LUT_INIT=16'b1100110010100000;
    LogicCell40 \RTD.cfg_tmp_i7_LC_6_8_6  (
            .in0(N__20935),
            .in1(N__21010),
            .in2(N__24199),
            .in3(N__22037),
            .lcout(\RTD.cfg_tmp_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41098),
            .ce(N__20767),
            .sr(N__20752));
    defparam \RTD.cfg_tmp_i0_LC_6_8_7 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i0_LC_6_8_7 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i0_LC_6_8_7 .LUT_INIT=16'b1101100010001000;
    LogicCell40 \RTD.cfg_tmp_i0_LC_6_8_7  (
            .in0(N__22031),
            .in1(N__20994),
            .in2(N__23737),
            .in3(N__20936),
            .lcout(\RTD.cfg_tmp_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41098),
            .ce(N__20767),
            .sr(N__20752));
    defparam \RTD.i1_3_lut_LC_6_9_2 .C_ON=1'b0;
    defparam \RTD.i1_3_lut_LC_6_9_2 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_3_lut_LC_6_9_2 .LUT_INIT=16'b0000101011111111;
    LogicCell40 \RTD.i1_3_lut_LC_6_9_2  (
            .in0(N__20945),
            .in1(_gnd_net_),
            .in2(N__22389),
            .in3(N__21152),
            .lcout(n18586),
            .ltout(n18586_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i0_LC_6_9_3 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i0_LC_6_9_3 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i0_LC_6_9_3 .LUT_INIT=16'b1100000010100000;
    LogicCell40 \RTD.cfg_buf_i0_LC_6_9_3  (
            .in0(N__20806),
            .in1(N__23732),
            .in2(N__20809),
            .in3(N__21153),
            .lcout(cfg_buf_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41079),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_4_lut_adj_23_LC_6_9_4 .C_ON=1'b0;
    defparam \RTD.i1_4_lut_adj_23_LC_6_9_4 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_4_lut_adj_23_LC_6_9_4 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \RTD.i1_4_lut_adj_23_LC_6_9_4  (
            .in0(N__23733),
            .in1(N__21114),
            .in2(N__29325),
            .in3(N__20805),
            .lcout(\RTD.n9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i18127_2_lut_LC_6_9_5 .C_ON=1'b0;
    defparam \RTD.i18127_2_lut_LC_6_9_5 .SEQ_MODE=4'b0000;
    defparam \RTD.i18127_2_lut_LC_6_9_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \RTD.i18127_2_lut_LC_6_9_5  (
            .in0(N__22223),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22355),
            .lcout(),
            .ltout(\RTD.n20722_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i30_4_lut_LC_6_9_6 .C_ON=1'b0;
    defparam \RTD.i30_4_lut_LC_6_9_6 .SEQ_MODE=4'b0000;
    defparam \RTD.i30_4_lut_LC_6_9_6 .LUT_INIT=16'b1100110000001010;
    LogicCell40 \RTD.i30_4_lut_LC_6_9_6  (
            .in0(N__20791),
            .in1(N__20779),
            .in2(N__20770),
            .in3(N__22025),
            .lcout(\RTD.n13198 ),
            .ltout(\RTD.n13198_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i12587_2_lut_LC_6_9_7 .C_ON=1'b0;
    defparam \RTD.i12587_2_lut_LC_6_9_7 .SEQ_MODE=4'b0000;
    defparam \RTD.i12587_2_lut_LC_6_9_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \RTD.i12587_2_lut_LC_6_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20755),
            .in3(N__22359),
            .lcout(\RTD.n14984 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i3_4_lut_LC_6_10_0 .C_ON=1'b0;
    defparam \RTD.i3_4_lut_LC_6_10_0 .SEQ_MODE=4'b0000;
    defparam \RTD.i3_4_lut_LC_6_10_0 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \RTD.i3_4_lut_LC_6_10_0  (
            .in0(N__41426),
            .in1(N__21213),
            .in2(N__23777),
            .in3(N__21195),
            .lcout(\RTD.n11_adj_1396 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i3_LC_6_10_1 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i3_LC_6_10_1 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i3_LC_6_10_1 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \RTD.cfg_buf_i3_LC_6_10_1  (
            .in0(N__21196),
            .in1(N__21159),
            .in2(N__23778),
            .in3(N__21181),
            .lcout(\RTD.cfg_buf_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41097),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i6_LC_6_10_2 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i6_LC_6_10_2 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i6_LC_6_10_2 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \RTD.cfg_buf_i6_LC_6_10_2  (
            .in0(N__21182),
            .in1(N__21115),
            .in2(N__29318),
            .in3(N__21160),
            .lcout(\RTD.cfg_buf_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__41097),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19496_LC_6_10_4.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19496_LC_6_10_4.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19496_LC_6_10_4.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_0__bdd_4_lut_19496_LC_6_10_4 (
            .in0(N__23767),
            .in1(N__57310),
            .in2(N__21103),
            .in3(N__56903),
            .lcout(),
            .ltout(n22099_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22099_bdd_4_lut_LC_6_10_5.C_ON=1'b0;
    defparam n22099_bdd_4_lut_LC_6_10_5.SEQ_MODE=4'b0000;
    defparam n22099_bdd_4_lut_LC_6_10_5.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22099_bdd_4_lut_LC_6_10_5 (
            .in0(N__57311),
            .in1(N__21065),
            .in2(N__21079),
            .in3(N__23290),
            .lcout(),
            .ltout(n22102_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18255_3_lut_LC_6_10_6.C_ON=1'b0;
    defparam i18255_3_lut_LC_6_10_6.SEQ_MODE=4'b0000;
    defparam i18255_3_lut_LC_6_10_6.LUT_INIT=16'b1110010011100100;
    LogicCell40 i18255_3_lut_LC_6_10_6 (
            .in0(N__47820),
            .in1(N__29524),
            .in2(N__21076),
            .in3(_gnd_net_),
            .lcout(n20850),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i19_LC_6_11_0 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i19_LC_6_11_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i19_LC_6_11_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i19_LC_6_11_0  (
            .in0(N__48319),
            .in1(N__48495),
            .in2(N__21277),
            .in3(N__21069),
            .lcout(buf_adcdata_vac_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55146),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_3_i19_3_lut_LC_6_11_1.C_ON=1'b0;
    defparam mux_130_Mux_3_i19_3_lut_LC_6_11_1.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_3_i19_3_lut_LC_6_11_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_130_Mux_3_i19_3_lut_LC_6_11_1 (
            .in0(N__23179),
            .in1(N__21474),
            .in2(_gnd_net_),
            .in3(N__56905),
            .lcout(),
            .ltout(n19_adj_1610_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_3_i22_3_lut_LC_6_11_2.C_ON=1'b0;
    defparam mux_130_Mux_3_i22_3_lut_LC_6_11_2.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_3_i22_3_lut_LC_6_11_2.LUT_INIT=16'b1111001111000000;
    LogicCell40 mux_130_Mux_3_i22_3_lut_LC_6_11_2 (
            .in0(_gnd_net_),
            .in1(N__47741),
            .in2(N__21049),
            .in3(N__21038),
            .lcout(n22_adj_1611),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i0_LC_6_11_3 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i0_LC_6_11_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i0_LC_6_11_3 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i0_LC_6_11_3  (
            .in0(N__50906),
            .in1(N__48997),
            .in2(N__21451),
            .in3(N__23450),
            .lcout(buf_adcdata_iac_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55146),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i21_LC_6_11_5 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i21_LC_6_11_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i21_LC_6_11_5 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i21_LC_6_11_5  (
            .in0(N__21557),
            .in1(N__48320),
            .in2(N__24142),
            .in3(N__37870),
            .lcout(cmd_rdadctmp_21_adj_1422),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55146),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i26_LC_6_12_1 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i26_LC_6_12_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i26_LC_6_12_1 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i26_LC_6_12_1  (
            .in0(N__37874),
            .in1(N__24235),
            .in2(N__48346),
            .in3(N__21290),
            .lcout(cmd_rdadctmp_26_adj_1417),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55161),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i30_LC_6_12_2 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i30_LC_6_12_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i30_LC_6_12_2 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i30_LC_6_12_2  (
            .in0(N__22619),
            .in1(N__48325),
            .in2(N__21345),
            .in3(N__37876),
            .lcout(cmd_rdadctmp_30_adj_1413),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55161),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i10_LC_6_12_3 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i10_LC_6_12_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i10_LC_6_12_3 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i10_LC_6_12_3  (
            .in0(N__21314),
            .in1(N__21252),
            .in2(N__50910),
            .in3(N__50514),
            .lcout(cmd_rdadctmp_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55161),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i24_LC_6_12_4 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i24_LC_6_12_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i24_LC_6_12_4 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i24_LC_6_12_4  (
            .in0(N__24251),
            .in1(N__48323),
            .in2(N__21237),
            .in3(N__37873),
            .lcout(cmd_rdadctmp_24_adj_1419),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55161),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i27_LC_6_12_6 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i27_LC_6_12_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i27_LC_6_12_6 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i27_LC_6_12_6  (
            .in0(N__21269),
            .in1(N__48324),
            .in2(N__21297),
            .in3(N__37875),
            .lcout(cmd_rdadctmp_27_adj_1416),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55161),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i1_LC_6_12_7 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i1_LC_6_12_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i1_LC_6_12_7 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_IAC.ADC_DATA_i1_LC_6_12_7  (
            .in0(N__48990),
            .in1(N__50936),
            .in2(N__23627),
            .in3(N__21253),
            .lcout(buf_adcdata_iac_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55161),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i23_LC_6_13_0 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i23_LC_6_13_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i23_LC_6_13_0 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i23_LC_6_13_0  (
            .in0(N__48196),
            .in1(N__21230),
            .in2(N__21420),
            .in3(N__37840),
            .lcout(cmd_rdadctmp_23_adj_1420),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55176),
            .ce(),
            .sr(_gnd_net_));
    defparam i18241_3_lut_LC_6_13_1.C_ON=1'b0;
    defparam i18241_3_lut_LC_6_13_1.SEQ_MODE=4'b0000;
    defparam i18241_3_lut_LC_6_13_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 i18241_3_lut_LC_6_13_1 (
            .in0(N__21672),
            .in1(N__24268),
            .in2(_gnd_net_),
            .in3(N__57485),
            .lcout(n20836),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i11_LC_6_13_2 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i11_LC_6_13_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i11_LC_6_13_2 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i11_LC_6_13_2  (
            .in0(N__48195),
            .in1(N__22838),
            .in2(N__22566),
            .in3(N__37838),
            .lcout(cmd_rdadctmp_11_adj_1432),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55176),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i3_LC_6_13_3 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i3_LC_6_13_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i3_LC_6_13_3 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i3_LC_6_13_3  (
            .in0(N__48493),
            .in1(N__48197),
            .in2(N__22845),
            .in3(N__21473),
            .lcout(buf_adcdata_vac_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55176),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i14_LC_6_13_4 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i14_LC_6_13_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i14_LC_6_13_4 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i14_LC_6_13_4  (
            .in0(N__48194),
            .in1(N__48494),
            .in2(N__21421),
            .in3(N__22677),
            .lcout(buf_adcdata_vac_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55176),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i8_LC_6_13_6 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i8_LC_6_13_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i8_LC_6_13_6 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i8_LC_6_13_6  (
            .in0(N__24286),
            .in1(N__50953),
            .in2(N__21446),
            .in3(N__50513),
            .lcout(cmd_rdadctmp_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55176),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i22_LC_6_13_7 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i22_LC_6_13_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i22_LC_6_13_7 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i22_LC_6_13_7  (
            .in0(N__37839),
            .in1(N__21413),
            .in2(N__21568),
            .in3(N__48198),
            .lcout(cmd_rdadctmp_22_adj_1421),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55176),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i8_LC_6_14_1 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i8_LC_6_14_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i8_LC_6_14_1 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \ADC_VAC.ADC_DATA_i8_LC_6_14_1  (
            .in0(N__48439),
            .in1(N__21387),
            .in2(N__48265),
            .in3(N__22726),
            .lcout(buf_adcdata_vac_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55191),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_5_i19_3_lut_LC_6_14_2.C_ON=1'b0;
    defparam mux_129_Mux_5_i19_3_lut_LC_6_14_2.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_5_i19_3_lut_LC_6_14_2.LUT_INIT=16'b1100110010101010;
    LogicCell40 mux_129_Mux_5_i19_3_lut_LC_6_14_2 (
            .in0(N__21533),
            .in1(N__23350),
            .in2(_gnd_net_),
            .in3(N__56907),
            .lcout(n19_adj_1487),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_0_i19_3_lut_LC_6_14_3.C_ON=1'b0;
    defparam mux_129_Mux_0_i19_3_lut_LC_6_14_3.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_0_i19_3_lut_LC_6_14_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_129_Mux_0_i19_3_lut_LC_6_14_3 (
            .in0(N__56908),
            .in1(N__26635),
            .in2(_gnd_net_),
            .in3(N__21386),
            .lcout(),
            .ltout(n19_adj_1479_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19393_LC_6_14_4.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19393_LC_6_14_4.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19393_LC_6_14_4.LUT_INIT=16'b1101100010101010;
    LogicCell40 comm_cmd_1__bdd_4_lut_19393_LC_6_14_4 (
            .in0(N__57448),
            .in1(N__21373),
            .in2(N__21349),
            .in3(N__47821),
            .lcout(n21973),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_6_i23_3_lut_LC_6_14_6.C_ON=1'b0;
    defparam mux_128_Mux_6_i23_3_lut_LC_6_14_6.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_6_i23_3_lut_LC_6_14_6.LUT_INIT=16'b1110111000100010;
    LogicCell40 mux_128_Mux_6_i23_3_lut_LC_6_14_6 (
            .in0(N__55962),
            .in1(N__56906),
            .in2(_gnd_net_),
            .in3(N__36664),
            .lcout(),
            .ltout(n23_adj_1512_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18247_4_lut_LC_6_14_7.C_ON=1'b0;
    defparam i18247_4_lut_LC_6_14_7.SEQ_MODE=4'b0000;
    defparam i18247_4_lut_LC_6_14_7.LUT_INIT=16'b0111010000110000;
    LogicCell40 i18247_4_lut_LC_6_14_7 (
            .in0(N__56909),
            .in1(N__57449),
            .in2(N__21586),
            .in3(N__45235),
            .lcout(n20842),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i4_LC_6_15_1 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i4_LC_6_15_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i4_LC_6_15_1 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i4_LC_6_15_1  (
            .in0(N__21513),
            .in1(N__48113),
            .in2(N__22879),
            .in3(N__37785),
            .lcout(cmd_rdadctmp_4_adj_1439),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55205),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i6_LC_6_15_2 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i6_LC_6_15_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i6_LC_6_15_2 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i6_LC_6_15_2  (
            .in0(N__37787),
            .in1(N__21579),
            .in2(N__48202),
            .in3(N__21502),
            .lcout(cmd_rdadctmp_6_adj_1437),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55205),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i13_LC_6_15_3 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i13_LC_6_15_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i13_LC_6_15_3 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC.ADC_DATA_i13_LC_6_15_3  (
            .in0(N__48437),
            .in1(N__48112),
            .in2(N__21541),
            .in3(N__21567),
            .lcout(buf_adcdata_vac_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55205),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i5_LC_6_15_4 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i5_LC_6_15_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i5_LC_6_15_4 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i5_LC_6_15_4  (
            .in0(N__37786),
            .in1(N__21501),
            .in2(N__21517),
            .in3(N__48117),
            .lcout(cmd_rdadctmp_5_adj_1438),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55205),
            .ce(),
            .sr(_gnd_net_));
    defparam i19061_2_lut_LC_6_15_5.C_ON=1'b0;
    defparam i19061_2_lut_LC_6_15_5.SEQ_MODE=4'b0000;
    defparam i19061_2_lut_LC_6_15_5.LUT_INIT=16'b1111111111001100;
    LogicCell40 i19061_2_lut_LC_6_15_5 (
            .in0(_gnd_net_),
            .in1(N__21493),
            .in2(_gnd_net_),
            .in3(N__56910),
            .lcout(n21109),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i18_LC_6_15_6 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i18_LC_6_15_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i18_LC_6_15_6 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i18_LC_6_15_6  (
            .in0(N__50491),
            .in1(N__21696),
            .in2(N__50909),
            .in3(N__21725),
            .lcout(cmd_rdadctmp_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55205),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i17_LC_6_15_7 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i17_LC_6_15_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i17_LC_6_15_7 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i17_LC_6_15_7  (
            .in0(N__21695),
            .in1(N__50830),
            .in2(N__45139),
            .in3(N__50492),
            .lcout(cmd_rdadctmp_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55205),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i21_LC_6_16_1 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i21_LC_6_16_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i21_LC_6_16_1 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i21_LC_6_16_1  (
            .in0(N__21776),
            .in1(N__50856),
            .in2(N__21802),
            .in3(N__50496),
            .lcout(cmd_rdadctmp_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55217),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i19_LC_6_16_3 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i19_LC_6_16_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i19_LC_6_16_3 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i19_LC_6_16_3  (
            .in0(N__21752),
            .in1(N__50855),
            .in2(N__21732),
            .in3(N__50495),
            .lcout(cmd_rdadctmp_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55217),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i10_LC_6_17_5 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i10_LC_6_17_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i10_LC_6_17_5 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i10_LC_6_17_5  (
            .in0(N__48892),
            .in1(N__50960),
            .in2(N__21736),
            .in3(N__25961),
            .lcout(buf_adcdata_iac_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55228),
            .ce(),
            .sr(_gnd_net_));
    defparam i18806_2_lut_LC_6_17_7.C_ON=1'b0;
    defparam i18806_2_lut_LC_6_17_7.SEQ_MODE=4'b0000;
    defparam i18806_2_lut_LC_6_17_7.LUT_INIT=16'b0000000011001100;
    LogicCell40 i18806_2_lut_LC_6_17_7 (
            .in0(_gnd_net_),
            .in1(N__21709),
            .in2(_gnd_net_),
            .in3(N__56912),
            .lcout(n21285),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i9_LC_6_18_3 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i9_LC_6_18_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i9_LC_6_18_3 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i9_LC_6_18_3  (
            .in0(N__48873),
            .in1(N__50821),
            .in2(N__21700),
            .in3(N__21671),
            .lcout(buf_adcdata_iac_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55238),
            .ce(),
            .sr(_gnd_net_));
    defparam \pll_main.i19651_1_lut_LC_7_1_7 .C_ON=1'b0;
    defparam \pll_main.i19651_1_lut_LC_7_1_7 .SEQ_MODE=4'b0000;
    defparam \pll_main.i19651_1_lut_LC_7_1_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pll_main.i19651_1_lut_LC_7_1_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56040),
            .lcout(DDS_MCLK1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.bit_cnt_i0_LC_7_4_5 .C_ON=1'b0;
    defparam \CLK_DDS.bit_cnt_i0_LC_7_4_5 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.bit_cnt_i0_LC_7_4_5 .LUT_INIT=16'b0000111101000000;
    LogicCell40 \CLK_DDS.bit_cnt_i0_LC_7_4_5  (
            .in0(N__28776),
            .in1(N__28607),
            .in2(N__28942),
            .in3(N__23233),
            .lcout(bit_cnt_0_adj_1449),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55076),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.CS_28_LC_7_5_3 .C_ON=1'b0;
    defparam \CLK_DDS.CS_28_LC_7_5_3 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.CS_28_LC_7_5_3 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \CLK_DDS.CS_28_LC_7_5_3  (
            .in0(N__28876),
            .in1(N__28773),
            .in2(_gnd_net_),
            .in3(N__28613),
            .lcout(DDS_CS1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55083),
            .ce(N__23269),
            .sr(_gnd_net_));
    defparam \CLK_DDS.SCLK_27_LC_7_7_4 .C_ON=1'b0;
    defparam \CLK_DDS.SCLK_27_LC_7_7_4 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.SCLK_27_LC_7_7_4 .LUT_INIT=16'b0101010011010001;
    LogicCell40 \CLK_DDS.SCLK_27_LC_7_7_4  (
            .in0(N__28750),
            .in1(N__28617),
            .in2(N__21603),
            .in3(N__28880),
            .lcout(DDS_SCK1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55096),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i2_2_lut_3_lut_LC_7_7_6 .C_ON=1'b0;
    defparam \RTD.i2_2_lut_3_lut_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \RTD.i2_2_lut_3_lut_LC_7_7_6 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \RTD.i2_2_lut_3_lut_LC_7_7_6  (
            .in0(N__22333),
            .in1(N__22195),
            .in2(_gnd_net_),
            .in3(N__22103),
            .lcout(\RTD.n20487 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.dds_state_i2_LC_7_9_1 .C_ON=1'b0;
    defparam \CLK_DDS.dds_state_i2_LC_7_9_1 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.dds_state_i2_LC_7_9_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \CLK_DDS.dds_state_i2_LC_7_9_1  (
            .in0(_gnd_net_),
            .in1(N__28941),
            .in2(_gnd_net_),
            .in3(N__28736),
            .lcout(dds_state_2_adj_1445),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55113),
            .ce(),
            .sr(_gnd_net_));
    defparam i18248_4_lut_LC_7_9_3.C_ON=1'b0;
    defparam i18248_4_lut_LC_7_9_3.SEQ_MODE=4'b0000;
    defparam i18248_4_lut_LC_7_9_3.LUT_INIT=16'b0011000010001000;
    LogicCell40 i18248_4_lut_LC_7_9_3 (
            .in0(N__21889),
            .in1(N__57187),
            .in2(N__31339),
            .in3(N__56982),
            .lcout(n20843),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.MOSI_31_LC_7_9_4 .C_ON=1'b0;
    defparam \CLK_DDS.MOSI_31_LC_7_9_4 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.MOSI_31_LC_7_9_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \CLK_DDS.MOSI_31_LC_7_9_4  (
            .in0(N__28940),
            .in1(N__27726),
            .in2(_gnd_net_),
            .in3(N__21867),
            .lcout(DDS_MOSI1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55113),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i1_LC_7_9_5.C_ON=1'b0;
    defparam buf_cfgRTD_i1_LC_7_9_5.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i1_LC_7_9_5.LUT_INIT=16'b0111010100100000;
    LogicCell40 buf_cfgRTD_i1_LC_7_9_5 (
            .in0(N__45331),
            .in1(N__52195),
            .in2(N__44146),
            .in3(N__23681),
            .lcout(buf_cfgRTD_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55113),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_217_LC_7_9_7.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_217_LC_7_9_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_217_LC_7_9_7.LUT_INIT=16'b0000000000100010;
    LogicCell40 i1_2_lut_3_lut_adj_217_LC_7_9_7 (
            .in0(N__41365),
            .in1(N__51298),
            .in2(_gnd_net_),
            .in3(N__54093),
            .lcout(n14_adj_1516),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22141_bdd_4_lut_LC_7_10_0.C_ON=1'b0;
    defparam n22141_bdd_4_lut_LC_7_10_0.SEQ_MODE=4'b0000;
    defparam n22141_bdd_4_lut_LC_7_10_0.LUT_INIT=16'b1100110011100010;
    LogicCell40 n22141_bdd_4_lut_LC_7_10_0 (
            .in0(N__22704),
            .in1(N__23404),
            .in2(N__23542),
            .in3(N__57191),
            .lcout(n20828),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22153_bdd_4_lut_LC_7_10_1.C_ON=1'b0;
    defparam n22153_bdd_4_lut_LC_7_10_1.SEQ_MODE=4'b0000;
    defparam n22153_bdd_4_lut_LC_7_10_1.LUT_INIT=16'b1100110011100010;
    LogicCell40 n22153_bdd_4_lut_LC_7_10_1 (
            .in0(N__21852),
            .in1(N__22501),
            .in2(N__23374),
            .in3(N__57188),
            .lcout(n22156),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19541_LC_7_10_2.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19541_LC_7_10_2.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19541_LC_7_10_2.LUT_INIT=16'b1110010010101010;
    LogicCell40 comm_cmd_0__bdd_4_lut_19541_LC_7_10_2 (
            .in0(N__56886),
            .in1(N__23717),
            .in2(N__21823),
            .in3(N__57192),
            .lcout(),
            .ltout(n22183_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22183_bdd_4_lut_LC_7_10_3.C_ON=1'b0;
    defparam n22183_bdd_4_lut_LC_7_10_3.SEQ_MODE=4'b0000;
    defparam n22183_bdd_4_lut_LC_7_10_3.LUT_INIT=16'b1111000010101100;
    LogicCell40 n22183_bdd_4_lut_LC_7_10_3 (
            .in0(N__23326),
            .in1(N__22596),
            .in2(N__22543),
            .in3(N__57190),
            .lcout(n20772),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22165_bdd_4_lut_LC_7_10_5.C_ON=1'b0;
    defparam n22165_bdd_4_lut_LC_7_10_5.SEQ_MODE=4'b0000;
    defparam n22165_bdd_4_lut_LC_7_10_5.LUT_INIT=16'b1100110011100010;
    LogicCell40 n22165_bdd_4_lut_LC_7_10_5 (
            .in0(N__22652),
            .in1(N__23635),
            .in2(N__23524),
            .in3(N__57189),
            .lcout(n20814),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_2_i30_3_lut_LC_7_10_7.C_ON=1'b0;
    defparam mux_130_Mux_2_i30_3_lut_LC_7_10_7.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_2_i30_3_lut_LC_7_10_7.LUT_INIT=16'b1111000010101010;
    LogicCell40 mux_130_Mux_2_i30_3_lut_LC_7_10_7 (
            .in0(N__22465),
            .in1(_gnd_net_),
            .in2(N__22540),
            .in3(N__56271),
            .lcout(n30_adj_1615),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19521_LC_7_11_0.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19521_LC_7_11_0.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19521_LC_7_11_0.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_0__bdd_4_lut_19521_LC_7_11_0 (
            .in0(N__41425),
            .in1(N__57182),
            .in2(N__22525),
            .in3(N__56865),
            .lcout(n22153),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i0_LC_7_11_1 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i0_LC_7_11_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i0_LC_7_11_1 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i0_LC_7_11_1  (
            .in0(N__48524),
            .in1(N__48179),
            .in2(N__22807),
            .in3(N__23477),
            .lcout(buf_adcdata_vac_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55134),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_2_i19_3_lut_LC_7_11_2.C_ON=1'b0;
    defparam mux_130_Mux_2_i19_3_lut_LC_7_11_2.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_2_i19_3_lut_LC_7_11_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_130_Mux_2_i19_3_lut_LC_7_11_2 (
            .in0(N__23308),
            .in1(N__22424),
            .in2(_gnd_net_),
            .in3(N__56867),
            .lcout(),
            .ltout(n19_adj_1613_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_2_i22_3_lut_LC_7_11_3.C_ON=1'b0;
    defparam mux_130_Mux_2_i22_3_lut_LC_7_11_3.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_2_i22_3_lut_LC_7_11_3.LUT_INIT=16'b1111000010101010;
    LogicCell40 mux_130_Mux_2_i22_3_lut_LC_7_11_3 (
            .in0(N__22491),
            .in1(_gnd_net_),
            .in2(N__22468),
            .in3(N__47742),
            .lcout(n22_adj_1614),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19501_LC_7_11_5.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19501_LC_7_11_5.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19501_LC_7_11_5.LUT_INIT=16'b1110010010101010;
    LogicCell40 comm_cmd_0__bdd_4_lut_19501_LC_7_11_5 (
            .in0(N__56866),
            .in1(N__24175),
            .in2(N__22459),
            .in3(N__57181),
            .lcout(n22135),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i2_LC_7_11_6 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i2_LC_7_11_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i2_LC_7_11_6 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i2_LC_7_11_6  (
            .in0(N__48178),
            .in1(N__48525),
            .in2(N__22570),
            .in3(N__22425),
            .lcout(buf_adcdata_vac_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55134),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i22_LC_7_12_0 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i22_LC_7_12_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i22_LC_7_12_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i22_LC_7_12_0  (
            .in0(N__48508),
            .in1(N__48176),
            .in2(N__22627),
            .in3(N__22703),
            .lcout(buf_adcdata_vac_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55147),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_6_i19_3_lut_LC_7_12_2.C_ON=1'b0;
    defparam mux_129_Mux_6_i19_3_lut_LC_7_12_2.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_6_i19_3_lut_LC_7_12_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_129_Mux_6_i19_3_lut_LC_7_12_2 (
            .in0(N__56883),
            .in1(N__23560),
            .in2(_gnd_net_),
            .in3(N__22673),
            .lcout(n19_adj_1482),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i17_LC_7_12_3 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i17_LC_7_12_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i17_LC_7_12_3 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC.ADC_DATA_i17_LC_7_12_3  (
            .in0(N__48173),
            .in1(N__48509),
            .in2(N__22656),
            .in3(N__24234),
            .lcout(buf_adcdata_vac_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55147),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i31_LC_7_12_4 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i31_LC_7_12_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i31_LC_7_12_4 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i31_LC_7_12_4  (
            .in0(N__22605),
            .in1(N__48177),
            .in2(N__22626),
            .in3(N__37844),
            .lcout(cmd_rdadctmp_31_adj_1412),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55147),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i23_LC_7_12_5 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i23_LC_7_12_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i23_LC_7_12_5 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC.ADC_DATA_i23_LC_7_12_5  (
            .in0(N__48174),
            .in1(N__48510),
            .in2(N__24338),
            .in3(N__22606),
            .lcout(buf_adcdata_vac_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55147),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i16_LC_7_12_6 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i16_LC_7_12_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i16_LC_7_12_6 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC.ADC_DATA_i16_LC_7_12_6  (
            .in0(N__48507),
            .in1(N__48175),
            .in2(N__22597),
            .in3(N__24255),
            .lcout(buf_adcdata_vac_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55147),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i18_LC_7_13_0 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i18_LC_7_13_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i18_LC_7_13_0 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i18_LC_7_13_0  (
            .in0(N__37834),
            .in1(N__22740),
            .in2(N__48262),
            .in3(N__24110),
            .lcout(cmd_rdadctmp_18_adj_1425),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55162),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i1_LC_7_13_1 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i1_LC_7_13_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i1_LC_7_13_1 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i1_LC_7_13_1  (
            .in0(N__48478),
            .in1(N__48181),
            .in2(N__22783),
            .in3(N__23960),
            .lcout(buf_adcdata_vac_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55162),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i9_LC_7_13_2 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i9_LC_7_13_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i9_LC_7_13_2 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC.ADC_DATA_i9_LC_7_13_2  (
            .in0(N__48180),
            .in1(N__48479),
            .in2(N__35276),
            .in3(N__22741),
            .lcout(buf_adcdata_vac_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55162),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i10_LC_7_13_3 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i10_LC_7_13_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i10_LC_7_13_3 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i10_LC_7_13_3  (
            .in0(N__22559),
            .in1(N__48182),
            .in2(N__22782),
            .in3(N__37832),
            .lcout(cmd_rdadctmp_10_adj_1433),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55162),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i19_LC_7_13_4 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i19_LC_7_13_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i19_LC_7_13_4 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i19_LC_7_13_4  (
            .in0(N__37835),
            .in1(N__24111),
            .in2(N__48263),
            .in3(N__24020),
            .lcout(cmd_rdadctmp_19_adj_1424),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55162),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i12_LC_7_13_5 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i12_LC_7_13_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i12_LC_7_13_5 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i12_LC_7_13_5  (
            .in0(N__47948),
            .in1(N__48183),
            .in2(N__22846),
            .in3(N__37833),
            .lcout(cmd_rdadctmp_12_adj_1431),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55162),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i8_LC_7_13_6 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i8_LC_7_13_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i8_LC_7_13_6 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i8_LC_7_13_6  (
            .in0(N__37836),
            .in1(N__22796),
            .in2(N__48264),
            .in3(N__22825),
            .lcout(cmd_rdadctmp_8_adj_1435),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55162),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i9_LC_7_13_7 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i9_LC_7_13_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i9_LC_7_13_7 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i9_LC_7_13_7  (
            .in0(N__22775),
            .in1(N__48184),
            .in2(N__22803),
            .in3(N__37837),
            .lcout(cmd_rdadctmp_9_adj_1434),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55162),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i0_LC_7_14_0 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i0_LC_7_14_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i0_LC_7_14_0 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i0_LC_7_14_0  (
            .in0(N__22905),
            .in1(N__48223),
            .in2(N__22765),
            .in3(N__37779),
            .lcout(cmd_rdadctmp_0_adj_1443),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55177),
            .ce(),
            .sr(_gnd_net_));
    defparam n21973_bdd_4_lut_LC_7_14_1.C_ON=1'b0;
    defparam n21973_bdd_4_lut_LC_7_14_1.SEQ_MODE=4'b0000;
    defparam n21973_bdd_4_lut_LC_7_14_1.LUT_INIT=16'b1100110011100010;
    LogicCell40 n21973_bdd_4_lut_LC_7_14_1 (
            .in0(N__27838),
            .in1(N__22747),
            .in2(N__24420),
            .in3(N__47822),
            .lcout(n21976),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i17_LC_7_14_3 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i17_LC_7_14_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i17_LC_7_14_3 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i17_LC_7_14_3  (
            .in0(N__37781),
            .in1(N__22725),
            .in2(N__48281),
            .in3(N__22739),
            .lcout(cmd_rdadctmp_17_adj_1426),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55177),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i16_LC_7_14_4 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i16_LC_7_14_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i16_LC_7_14_4 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i16_LC_7_14_4  (
            .in0(N__22724),
            .in1(N__48224),
            .in2(N__45205),
            .in3(N__37780),
            .lcout(cmd_rdadctmp_16_adj_1427),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55177),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i2_LC_7_14_5 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i2_LC_7_14_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i2_LC_7_14_5 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i2_LC_7_14_5  (
            .in0(N__37783),
            .in1(N__22897),
            .in2(N__48282),
            .in3(N__22887),
            .lcout(cmd_rdadctmp_2_adj_1441),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55177),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i1_LC_7_14_6 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i1_LC_7_14_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i1_LC_7_14_6 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i1_LC_7_14_6  (
            .in0(N__22896),
            .in1(N__48225),
            .in2(N__22909),
            .in3(N__37782),
            .lcout(cmd_rdadctmp_1_adj_1442),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55177),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i3_LC_7_14_7 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i3_LC_7_14_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i3_LC_7_14_7 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i3_LC_7_14_7  (
            .in0(N__37784),
            .in1(N__22888),
            .in2(N__48283),
            .in3(N__22875),
            .lcout(cmd_rdadctmp_3_adj_1440),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55177),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i1_3_lut_LC_7_15_0 .C_ON=1'b0;
    defparam \ADC_VAC.i1_3_lut_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i1_3_lut_LC_7_15_0 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \ADC_VAC.i1_3_lut_LC_7_15_0  (
            .in0(N__48040),
            .in1(N__22993),
            .in2(_gnd_net_),
            .in3(N__22864),
            .lcout(n12643),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.adc_state_i2_LC_7_15_1 .C_ON=1'b0;
    defparam \ADC_VAC.adc_state_i2_LC_7_15_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.adc_state_i2_LC_7_15_1 .LUT_INIT=16'b0110011000100010;
    LogicCell40 \ADC_VAC.adc_state_i2_LC_7_15_1  (
            .in0(N__29766),
            .in1(N__29845),
            .in2(_gnd_net_),
            .in3(N__48042),
            .lcout(DTRIG_N_910_adj_1444),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55192),
            .ce(N__22951),
            .sr(_gnd_net_));
    defparam \ADC_VAC.adc_state_i1_LC_7_15_2 .C_ON=1'b0;
    defparam \ADC_VAC.adc_state_i1_LC_7_15_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.adc_state_i1_LC_7_15_2 .LUT_INIT=16'b0000000011110101;
    LogicCell40 \ADC_VAC.adc_state_i1_LC_7_15_2  (
            .in0(N__48041),
            .in1(_gnd_net_),
            .in2(N__29858),
            .in3(N__29767),
            .lcout(adc_state_1_adj_1410),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55192),
            .ce(N__22951),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i1_4_lut_adj_4_LC_7_15_4 .C_ON=1'b0;
    defparam \ADC_VAC.i1_4_lut_adj_4_LC_7_15_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i1_4_lut_adj_4_LC_7_15_4 .LUT_INIT=16'b0001000000010100;
    LogicCell40 \ADC_VAC.i1_4_lut_adj_4_LC_7_15_4  (
            .in0(N__48039),
            .in1(N__29765),
            .in2(N__29857),
            .in3(N__22994),
            .lcout(\ADC_VAC.n12556 ),
            .ltout(\ADC_VAC.n12556_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i12432_2_lut_LC_7_15_5 .C_ON=1'b0;
    defparam \ADC_VAC.i12432_2_lut_LC_7_15_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i12432_2_lut_LC_7_15_5 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \ADC_VAC.i12432_2_lut_LC_7_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22855),
            .in3(N__29841),
            .lcout(\ADC_VAC.n14829 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_118_LC_7_15_7.C_ON=1'b0;
    defparam i1_2_lut_adj_118_LC_7_15_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_118_LC_7_15_7.LUT_INIT=16'b0011001100000000;
    LogicCell40 i1_2_lut_adj_118_LC_7_15_7 (
            .in0(_gnd_net_),
            .in1(N__29764),
            .in2(_gnd_net_),
            .in3(N__29837),
            .lcout(n20540),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i1_2_lut_adj_3_LC_7_16_0 .C_ON=1'b0;
    defparam \ADC_VAC.i1_2_lut_adj_3_LC_7_16_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i1_2_lut_adj_3_LC_7_16_0 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \ADC_VAC.i1_2_lut_adj_3_LC_7_16_0  (
            .in0(N__29787),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22852),
            .lcout(\ADC_VAC.n20668 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i1_4_lut_LC_7_16_1 .C_ON=1'b0;
    defparam \ADC_VAC.i1_4_lut_LC_7_16_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i1_4_lut_LC_7_16_1 .LUT_INIT=16'b1100110111101111;
    LogicCell40 \ADC_VAC.i1_4_lut_LC_7_16_1  (
            .in0(N__29846),
            .in1(N__48035),
            .in2(N__22999),
            .in3(N__30141),
            .lcout(\ADC_VAC.n20667 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i18152_4_lut_LC_7_16_2 .C_ON=1'b0;
    defparam \ADC_VAC.i18152_4_lut_LC_7_16_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i18152_4_lut_LC_7_16_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VAC.i18152_4_lut_LC_7_16_2  (
            .in0(N__23104),
            .in1(N__23118),
            .in2(N__22927),
            .in3(N__23133),
            .lcout(),
            .ltout(\ADC_VAC.n20747_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i18168_4_lut_LC_7_16_3 .C_ON=1'b0;
    defparam \ADC_VAC.i18168_4_lut_LC_7_16_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i18168_4_lut_LC_7_16_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VAC.i18168_4_lut_LC_7_16_3  (
            .in0(N__23070),
            .in1(N__22941),
            .in2(N__23017),
            .in3(N__23052),
            .lcout(),
            .ltout(\ADC_VAC.n20763_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i19024_4_lut_LC_7_16_4 .C_ON=1'b0;
    defparam \ADC_VAC.i19024_4_lut_LC_7_16_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i19024_4_lut_LC_7_16_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \ADC_VAC.i19024_4_lut_LC_7_16_4  (
            .in0(N__48037),
            .in1(N__23085),
            .in2(N__23014),
            .in3(N__29791),
            .lcout(),
            .ltout(\ADC_VAC.n21031_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.adc_state_i0_LC_7_16_5 .C_ON=1'b0;
    defparam \ADC_VAC.adc_state_i0_LC_7_16_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.adc_state_i0_LC_7_16_5 .LUT_INIT=16'b0011000001110100;
    LogicCell40 \ADC_VAC.adc_state_i0_LC_7_16_5  (
            .in0(N__29792),
            .in1(N__29862),
            .in2(N__23011),
            .in3(N__48038),
            .lcout(adc_state_0_adj_1411),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55206),
            .ce(N__23008),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i30_4_lut_LC_7_16_6 .C_ON=1'b0;
    defparam \ADC_VAC.i30_4_lut_LC_7_16_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i30_4_lut_LC_7_16_6 .LUT_INIT=16'b1011000110000001;
    LogicCell40 \ADC_VAC.i30_4_lut_LC_7_16_6  (
            .in0(N__30142),
            .in1(N__29847),
            .in2(N__29793),
            .in3(N__22998),
            .lcout(),
            .ltout(\ADC_VAC.n17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i19101_2_lut_LC_7_16_7 .C_ON=1'b0;
    defparam \ADC_VAC.i19101_2_lut_LC_7_16_7 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i19101_2_lut_LC_7_16_7 .LUT_INIT=16'b1111111100001111;
    LogicCell40 \ADC_VAC.i19101_2_lut_LC_7_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22954),
            .in3(N__48036),
            .lcout(\ADC_VAC.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.bit_cnt_i0_LC_7_17_0 .C_ON=1'b1;
    defparam \ADC_VAC.bit_cnt_i0_LC_7_17_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i0_LC_7_17_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i0_LC_7_17_0  (
            .in0(_gnd_net_),
            .in1(N__22942),
            .in2(_gnd_net_),
            .in3(N__22930),
            .lcout(\ADC_VAC.bit_cnt_0 ),
            .ltout(),
            .carryin(bfn_7_17_0_),
            .carryout(\ADC_VAC.n19357 ),
            .clk(N__55218),
            .ce(N__23041),
            .sr(N__23029));
    defparam \ADC_VAC.bit_cnt_i1_LC_7_17_1 .C_ON=1'b1;
    defparam \ADC_VAC.bit_cnt_i1_LC_7_17_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i1_LC_7_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i1_LC_7_17_1  (
            .in0(_gnd_net_),
            .in1(N__22926),
            .in2(_gnd_net_),
            .in3(N__22912),
            .lcout(\ADC_VAC.bit_cnt_1 ),
            .ltout(),
            .carryin(\ADC_VAC.n19357 ),
            .carryout(\ADC_VAC.n19358 ),
            .clk(N__55218),
            .ce(N__23041),
            .sr(N__23029));
    defparam \ADC_VAC.bit_cnt_i2_LC_7_17_2 .C_ON=1'b1;
    defparam \ADC_VAC.bit_cnt_i2_LC_7_17_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i2_LC_7_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i2_LC_7_17_2  (
            .in0(_gnd_net_),
            .in1(N__23134),
            .in2(_gnd_net_),
            .in3(N__23122),
            .lcout(\ADC_VAC.bit_cnt_2 ),
            .ltout(),
            .carryin(\ADC_VAC.n19358 ),
            .carryout(\ADC_VAC.n19359 ),
            .clk(N__55218),
            .ce(N__23041),
            .sr(N__23029));
    defparam \ADC_VAC.bit_cnt_i3_LC_7_17_3 .C_ON=1'b1;
    defparam \ADC_VAC.bit_cnt_i3_LC_7_17_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i3_LC_7_17_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i3_LC_7_17_3  (
            .in0(_gnd_net_),
            .in1(N__23119),
            .in2(_gnd_net_),
            .in3(N__23107),
            .lcout(\ADC_VAC.bit_cnt_3 ),
            .ltout(),
            .carryin(\ADC_VAC.n19359 ),
            .carryout(\ADC_VAC.n19360 ),
            .clk(N__55218),
            .ce(N__23041),
            .sr(N__23029));
    defparam \ADC_VAC.bit_cnt_i4_LC_7_17_4 .C_ON=1'b1;
    defparam \ADC_VAC.bit_cnt_i4_LC_7_17_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i4_LC_7_17_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i4_LC_7_17_4  (
            .in0(_gnd_net_),
            .in1(N__23103),
            .in2(_gnd_net_),
            .in3(N__23089),
            .lcout(\ADC_VAC.bit_cnt_4 ),
            .ltout(),
            .carryin(\ADC_VAC.n19360 ),
            .carryout(\ADC_VAC.n19361 ),
            .clk(N__55218),
            .ce(N__23041),
            .sr(N__23029));
    defparam \ADC_VAC.bit_cnt_i5_LC_7_17_5 .C_ON=1'b1;
    defparam \ADC_VAC.bit_cnt_i5_LC_7_17_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i5_LC_7_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i5_LC_7_17_5  (
            .in0(_gnd_net_),
            .in1(N__23086),
            .in2(_gnd_net_),
            .in3(N__23074),
            .lcout(\ADC_VAC.bit_cnt_5 ),
            .ltout(),
            .carryin(\ADC_VAC.n19361 ),
            .carryout(\ADC_VAC.n19362 ),
            .clk(N__55218),
            .ce(N__23041),
            .sr(N__23029));
    defparam \ADC_VAC.bit_cnt_i6_LC_7_17_6 .C_ON=1'b1;
    defparam \ADC_VAC.bit_cnt_i6_LC_7_17_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i6_LC_7_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i6_LC_7_17_6  (
            .in0(_gnd_net_),
            .in1(N__23071),
            .in2(_gnd_net_),
            .in3(N__23059),
            .lcout(\ADC_VAC.bit_cnt_6 ),
            .ltout(),
            .carryin(\ADC_VAC.n19362 ),
            .carryout(\ADC_VAC.n19363 ),
            .clk(N__55218),
            .ce(N__23041),
            .sr(N__23029));
    defparam \ADC_VAC.bit_cnt_i7_LC_7_17_7 .C_ON=1'b0;
    defparam \ADC_VAC.bit_cnt_i7_LC_7_17_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i7_LC_7_17_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i7_LC_7_17_7  (
            .in0(_gnd_net_),
            .in1(N__23053),
            .in2(_gnd_net_),
            .in3(N__23056),
            .lcout(\ADC_VAC.bit_cnt_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55218),
            .ce(N__23041),
            .sr(N__23029));
    defparam \ADC_IAC.i1_3_lut_LC_7_18_0 .C_ON=1'b0;
    defparam \ADC_IAC.i1_3_lut_LC_7_18_0 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i1_3_lut_LC_7_18_0 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \ADC_IAC.i1_3_lut_LC_7_18_0  (
            .in0(N__25007),
            .in1(N__50645),
            .in2(_gnd_net_),
            .in3(N__24657),
            .lcout(n12542),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.adc_state_i2_LC_7_18_1 .C_ON=1'b0;
    defparam \ADC_IAC.adc_state_i2_LC_7_18_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.adc_state_i2_LC_7_18_1 .LUT_INIT=16'b0011001110001000;
    LogicCell40 \ADC_IAC.adc_state_i2_LC_7_18_1  (
            .in0(N__50647),
            .in1(N__29999),
            .in2(_gnd_net_),
            .in3(N__29930),
            .lcout(DTRIG_N_910),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55229),
            .ce(N__24955),
            .sr(_gnd_net_));
    defparam \ADC_IAC.adc_state_i1_LC_7_18_2 .C_ON=1'b0;
    defparam \ADC_IAC.adc_state_i1_LC_7_18_2 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.adc_state_i1_LC_7_18_2 .LUT_INIT=16'b0101000001010101;
    LogicCell40 \ADC_IAC.adc_state_i1_LC_7_18_2  (
            .in0(N__29931),
            .in1(_gnd_net_),
            .in2(N__30013),
            .in3(N__50648),
            .lcout(adc_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55229),
            .ce(N__24955),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i1_2_lut_LC_7_18_3 .C_ON=1'b0;
    defparam \ADC_IAC.i1_2_lut_LC_7_18_3 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i1_2_lut_LC_7_18_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \ADC_IAC.i1_2_lut_LC_7_18_3  (
            .in0(_gnd_net_),
            .in1(N__29990),
            .in2(_gnd_net_),
            .in3(N__29927),
            .lcout(n20553),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i1_4_lut_adj_6_LC_7_18_4 .C_ON=1'b0;
    defparam \ADC_IAC.i1_4_lut_adj_6_LC_7_18_4 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i1_4_lut_adj_6_LC_7_18_4 .LUT_INIT=16'b0000000001010010;
    LogicCell40 \ADC_IAC.i1_4_lut_adj_6_LC_7_18_4  (
            .in0(N__29928),
            .in1(N__25008),
            .in2(N__30012),
            .in3(N__50646),
            .lcout(\ADC_IAC.n12459 ),
            .ltout(\ADC_IAC.n12459_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i12394_2_lut_LC_7_18_5 .C_ON=1'b0;
    defparam \ADC_IAC.i12394_2_lut_LC_7_18_5 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i12394_2_lut_LC_7_18_5 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \ADC_IAC.i12394_2_lut_LC_7_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23155),
            .in3(N__29995),
            .lcout(\ADC_IAC.n14791 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_83_LC_7_18_7.C_ON=1'b0;
    defparam i1_2_lut_adj_83_LC_7_18_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_83_LC_7_18_7.LUT_INIT=16'b0000000011001100;
    LogicCell40 i1_2_lut_adj_83_LC_7_18_7 (
            .in0(_gnd_net_),
            .in1(N__29994),
            .in2(_gnd_net_),
            .in3(N__29929),
            .lcout(n20543),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.bit_cnt_i0_LC_7_19_0 .C_ON=1'b1;
    defparam \ADC_IAC.bit_cnt_i0_LC_7_19_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i0_LC_7_19_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i0_LC_7_19_0  (
            .in0(_gnd_net_),
            .in1(N__24745),
            .in2(_gnd_net_),
            .in3(N__23152),
            .lcout(\ADC_IAC.bit_cnt_0 ),
            .ltout(),
            .carryin(bfn_7_19_0_),
            .carryout(\ADC_IAC.n19350 ),
            .clk(N__55239),
            .ce(N__23254),
            .sr(N__23239));
    defparam \ADC_IAC.bit_cnt_i1_LC_7_19_1 .C_ON=1'b1;
    defparam \ADC_IAC.bit_cnt_i1_LC_7_19_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i1_LC_7_19_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i1_LC_7_19_1  (
            .in0(_gnd_net_),
            .in1(N__24783),
            .in2(_gnd_net_),
            .in3(N__23149),
            .lcout(\ADC_IAC.bit_cnt_1 ),
            .ltout(),
            .carryin(\ADC_IAC.n19350 ),
            .carryout(\ADC_IAC.n19351 ),
            .clk(N__55239),
            .ce(N__23254),
            .sr(N__23239));
    defparam \ADC_IAC.bit_cnt_i2_LC_7_19_2 .C_ON=1'b1;
    defparam \ADC_IAC.bit_cnt_i2_LC_7_19_2 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i2_LC_7_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i2_LC_7_19_2  (
            .in0(_gnd_net_),
            .in1(N__24769),
            .in2(_gnd_net_),
            .in3(N__23146),
            .lcout(\ADC_IAC.bit_cnt_2 ),
            .ltout(),
            .carryin(\ADC_IAC.n19351 ),
            .carryout(\ADC_IAC.n19352 ),
            .clk(N__55239),
            .ce(N__23254),
            .sr(N__23239));
    defparam \ADC_IAC.bit_cnt_i3_LC_7_19_3 .C_ON=1'b1;
    defparam \ADC_IAC.bit_cnt_i3_LC_7_19_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i3_LC_7_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i3_LC_7_19_3  (
            .in0(_gnd_net_),
            .in1(N__24796),
            .in2(_gnd_net_),
            .in3(N__23143),
            .lcout(\ADC_IAC.bit_cnt_3 ),
            .ltout(),
            .carryin(\ADC_IAC.n19352 ),
            .carryout(\ADC_IAC.n19353 ),
            .clk(N__55239),
            .ce(N__23254),
            .sr(N__23239));
    defparam \ADC_IAC.bit_cnt_i4_LC_7_19_4 .C_ON=1'b1;
    defparam \ADC_IAC.bit_cnt_i4_LC_7_19_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i4_LC_7_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i4_LC_7_19_4  (
            .in0(_gnd_net_),
            .in1(N__24808),
            .in2(_gnd_net_),
            .in3(N__23140),
            .lcout(\ADC_IAC.bit_cnt_4 ),
            .ltout(),
            .carryin(\ADC_IAC.n19353 ),
            .carryout(\ADC_IAC.n19354 ),
            .clk(N__55239),
            .ce(N__23254),
            .sr(N__23239));
    defparam \ADC_IAC.bit_cnt_i5_LC_7_19_5 .C_ON=1'b1;
    defparam \ADC_IAC.bit_cnt_i5_LC_7_19_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i5_LC_7_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i5_LC_7_19_5  (
            .in0(_gnd_net_),
            .in1(N__25041),
            .in2(_gnd_net_),
            .in3(N__23137),
            .lcout(\ADC_IAC.bit_cnt_5 ),
            .ltout(),
            .carryin(\ADC_IAC.n19354 ),
            .carryout(\ADC_IAC.n19355 ),
            .clk(N__55239),
            .ce(N__23254),
            .sr(N__23239));
    defparam \ADC_IAC.bit_cnt_i6_LC_7_19_6 .C_ON=1'b1;
    defparam \ADC_IAC.bit_cnt_i6_LC_7_19_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i6_LC_7_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i6_LC_7_19_6  (
            .in0(_gnd_net_),
            .in1(N__24757),
            .in2(_gnd_net_),
            .in3(N__23260),
            .lcout(\ADC_IAC.bit_cnt_6 ),
            .ltout(),
            .carryin(\ADC_IAC.n19355 ),
            .carryout(\ADC_IAC.n19356 ),
            .clk(N__55239),
            .ce(N__23254),
            .sr(N__23239));
    defparam \ADC_IAC.bit_cnt_i7_LC_7_19_7 .C_ON=1'b0;
    defparam \ADC_IAC.bit_cnt_i7_LC_7_19_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i7_LC_7_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i7_LC_7_19_7  (
            .in0(_gnd_net_),
            .in1(N__24730),
            .in2(_gnd_net_),
            .in3(N__23257),
            .lcout(\ADC_IAC.bit_cnt_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55239),
            .ce(N__23254),
            .sr(N__23239));
    defparam \ADC_VDC.i1_2_lut_adj_42_LC_8_4_3 .C_ON=1'b0;
    defparam \ADC_VDC.i1_2_lut_adj_42_LC_8_4_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_2_lut_adj_42_LC_8_4_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ADC_VDC.i1_2_lut_adj_42_LC_8_4_3  (
            .in0(_gnd_net_),
            .in1(N__34588),
            .in2(_gnd_net_),
            .in3(N__34361),
            .lcout(\ADC_VDC.n20345 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19022_2_lut_LC_8_4_5.C_ON=1'b0;
    defparam i19022_2_lut_LC_8_4_5.SEQ_MODE=4'b0000;
    defparam i19022_2_lut_LC_8_4_5.LUT_INIT=16'b1100110000000000;
    LogicCell40 i19022_2_lut_LC_8_4_5 (
            .in0(_gnd_net_),
            .in1(N__23229),
            .in2(_gnd_net_),
            .in3(N__23205),
            .lcout(n21206),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i9_LC_8_5_0 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i9_LC_8_5_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i9_LC_8_5_0 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i9_LC_8_5_0  (
            .in0(N__34365),
            .in1(N__25078),
            .in2(N__26884),
            .in3(N__26509),
            .lcout(cmd_rdadctmp_9_adj_1463),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32904),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i3_LC_8_5_1 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i3_LC_8_5_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i3_LC_8_5_1 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i3_LC_8_5_1  (
            .in0(N__28361),
            .in1(N__34629),
            .in2(N__23172),
            .in3(N__25222),
            .lcout(buf_adcdata_vdc_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32904),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i7_LC_8_5_2 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i7_LC_8_5_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i7_LC_8_5_2 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i7_LC_8_5_2  (
            .in0(N__34364),
            .in1(N__26528),
            .in2(N__26883),
            .in3(N__25122),
            .lcout(cmd_rdadctmp_7_adj_1465),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32904),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i10_LC_8_5_3 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i10_LC_8_5_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i10_LC_8_5_3 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i10_LC_8_5_3  (
            .in0(N__25077),
            .in1(N__34366),
            .in2(N__26988),
            .in3(N__26850),
            .lcout(cmd_rdadctmp_10_adj_1462),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32904),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i6_LC_8_5_4 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i6_LC_8_5_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i6_LC_8_5_4 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i6_LC_8_5_4  (
            .in0(N__34363),
            .in1(N__25121),
            .in2(N__26882),
            .in3(N__25149),
            .lcout(cmd_rdadctmp_6_adj_1466),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32904),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.i23_4_lut_LC_8_5_5 .C_ON=1'b0;
    defparam \CLK_DDS.i23_4_lut_LC_8_5_5 .SEQ_MODE=4'b0000;
    defparam \CLK_DDS.i23_4_lut_LC_8_5_5 .LUT_INIT=16'b1100110110011001;
    LogicCell40 \CLK_DDS.i23_4_lut_LC_8_5_5  (
            .in0(N__28943),
            .in1(N__28775),
            .in2(N__28677),
            .in3(N__28611),
            .lcout(\CLK_DDS.n9_adj_1386 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i5_LC_8_5_6 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i5_LC_8_5_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i5_LC_8_5_6 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i5_LC_8_5_6  (
            .in0(N__34362),
            .in1(N__25148),
            .in2(N__26881),
            .in3(N__26569),
            .lcout(cmd_rdadctmp_5_adj_1467),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32904),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i15_LC_8_5_7 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i15_LC_8_5_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i15_LC_8_5_7 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i15_LC_8_5_7  (
            .in0(N__26450),
            .in1(N__34367),
            .in2(N__25252),
            .in3(N__26851),
            .lcout(cmd_rdadctmp_15_adj_1457),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32904),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i14_LC_8_6_0 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i14_LC_8_6_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i14_LC_8_6_0 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i14_LC_8_6_0  (
            .in0(N__34370),
            .in1(N__25287),
            .in2(N__25248),
            .in3(N__26888),
            .lcout(cmd_rdadctmp_14_adj_1458),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32886),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i0_LC_8_6_1 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i0_LC_8_6_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i0_LC_8_6_1 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i0_LC_8_6_1  (
            .in0(N__28362),
            .in1(N__34631),
            .in2(N__23499),
            .in3(N__25318),
            .lcout(buf_adcdata_vdc_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32886),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i18_LC_8_6_2 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i18_LC_8_6_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i18_LC_8_6_2 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i18_LC_8_6_2  (
            .in0(N__34371),
            .in1(N__25193),
            .in2(N__26485),
            .in3(N__26889),
            .lcout(cmd_rdadctmp_18_adj_1454),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32886),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i1_LC_8_6_3 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i1_LC_8_6_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i1_LC_8_6_3 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i1_LC_8_6_3  (
            .in0(N__28364),
            .in1(N__34633),
            .in2(N__23985),
            .in3(N__25303),
            .lcout(buf_adcdata_vdc_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32886),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i19_LC_8_6_4 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i19_LC_8_6_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i19_LC_8_6_4 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i19_LC_8_6_4  (
            .in0(N__34372),
            .in1(N__26915),
            .in2(N__25198),
            .in3(N__26890),
            .lcout(cmd_rdadctmp_19_adj_1453),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32886),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i10_LC_8_6_5 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i10_LC_8_6_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i10_LC_8_6_5 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i10_LC_8_6_5  (
            .in0(N__28363),
            .in1(N__34632),
            .in2(N__24072),
            .in3(N__25444),
            .lcout(buf_adcdata_vdc_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32886),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i21_LC_8_6_6 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i21_LC_8_6_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i21_LC_8_6_6 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i21_LC_8_6_6  (
            .in0(N__34373),
            .in1(N__25463),
            .in2(N__26773),
            .in3(N__26891),
            .lcout(cmd_rdadctmp_21_adj_1451),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32886),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i13_LC_8_6_7 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i13_LC_8_6_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i13_LC_8_6_7 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i13_LC_8_6_7  (
            .in0(N__25286),
            .in1(N__26363),
            .in2(N__26895),
            .in3(N__34374),
            .lcout(cmd_rdadctmp_13_adj_1459),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32886),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i22_LC_8_7_2 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i22_LC_8_7_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i22_LC_8_7_2 .LUT_INIT=16'b0011101000001010;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i22_LC_8_7_2  (
            .in0(N__25424),
            .in1(N__34369),
            .in2(N__26896),
            .in3(N__25464),
            .lcout(cmd_rdadctmp_22_adj_1450),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32872),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i21_LC_8_8_0 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i21_LC_8_8_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i21_LC_8_8_0 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \ADC_VDC.ADC_DATA_i21_LC_8_8_0  (
            .in0(N__25519),
            .in1(N__34640),
            .in2(N__23367),
            .in3(N__28397),
            .lcout(buf_adcdata_vdc_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32908),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i20_LC_8_8_1 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i20_LC_8_8_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i20_LC_8_8_1 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \ADC_VDC.ADC_DATA_i20_LC_8_8_1  (
            .in0(N__34636),
            .in1(N__28419),
            .in2(N__25668),
            .in3(N__25534),
            .lcout(buf_adcdata_vdc_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32908),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i13_LC_8_8_2 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i13_LC_8_8_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i13_LC_8_8_2 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i13_LC_8_8_2  (
            .in0(N__28414),
            .in1(N__34637),
            .in2(N__23343),
            .in3(N__25378),
            .lcout(buf_adcdata_vdc_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32908),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i18_LC_8_8_3 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i18_LC_8_8_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i18_LC_8_8_3 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \ADC_VDC.ADC_DATA_i18_LC_8_8_3  (
            .in0(N__34635),
            .in1(N__28418),
            .in2(N__23874),
            .in3(N__25564),
            .lcout(buf_adcdata_vdc_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32908),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i16_LC_8_8_4 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i16_LC_8_8_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i16_LC_8_8_4 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i16_LC_8_8_4  (
            .in0(N__28415),
            .in1(N__34638),
            .in2(N__23325),
            .in3(N__25333),
            .lcout(buf_adcdata_vdc_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32908),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i2_LC_8_8_5 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i2_LC_8_8_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i2_LC_8_8_5 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \ADC_VDC.ADC_DATA_i2_LC_8_8_5  (
            .in0(N__25270),
            .in1(N__28420),
            .in2(N__23307),
            .in3(N__34641),
            .lcout(buf_adcdata_vdc_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32908),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i19_LC_8_8_6 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i19_LC_8_8_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i19_LC_8_8_6 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i19_LC_8_8_6  (
            .in0(N__28416),
            .in1(N__34639),
            .in2(N__23286),
            .in3(N__25549),
            .lcout(buf_adcdata_vdc_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32908),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i15_LC_8_8_7 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i15_LC_8_8_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i15_LC_8_8_7 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \ADC_VDC.ADC_DATA_i15_LC_8_8_7  (
            .in0(N__34634),
            .in1(N__28417),
            .in2(N__23577),
            .in3(N__25348),
            .lcout(buf_adcdata_vdc_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32908),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i14_LC_8_9_1 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i14_LC_8_9_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i14_LC_8_9_1 .LUT_INIT=16'b0010111100100000;
    LogicCell40 \ADC_VDC.ADC_DATA_i14_LC_8_9_1  (
            .in0(N__25363),
            .in1(N__34627),
            .in2(N__28398),
            .in3(N__23553),
            .lcout(buf_adcdata_vdc_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32885),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i22_LC_8_9_2 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i22_LC_8_9_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i22_LC_8_9_2 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \ADC_VDC.ADC_DATA_i22_LC_8_9_2  (
            .in0(N__34625),
            .in1(N__28390),
            .in2(N__23541),
            .in3(N__25504),
            .lcout(buf_adcdata_vdc_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32885),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i17_LC_8_9_3 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i17_LC_8_9_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i17_LC_8_9_3 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i17_LC_8_9_3  (
            .in0(N__28388),
            .in1(N__34626),
            .in2(N__23523),
            .in3(N__25579),
            .lcout(buf_adcdata_vdc_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32885),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_0_i19_3_lut_LC_8_9_4.C_ON=1'b0;
    defparam mux_130_Mux_0_i19_3_lut_LC_8_9_4.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_0_i19_3_lut_LC_8_9_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_130_Mux_0_i19_3_lut_LC_8_9_4 (
            .in0(N__23500),
            .in1(N__23478),
            .in2(_gnd_net_),
            .in3(N__56960),
            .lcout(),
            .ltout(n19_adj_1477_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_0_i22_3_lut_LC_8_9_5.C_ON=1'b0;
    defparam mux_130_Mux_0_i22_3_lut_LC_8_9_5.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_0_i22_3_lut_LC_8_9_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 mux_130_Mux_0_i22_3_lut_LC_8_9_5 (
            .in0(_gnd_net_),
            .in1(N__23457),
            .in2(N__23431),
            .in3(N__47774),
            .lcout(n22_adj_1476),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19506_LC_8_9_6.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19506_LC_8_9_6.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19506_LC_8_9_6.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_0__bdd_4_lut_19506_LC_8_9_6 (
            .in0(N__29317),
            .in1(N__57183),
            .in2(N__23428),
            .in3(N__56959),
            .lcout(n22141),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i23_LC_8_9_7 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i23_LC_8_9_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i23_LC_8_9_7 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \ADC_VDC.ADC_DATA_i23_LC_8_9_7  (
            .in0(N__28389),
            .in1(N__27055),
            .in2(N__24309),
            .in3(N__34628),
            .lcout(buf_adcdata_vdc_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32885),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19388_LC_8_10_0.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19388_LC_8_10_0.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19388_LC_8_10_0.LUT_INIT=16'b1101101010001010;
    LogicCell40 comm_cmd_0__bdd_4_lut_19388_LC_8_10_0 (
            .in0(N__56885),
            .in1(N__23398),
            .in2(N__57465),
            .in3(N__23805),
            .lcout(),
            .ltout(n21931_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n21931_bdd_4_lut_LC_8_10_1.C_ON=1'b0;
    defparam n21931_bdd_4_lut_LC_8_10_1.SEQ_MODE=4'b0000;
    defparam n21931_bdd_4_lut_LC_8_10_1.LUT_INIT=16'b1111000010101100;
    LogicCell40 n21931_bdd_4_lut_LC_8_10_1 (
            .in0(N__23878),
            .in1(N__23857),
            .in2(N__23830),
            .in3(N__57345),
            .lcout(n21934),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i2_LC_8_10_2.C_ON=1'b0;
    defparam buf_cfgRTD_i2_LC_8_10_2.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i2_LC_8_10_2.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_cfgRTD_i2_LC_8_10_2 (
            .in0(N__52190),
            .in1(N__45329),
            .in2(N__38729),
            .in3(N__23806),
            .lcout(buf_cfgRTD_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55114),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i3_LC_8_10_3.C_ON=1'b0;
    defparam buf_cfgRTD_i3_LC_8_10_3.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i3_LC_8_10_3.LUT_INIT=16'b0111010100100000;
    LogicCell40 buf_cfgRTD_i3_LC_8_10_3 (
            .in0(N__45330),
            .in1(N__52191),
            .in2(N__43760),
            .in3(N__23763),
            .lcout(buf_cfgRTD_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55114),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i0_LC_8_10_4.C_ON=1'b0;
    defparam buf_cfgRTD_i0_LC_8_10_4.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i0_LC_8_10_4.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_cfgRTD_i0_LC_8_10_4 (
            .in0(N__52189),
            .in1(N__45328),
            .in2(N__43504),
            .in3(N__23718),
            .lcout(buf_cfgRTD_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55114),
            .ce(),
            .sr(_gnd_net_));
    defparam i12100_2_lut_LC_8_10_5.C_ON=1'b0;
    defparam i12100_2_lut_LC_8_10_5.SEQ_MODE=4'b0000;
    defparam i12100_2_lut_LC_8_10_5.LUT_INIT=16'b0101010100000000;
    LogicCell40 i12100_2_lut_LC_8_10_5 (
            .in0(N__54721),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54091),
            .lcout(n14490),
            .ltout(n14490_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i1_LC_8_10_6.C_ON=1'b0;
    defparam comm_cmd_i1_LC_8_10_6.SEQ_MODE=4'b1000;
    defparam comm_cmd_i1_LC_8_10_6.LUT_INIT=16'b1100000010101010;
    LogicCell40 comm_cmd_i1_LC_8_10_6 (
            .in0(N__57346),
            .in1(N__35991),
            .in2(N__23701),
            .in3(N__30939),
            .lcout(comm_cmd_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55114),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19526_LC_8_10_7.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19526_LC_8_10_7.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19526_LC_8_10_7.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_0__bdd_4_lut_19526_LC_8_10_7 (
            .in0(N__23680),
            .in1(N__57341),
            .in2(N__23659),
            .in3(N__56884),
            .lcout(n22165),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_1_i22_3_lut_LC_8_11_0.C_ON=1'b0;
    defparam mux_130_Mux_1_i22_3_lut_LC_8_11_0.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_1_i22_3_lut_LC_8_11_0.LUT_INIT=16'b1110111001000100;
    LogicCell40 mux_130_Mux_1_i22_3_lut_LC_8_11_0 (
            .in0(N__47743),
            .in1(N__23629),
            .in2(_gnd_net_),
            .in3(N__23941),
            .lcout(),
            .ltout(n22_adj_1618_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_1_i30_3_lut_LC_8_11_1.C_ON=1'b0;
    defparam mux_130_Mux_1_i30_3_lut_LC_8_11_1.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_1_i30_3_lut_LC_8_11_1.LUT_INIT=16'b1100110011110000;
    LogicCell40 mux_130_Mux_1_i30_3_lut_LC_8_11_1 (
            .in0(_gnd_net_),
            .in1(N__23596),
            .in2(N__23584),
            .in3(N__56345),
            .lcout(n30_adj_1619),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18186_4_lut_LC_8_11_2.C_ON=1'b0;
    defparam i18186_4_lut_LC_8_11_2.SEQ_MODE=4'b0000;
    defparam i18186_4_lut_LC_8_11_2.LUT_INIT=16'b1111110110101000;
    LogicCell40 i18186_4_lut_LC_8_11_2 (
            .in0(N__57186),
            .in1(N__56685),
            .in2(N__24004),
            .in3(N__41449),
            .lcout(),
            .ltout(n20781_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_2__bdd_4_lut_19360_LC_8_11_3.C_ON=1'b0;
    defparam comm_cmd_2__bdd_4_lut_19360_LC_8_11_3.SEQ_MODE=4'b0000;
    defparam comm_cmd_2__bdd_4_lut_19360_LC_8_11_3.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_cmd_2__bdd_4_lut_19360_LC_8_11_3 (
            .in0(N__23932),
            .in1(N__47744),
            .in2(N__23989),
            .in3(N__56346),
            .lcout(n21943),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_1_i19_3_lut_LC_8_11_4.C_ON=1'b0;
    defparam mux_130_Mux_1_i19_3_lut_LC_8_11_4.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_1_i19_3_lut_LC_8_11_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_130_Mux_1_i19_3_lut_LC_8_11_4 (
            .in0(N__23986),
            .in1(N__23961),
            .in2(_gnd_net_),
            .in3(N__56684),
            .lcout(n19_adj_1617),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19536_LC_8_11_5.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19536_LC_8_11_5.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19536_LC_8_11_5.LUT_INIT=16'b1110010010101010;
    LogicCell40 comm_cmd_0__bdd_4_lut_19536_LC_8_11_5 (
            .in0(N__56683),
            .in1(N__41899),
            .in2(N__30463),
            .in3(N__57184),
            .lcout(),
            .ltout(n22171_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22171_bdd_4_lut_LC_8_11_6.C_ON=1'b0;
    defparam n22171_bdd_4_lut_LC_8_11_6.SEQ_MODE=4'b0000;
    defparam n22171_bdd_4_lut_LC_8_11_6.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22171_bdd_4_lut_LC_8_11_6 (
            .in0(N__57185),
            .in1(N__50299),
            .in2(N__23935),
            .in3(N__31537),
            .lcout(n20775),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15210_2_lut_3_lut_LC_8_12_0.C_ON=1'b0;
    defparam i15210_2_lut_3_lut_LC_8_12_0.SEQ_MODE=4'b0000;
    defparam i15210_2_lut_3_lut_LC_8_12_0.LUT_INIT=16'b0000000000100010;
    LogicCell40 i15210_2_lut_3_lut_LC_8_12_0 (
            .in0(N__30803),
            .in1(N__51284),
            .in2(_gnd_net_),
            .in3(N__54092),
            .lcout(n14_adj_1523),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_2__bdd_4_lut_19433_LC_8_12_2.C_ON=1'b0;
    defparam comm_cmd_2__bdd_4_lut_19433_LC_8_12_2.SEQ_MODE=4'b0000;
    defparam comm_cmd_2__bdd_4_lut_19433_LC_8_12_2.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_cmd_2__bdd_4_lut_19433_LC_8_12_2 (
            .in0(N__23923),
            .in1(N__47789),
            .in2(N__23911),
            .in3(N__56338),
            .lcout(),
            .ltout(n22051_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22051_bdd_4_lut_LC_8_12_3.C_ON=1'b0;
    defparam n22051_bdd_4_lut_LC_8_12_3.SEQ_MODE=4'b0000;
    defparam n22051_bdd_4_lut_LC_8_12_3.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22051_bdd_4_lut_LC_8_12_3 (
            .in0(N__56339),
            .in1(N__24205),
            .in2(N__23899),
            .in3(N__23896),
            .lcout(n22054),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n21967_bdd_4_lut_LC_8_12_5.C_ON=1'b0;
    defparam n21967_bdd_4_lut_LC_8_12_5.SEQ_MODE=4'b0000;
    defparam n21967_bdd_4_lut_LC_8_12_5.LUT_INIT=16'b1110111001010000;
    LogicCell40 n21967_bdd_4_lut_LC_8_12_5 (
            .in0(N__56340),
            .in1(N__23887),
            .in2(N__26008),
            .in3(N__25612),
            .lcout(n21970),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i25_LC_8_12_6 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i25_LC_8_12_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i25_LC_8_12_6 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i25_LC_8_12_6  (
            .in0(N__37869),
            .in1(N__24256),
            .in2(N__48280),
            .in3(N__24230),
            .lcout(cmd_rdadctmp_25_adj_1418),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55135),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i20_LC_8_12_7 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i20_LC_8_12_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i20_LC_8_12_7 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i20_LC_8_12_7  (
            .in0(N__24128),
            .in1(N__48219),
            .in2(N__24031),
            .in3(N__37868),
            .lcout(cmd_rdadctmp_20_adj_1423),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55135),
            .ce(),
            .sr(_gnd_net_));
    defparam n22039_bdd_4_lut_LC_8_13_0.C_ON=1'b0;
    defparam n22039_bdd_4_lut_LC_8_13_0.SEQ_MODE=4'b0000;
    defparam n22039_bdd_4_lut_LC_8_13_0.LUT_INIT=16'b1100110010111000;
    LogicCell40 n22039_bdd_4_lut_LC_8_13_0 (
            .in0(N__27613),
            .in1(N__24214),
            .in2(N__32272),
            .in3(N__57440),
            .lcout(n22042),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i7_LC_8_13_1.C_ON=1'b0;
    defparam buf_cfgRTD_i7_LC_8_13_1.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i7_LC_8_13_1.LUT_INIT=16'b1011101110001000;
    LogicCell40 buf_cfgRTD_i7_LC_8_13_1 (
            .in0(N__45727),
            .in1(N__45327),
            .in2(_gnd_net_),
            .in3(N__24166),
            .lcout(buf_cfgRTD_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55148),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i12_LC_8_13_2 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i12_LC_8_13_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i12_LC_8_13_2 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \ADC_VAC.ADC_DATA_i12_LC_8_13_2  (
            .in0(N__24090),
            .in1(N__48480),
            .in2(N__24138),
            .in3(N__48217),
            .lcout(buf_adcdata_vac_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55148),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i10_LC_8_13_3 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i10_LC_8_13_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i10_LC_8_13_3 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i10_LC_8_13_3  (
            .in0(N__48216),
            .in1(N__24112),
            .in2(N__48511),
            .in3(N__24045),
            .lcout(buf_adcdata_vac_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55148),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_4_i19_3_lut_LC_8_13_5.C_ON=1'b0;
    defparam mux_129_Mux_4_i19_3_lut_LC_8_13_5.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_4_i19_3_lut_LC_8_13_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_129_Mux_4_i19_3_lut_LC_8_13_5 (
            .in0(N__26734),
            .in1(N__24089),
            .in2(_gnd_net_),
            .in3(N__56725),
            .lcout(n19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_2_i19_3_lut_LC_8_13_7.C_ON=1'b0;
    defparam mux_129_Mux_2_i19_3_lut_LC_8_13_7.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_2_i19_3_lut_LC_8_13_7.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_129_Mux_2_i19_3_lut_LC_8_13_7 (
            .in0(N__24076),
            .in1(N__24044),
            .in2(_gnd_net_),
            .in3(N__56726),
            .lcout(n19_adj_1505),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i11_LC_8_14_0 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i11_LC_8_14_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i11_LC_8_14_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i11_LC_8_14_0  (
            .in0(N__48438),
            .in1(N__48218),
            .in2(N__24030),
            .in3(N__25893),
            .lcout(buf_adcdata_vac_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55163),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_7_i26_3_lut_LC_8_14_1.C_ON=1'b0;
    defparam mux_128_Mux_7_i26_3_lut_LC_8_14_1.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_7_i26_3_lut_LC_8_14_1.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_128_Mux_7_i26_3_lut_LC_8_14_1 (
            .in0(N__31306),
            .in1(N__56639),
            .in2(_gnd_net_),
            .in3(N__30100),
            .lcout(),
            .ltout(n26_adj_1511_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18239_4_lut_LC_8_14_2.C_ON=1'b0;
    defparam i18239_4_lut_LC_8_14_2.SEQ_MODE=4'b0000;
    defparam i18239_4_lut_LC_8_14_2.LUT_INIT=16'b0100010011110000;
    LogicCell40 i18239_4_lut_LC_8_14_2 (
            .in0(N__56641),
            .in1(N__24394),
            .in2(N__24376),
            .in3(N__57436),
            .lcout(),
            .ltout(n20834_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_2__bdd_4_lut_19442_LC_8_14_3.C_ON=1'b0;
    defparam comm_cmd_2__bdd_4_lut_19442_LC_8_14_3.SEQ_MODE=4'b0000;
    defparam comm_cmd_2__bdd_4_lut_19442_LC_8_14_3.LUT_INIT=16'b1111010110001000;
    LogicCell40 comm_cmd_2__bdd_4_lut_19442_LC_8_14_3 (
            .in0(N__56334),
            .in1(N__29032),
            .in2(N__24373),
            .in3(N__47753),
            .lcout(),
            .ltout(n22057_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22057_bdd_4_lut_LC_8_14_4.C_ON=1'b0;
    defparam n22057_bdd_4_lut_LC_8_14_4.SEQ_MODE=4'b0000;
    defparam n22057_bdd_4_lut_LC_8_14_4.LUT_INIT=16'b1111000011001010;
    LogicCell40 n22057_bdd_4_lut_LC_8_14_4 (
            .in0(N__27892),
            .in1(N__24292),
            .in2(N__24370),
            .in3(N__56335),
            .lcout(n22060),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19020_2_lut_LC_8_14_5.C_ON=1'b0;
    defparam i19020_2_lut_LC_8_14_5.SEQ_MODE=4'b0000;
    defparam i19020_2_lut_LC_8_14_5.LUT_INIT=16'b1111111111001100;
    LogicCell40 i19020_2_lut_LC_8_14_5 (
            .in0(_gnd_net_),
            .in1(N__24367),
            .in2(_gnd_net_),
            .in3(N__56640),
            .lcout(n21261),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22135_bdd_4_lut_LC_8_14_6.C_ON=1'b0;
    defparam n22135_bdd_4_lut_LC_8_14_6.SEQ_MODE=4'b0000;
    defparam n22135_bdd_4_lut_LC_8_14_6.LUT_INIT=16'b1010111010100100;
    LogicCell40 n22135_bdd_4_lut_LC_8_14_6 (
            .in0(N__24355),
            .in1(N__24342),
            .in2(N__57524),
            .in3(N__24310),
            .lcout(n20831),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i7_LC_8_15_0 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i7_LC_8_15_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i7_LC_8_15_0 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i7_LC_8_15_0  (
            .in0(N__50500),
            .in1(N__24279),
            .in2(N__24562),
            .in3(N__50921),
            .lcout(cmd_rdadctmp_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55178),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i21_LC_8_15_1 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i21_LC_8_15_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i21_LC_8_15_1 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i21_LC_8_15_1  (
            .in0(N__50919),
            .in1(N__48975),
            .in2(N__24646),
            .in3(N__27287),
            .lcout(buf_adcdata_iac_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55178),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_1_i16_3_lut_LC_8_15_3.C_ON=1'b0;
    defparam mux_129_Mux_1_i16_3_lut_LC_8_15_3.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_1_i16_3_lut_LC_8_15_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_129_Mux_1_i16_3_lut_LC_8_15_3 (
            .in0(N__31932),
            .in1(N__32239),
            .in2(_gnd_net_),
            .in3(N__56698),
            .lcout(n16_adj_1507),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i8_LC_8_15_4.C_ON=1'b0;
    defparam data_index_i8_LC_8_15_4.SEQ_MODE=4'b1000;
    defparam data_index_i8_LC_8_15_4.LUT_INIT=16'b0101110100001000;
    LogicCell40 data_index_i8_LC_8_15_4 (
            .in0(N__54718),
            .in1(N__24433),
            .in2(N__52167),
            .in3(N__42382),
            .lcout(data_index_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55178),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i6_LC_8_15_5 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i6_LC_8_15_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i6_LC_8_15_5 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i6_LC_8_15_5  (
            .in0(N__50920),
            .in1(N__24558),
            .in2(N__24718),
            .in3(N__50501),
            .lcout(cmd_rdadctmp_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55178),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_354_Mux_8_i15_4_lut_LC_8_15_6.C_ON=1'b0;
    defparam comm_state_3__I_0_354_Mux_8_i15_4_lut_LC_8_15_6.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_354_Mux_8_i15_4_lut_LC_8_15_6.LUT_INIT=16'b0101110100001000;
    LogicCell40 comm_state_3__I_0_354_Mux_8_i15_4_lut_LC_8_15_6 (
            .in0(N__54717),
            .in1(N__24432),
            .in2(N__52166),
            .in3(N__42381),
            .lcout(data_index_9_N_212_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_6__I_0_368_i8_2_lut_LC_8_15_7.C_ON=1'b0;
    defparam comm_cmd_6__I_0_368_i8_2_lut_LC_8_15_7.SEQ_MODE=4'b0000;
    defparam comm_cmd_6__I_0_368_i8_2_lut_LC_8_15_7.LUT_INIT=16'b1111111100110011;
    LogicCell40 comm_cmd_6__I_0_368_i8_2_lut_LC_8_15_7 (
            .in0(_gnd_net_),
            .in1(N__57388),
            .in2(_gnd_net_),
            .in3(N__47748),
            .lcout(n8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i19_LC_8_16_1 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i19_LC_8_16_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i19_LC_8_16_1 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i19_LC_8_16_1  (
            .in0(N__50759),
            .in1(N__48968),
            .in2(N__24616),
            .in3(N__26069),
            .lcout(buf_adcdata_iac_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55193),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i23_LC_8_16_3 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i23_LC_8_16_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i23_LC_8_16_3 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i23_LC_8_16_3  (
            .in0(N__50469),
            .in1(N__24454),
            .in2(N__50837),
            .in3(N__25856),
            .lcout(cmd_rdadctmp_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55193),
            .ce(),
            .sr(_gnd_net_));
    defparam i6362_3_lut_LC_8_16_5.C_ON=1'b0;
    defparam i6362_3_lut_LC_8_16_5.SEQ_MODE=4'b0000;
    defparam i6362_3_lut_LC_8_16_5.LUT_INIT=16'b1100110010101010;
    LogicCell40 i6362_3_lut_LC_8_16_5 (
            .in0(N__43487),
            .in1(N__42396),
            .in2(_gnd_net_),
            .in3(N__43300),
            .lcout(n8_adj_1534),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i7_LC_8_16_6.C_ON=1'b0;
    defparam data_index_i7_LC_8_16_6.SEQ_MODE=4'b1000;
    defparam data_index_i7_LC_8_16_6.LUT_INIT=16'b0101110100001000;
    LogicCell40 data_index_i7_LC_8_16_6 (
            .in0(N__54724),
            .in1(N__30078),
            .in2(N__52170),
            .in3(N__42439),
            .lcout(data_index_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55193),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i8_LC_8_17_0 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i8_LC_8_17_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i8_LC_8_17_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i8_LC_8_17_0  (
            .in0(N__50746),
            .in1(N__48894),
            .in2(N__45138),
            .in3(N__24413),
            .lcout(buf_adcdata_iac_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55207),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i27_LC_8_17_2 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i27_LC_8_17_2 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i27_LC_8_17_2 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i27_LC_8_17_2  (
            .in0(N__50415),
            .in1(N__27757),
            .in2(N__50834),
            .in3(N__24611),
            .lcout(cmd_rdadctmp_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55207),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i1_LC_8_17_3 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i1_LC_8_17_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i1_LC_8_17_3 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i1_LC_8_17_3  (
            .in0(N__24666),
            .in1(N__24574),
            .in2(N__50470),
            .in3(N__50749),
            .lcout(cmd_rdadctmp_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55207),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i5_LC_8_17_4 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i5_LC_8_17_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i5_LC_8_17_4 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i5_LC_8_17_4  (
            .in0(N__50417),
            .in1(N__24886),
            .in2(N__50836),
            .in3(N__24711),
            .lcout(cmd_rdadctmp_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55207),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i22_LC_8_17_5 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i22_LC_8_17_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i22_LC_8_17_5 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i22_LC_8_17_5  (
            .in0(N__48893),
            .in1(N__50747),
            .in2(N__24904),
            .in3(N__24683),
            .lcout(buf_adcdata_iac_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55207),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i2_LC_8_17_6 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i2_LC_8_17_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i2_LC_8_17_6 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i2_LC_8_17_6  (
            .in0(N__50416),
            .in1(N__24667),
            .in2(N__50835),
            .in3(N__24870),
            .lcout(cmd_rdadctmp_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55207),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i30_LC_8_17_7 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i30_LC_8_17_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i30_LC_8_17_7 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i30_LC_8_17_7  (
            .in0(N__24899),
            .in1(N__50748),
            .in2(N__24644),
            .in3(N__50418),
            .lcout(cmd_rdadctmp_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55207),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.CS_37_LC_8_18_0 .C_ON=1'b0;
    defparam \ADC_IAC.CS_37_LC_8_18_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.CS_37_LC_8_18_0 .LUT_INIT=16'b0101010001010101;
    LogicCell40 \ADC_IAC.CS_37_LC_8_18_0  (
            .in0(N__24820),
            .in1(N__50714),
            .in2(N__25012),
            .in3(N__24658),
            .lcout(IAC_CS),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55219),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i29_LC_8_18_1 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i29_LC_8_18_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i29_LC_8_18_1 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i29_LC_8_18_1  (
            .in0(N__50712),
            .in1(N__50458),
            .in2(N__24645),
            .in3(N__28157),
            .lcout(cmd_rdadctmp_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55219),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i28_LC_8_18_2 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i28_LC_8_18_2 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i28_LC_8_18_2 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i28_LC_8_18_2  (
            .in0(N__50454),
            .in1(N__50715),
            .in2(N__28161),
            .in3(N__24612),
            .lcout(cmd_rdadctmp_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55219),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i0_LC_8_18_3 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i0_LC_8_18_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i0_LC_8_18_3 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i0_LC_8_18_3  (
            .in0(N__50711),
            .in1(N__50457),
            .in2(N__24595),
            .in3(N__24573),
            .lcout(cmd_rdadctmp_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55219),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i31_LC_8_18_4 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i31_LC_8_18_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i31_LC_8_18_4 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i31_LC_8_18_4  (
            .in0(N__50455),
            .in1(N__50716),
            .in2(N__26292),
            .in3(N__24903),
            .lcout(cmd_rdadctmp_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55219),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i4_LC_8_18_5 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i4_LC_8_18_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i4_LC_8_18_5 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i4_LC_8_18_5  (
            .in0(N__50713),
            .in1(N__50459),
            .in2(N__24859),
            .in3(N__24885),
            .lcout(cmd_rdadctmp_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55219),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i3_LC_8_18_6 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i3_LC_8_18_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i3_LC_8_18_6 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i3_LC_8_18_6  (
            .in0(N__50456),
            .in1(N__24855),
            .in2(N__24874),
            .in3(N__50717),
            .lcout(cmd_rdadctmp_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55219),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_207_LC_8_18_7.C_ON=1'b0;
    defparam i1_4_lut_adj_207_LC_8_18_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_207_LC_8_18_7.LUT_INIT=16'b0000111100000110;
    LogicCell40 i1_4_lut_adj_207_LC_8_18_7 (
            .in0(N__50710),
            .in1(N__30005),
            .in2(N__24837),
            .in3(N__29936),
            .lcout(n14_adj_1581),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i1_2_lut_adj_5_LC_8_19_0 .C_ON=1'b0;
    defparam \ADC_IAC.i1_2_lut_adj_5_LC_8_19_0 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i1_2_lut_adj_5_LC_8_19_0 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \ADC_IAC.i1_2_lut_adj_5_LC_8_19_0  (
            .in0(_gnd_net_),
            .in1(N__29934),
            .in2(_gnd_net_),
            .in3(N__24814),
            .lcout(\ADC_IAC.n20670 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i1_4_lut_LC_8_19_1 .C_ON=1'b0;
    defparam \ADC_IAC.i1_4_lut_LC_8_19_1 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i1_4_lut_LC_8_19_1 .LUT_INIT=16'b1010101111101111;
    LogicCell40 \ADC_IAC.i1_4_lut_LC_8_19_1  (
            .in0(N__50649),
            .in1(N__30003),
            .in2(N__24997),
            .in3(N__30139),
            .lcout(\ADC_IAC.n20669 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i18158_4_lut_LC_8_19_2 .C_ON=1'b0;
    defparam \ADC_IAC.i18158_4_lut_LC_8_19_2 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i18158_4_lut_LC_8_19_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_IAC.i18158_4_lut_LC_8_19_2  (
            .in0(N__24807),
            .in1(N__24795),
            .in2(N__24784),
            .in3(N__24768),
            .lcout(),
            .ltout(\ADC_IAC.n20753_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i18170_4_lut_LC_8_19_3 .C_ON=1'b0;
    defparam \ADC_IAC.i18170_4_lut_LC_8_19_3 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i18170_4_lut_LC_8_19_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_IAC.i18170_4_lut_LC_8_19_3  (
            .in0(N__24756),
            .in1(N__24744),
            .in2(N__24733),
            .in3(N__24729),
            .lcout(),
            .ltout(\ADC_IAC.n20765_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i18788_4_lut_LC_8_19_4 .C_ON=1'b0;
    defparam \ADC_IAC.i18788_4_lut_LC_8_19_4 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i18788_4_lut_LC_8_19_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \ADC_IAC.i18788_4_lut_LC_8_19_4  (
            .in0(N__25042),
            .in1(N__50651),
            .in2(N__25027),
            .in3(N__29933),
            .lcout(),
            .ltout(\ADC_IAC.n21007_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.adc_state_i0_LC_8_19_5 .C_ON=1'b0;
    defparam \ADC_IAC.adc_state_i0_LC_8_19_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.adc_state_i0_LC_8_19_5 .LUT_INIT=16'b0001000111110000;
    LogicCell40 \ADC_IAC.adc_state_i0_LC_8_19_5  (
            .in0(N__29935),
            .in1(N__50724),
            .in2(N__25024),
            .in3(N__30004),
            .lcout(adc_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55230),
            .ce(N__25021),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i30_4_lut_LC_8_19_6 .C_ON=1'b0;
    defparam \ADC_IAC.i30_4_lut_LC_8_19_6 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i30_4_lut_LC_8_19_6 .LUT_INIT=16'b1010110000000101;
    LogicCell40 \ADC_IAC.i30_4_lut_LC_8_19_6  (
            .in0(N__30140),
            .in1(N__24989),
            .in2(N__30014),
            .in3(N__29932),
            .lcout(),
            .ltout(\ADC_IAC.n17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i19104_2_lut_LC_8_19_7 .C_ON=1'b0;
    defparam \ADC_IAC.i19104_2_lut_LC_8_19_7 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i19104_2_lut_LC_8_19_7 .LUT_INIT=16'b1010111110101111;
    LogicCell40 \ADC_IAC.i19104_2_lut_LC_8_19_7  (
            .in0(N__50650),
            .in1(_gnd_net_),
            .in2(N__24958),
            .in3(_gnd_net_),
            .lcout(\ADC_IAC.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i23_LC_9_4_2 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i23_LC_9_4_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i23_LC_9_4_2 .LUT_INIT=16'b1110001000101110;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i23_LC_9_4_2  (
            .in0(N__25429),
            .in1(N__34121),
            .in2(N__25401),
            .in3(N__26308),
            .lcout(\ADC_VDC.cmd_rdadctmp_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32806),
            .ce(N__26545),
            .sr(N__24946));
    defparam \comm_spi.RESET_I_0_102_2_lut_LC_9_4_5 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_102_2_lut_LC_9_4_5 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_102_2_lut_LC_9_4_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \comm_spi.RESET_I_0_102_2_lut_LC_9_4_5  (
            .in0(_gnd_net_),
            .in1(N__48744),
            .in2(_gnd_net_),
            .in3(N__55474),
            .lcout(\comm_spi.data_tx_7__N_772 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadcbuf_i0_LC_9_5_0 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i0_LC_9_5_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i0_LC_9_5_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i0_LC_9_5_0  (
            .in0(_gnd_net_),
            .in1(N__24931),
            .in2(N__26611),
            .in3(_gnd_net_),
            .lcout(\ADC_VDC.cmd_rdadcbuf_0 ),
            .ltout(),
            .carryin(bfn_9_5_0_),
            .carryout(\ADC_VDC.n19364 ),
            .clk(N__32842),
            .ce(N__29162),
            .sr(N__29103));
    defparam \ADC_VDC.cmd_rdadcbuf_i1_LC_9_5_1 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i1_LC_9_5_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i1_LC_9_5_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i1_LC_9_5_1  (
            .in0(_gnd_net_),
            .in1(N__24925),
            .in2(N__26410),
            .in3(N__24919),
            .lcout(\ADC_VDC.cmd_rdadcbuf_1 ),
            .ltout(),
            .carryin(\ADC_VDC.n19364 ),
            .carryout(\ADC_VDC.n19365 ),
            .clk(N__32842),
            .ce(N__29162),
            .sr(N__29103));
    defparam \ADC_VDC.cmd_rdadcbuf_i2_LC_9_5_2 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i2_LC_9_5_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i2_LC_9_5_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i2_LC_9_5_2  (
            .in0(_gnd_net_),
            .in1(N__26388),
            .in2(N__24916),
            .in3(N__24907),
            .lcout(\ADC_VDC.cmd_rdadcbuf_2 ),
            .ltout(),
            .carryin(\ADC_VDC.n19365 ),
            .carryout(\ADC_VDC.n19366 ),
            .clk(N__32842),
            .ce(N__29162),
            .sr(N__29103));
    defparam \ADC_VDC.cmd_rdadcbuf_i3_LC_9_5_3 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i3_LC_9_5_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i3_LC_9_5_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i3_LC_9_5_3  (
            .in0(_gnd_net_),
            .in1(N__25168),
            .in2(N__26590),
            .in3(N__25162),
            .lcout(\ADC_VDC.cmd_rdadcbuf_3 ),
            .ltout(),
            .carryin(\ADC_VDC.n19366 ),
            .carryout(\ADC_VDC.n19367 ),
            .clk(N__32842),
            .ce(N__29162),
            .sr(N__29103));
    defparam \ADC_VDC.cmd_rdadcbuf_i4_LC_9_5_4 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i4_LC_9_5_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i4_LC_9_5_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i4_LC_9_5_4  (
            .in0(_gnd_net_),
            .in1(N__25159),
            .in2(N__26568),
            .in3(N__25153),
            .lcout(\ADC_VDC.cmd_rdadcbuf_4 ),
            .ltout(),
            .carryin(\ADC_VDC.n19367 ),
            .carryout(\ADC_VDC.n19368 ),
            .clk(N__32842),
            .ce(N__29162),
            .sr(N__29103));
    defparam \ADC_VDC.cmd_rdadcbuf_i5_LC_9_5_5 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i5_LC_9_5_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i5_LC_9_5_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i5_LC_9_5_5  (
            .in0(_gnd_net_),
            .in1(N__25132),
            .in2(N__25150),
            .in3(N__25126),
            .lcout(\ADC_VDC.cmd_rdadcbuf_5 ),
            .ltout(),
            .carryin(\ADC_VDC.n19368 ),
            .carryout(\ADC_VDC.n19369 ),
            .clk(N__32842),
            .ce(N__29162),
            .sr(N__29103));
    defparam \ADC_VDC.cmd_rdadcbuf_i6_LC_9_5_6 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i6_LC_9_5_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i6_LC_9_5_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i6_LC_9_5_6  (
            .in0(_gnd_net_),
            .in1(N__25105),
            .in2(N__25123),
            .in3(N__25099),
            .lcout(\ADC_VDC.cmd_rdadcbuf_6 ),
            .ltout(),
            .carryin(\ADC_VDC.n19369 ),
            .carryout(\ADC_VDC.n19370 ),
            .clk(N__32842),
            .ce(N__29162),
            .sr(N__29103));
    defparam \ADC_VDC.cmd_rdadcbuf_i7_LC_9_5_7 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i7_LC_9_5_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i7_LC_9_5_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i7_LC_9_5_7  (
            .in0(_gnd_net_),
            .in1(N__25096),
            .in2(N__26533),
            .in3(N__25090),
            .lcout(\ADC_VDC.cmd_rdadcbuf_7 ),
            .ltout(),
            .carryin(\ADC_VDC.n19370 ),
            .carryout(\ADC_VDC.n19371 ),
            .clk(N__32842),
            .ce(N__29162),
            .sr(N__29103));
    defparam \ADC_VDC.cmd_rdadcbuf_i8_LC_9_6_0 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i8_LC_9_6_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i8_LC_9_6_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i8_LC_9_6_0  (
            .in0(_gnd_net_),
            .in1(N__25087),
            .in2(N__26508),
            .in3(N__25081),
            .lcout(\ADC_VDC.cmd_rdadcbuf_8 ),
            .ltout(),
            .carryin(bfn_9_6_0_),
            .carryout(\ADC_VDC.n19372 ),
            .clk(N__32903),
            .ce(N__29179),
            .sr(N__29108));
    defparam \ADC_VDC.cmd_rdadcbuf_i9_LC_9_6_1 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i9_LC_9_6_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i9_LC_9_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i9_LC_9_6_1  (
            .in0(_gnd_net_),
            .in1(N__25076),
            .in2(N__25063),
            .in3(N__25054),
            .lcout(\ADC_VDC.cmd_rdadcbuf_9 ),
            .ltout(),
            .carryin(\ADC_VDC.n19372 ),
            .carryout(\ADC_VDC.n19373 ),
            .clk(N__32903),
            .ce(N__29179),
            .sr(N__29108));
    defparam \ADC_VDC.cmd_rdadcbuf_i10_LC_9_6_2 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i10_LC_9_6_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i10_LC_9_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i10_LC_9_6_2  (
            .in0(_gnd_net_),
            .in1(N__25051),
            .in2(N__26984),
            .in3(N__25045),
            .lcout(\ADC_VDC.cmd_rdadcbuf_10 ),
            .ltout(),
            .carryin(\ADC_VDC.n19373 ),
            .carryout(\ADC_VDC.n19374 ),
            .clk(N__32903),
            .ce(N__29179),
            .sr(N__29108));
    defparam \ADC_VDC.cmd_rdadcbuf_i11_LC_9_6_3 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i11_LC_9_6_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i11_LC_9_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i11_LC_9_6_3  (
            .in0(_gnd_net_),
            .in1(N__25317),
            .in2(N__26959),
            .in3(N__25306),
            .lcout(cmd_rdadcbuf_11),
            .ltout(),
            .carryin(\ADC_VDC.n19374 ),
            .carryout(\ADC_VDC.n19375 ),
            .clk(N__32903),
            .ce(N__29179),
            .sr(N__29108));
    defparam \ADC_VDC.cmd_rdadcbuf_i12_LC_9_6_4 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i12_LC_9_6_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i12_LC_9_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i12_LC_9_6_4  (
            .in0(_gnd_net_),
            .in1(N__25302),
            .in2(N__26365),
            .in3(N__25291),
            .lcout(cmd_rdadcbuf_12),
            .ltout(),
            .carryin(\ADC_VDC.n19375 ),
            .carryout(\ADC_VDC.n19376 ),
            .clk(N__32903),
            .ce(N__29179),
            .sr(N__29108));
    defparam \ADC_VDC.cmd_rdadcbuf_i13_LC_9_6_5 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i13_LC_9_6_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i13_LC_9_6_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i13_LC_9_6_5  (
            .in0(_gnd_net_),
            .in1(N__25266),
            .in2(N__25288),
            .in3(N__25255),
            .lcout(cmd_rdadcbuf_13),
            .ltout(),
            .carryin(\ADC_VDC.n19376 ),
            .carryout(\ADC_VDC.n19377 ),
            .clk(N__32903),
            .ce(N__29179),
            .sr(N__29108));
    defparam \ADC_VDC.cmd_rdadcbuf_i14_LC_9_6_6 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i14_LC_9_6_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i14_LC_9_6_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i14_LC_9_6_6  (
            .in0(_gnd_net_),
            .in1(N__25221),
            .in2(N__25247),
            .in3(N__25210),
            .lcout(cmd_rdadcbuf_14),
            .ltout(),
            .carryin(\ADC_VDC.n19377 ),
            .carryout(\ADC_VDC.n19378 ),
            .clk(N__32903),
            .ce(N__29179),
            .sr(N__29108));
    defparam \ADC_VDC.cmd_rdadcbuf_i15_LC_9_6_7 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i15_LC_9_6_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i15_LC_9_6_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i15_LC_9_6_7  (
            .in0(_gnd_net_),
            .in1(N__26670),
            .in2(N__26451),
            .in3(N__25207),
            .lcout(cmd_rdadcbuf_15),
            .ltout(),
            .carryin(\ADC_VDC.n19378 ),
            .carryout(\ADC_VDC.n19379 ),
            .clk(N__32903),
            .ce(N__29179),
            .sr(N__29108));
    defparam \ADC_VDC.cmd_rdadcbuf_i16_LC_9_7_0 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i16_LC_9_7_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i16_LC_9_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i16_LC_9_7_0  (
            .in0(_gnd_net_),
            .in1(N__27087),
            .in2(N__26428),
            .in3(N__25204),
            .lcout(cmd_rdadcbuf_16),
            .ltout(),
            .carryin(bfn_9_7_0_),
            .carryout(\ADC_VDC.n19380 ),
            .clk(N__32896),
            .ce(N__29191),
            .sr(N__29104));
    defparam \ADC_VDC.cmd_rdadcbuf_i17_LC_9_7_1 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i17_LC_9_7_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i17_LC_9_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i17_LC_9_7_1  (
            .in0(_gnd_net_),
            .in1(N__27102),
            .in2(N__26481),
            .in3(N__25201),
            .lcout(cmd_rdadcbuf_17),
            .ltout(),
            .carryin(\ADC_VDC.n19380 ),
            .carryout(\ADC_VDC.n19381 ),
            .clk(N__32896),
            .ce(N__29191),
            .sr(N__29104));
    defparam \ADC_VDC.cmd_rdadcbuf_i18_LC_9_7_2 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i18_LC_9_7_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i18_LC_9_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i18_LC_9_7_2  (
            .in0(_gnd_net_),
            .in1(N__27114),
            .in2(N__25197),
            .in3(N__25174),
            .lcout(cmd_rdadcbuf_18),
            .ltout(),
            .carryin(\ADC_VDC.n19381 ),
            .carryout(\ADC_VDC.n19382 ),
            .clk(N__32896),
            .ce(N__29191),
            .sr(N__29104));
    defparam \ADC_VDC.cmd_rdadcbuf_i19_LC_9_7_3 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i19_LC_9_7_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i19_LC_9_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i19_LC_9_7_3  (
            .in0(_gnd_net_),
            .in1(N__26646),
            .in2(N__26919),
            .in3(N__25171),
            .lcout(cmd_rdadcbuf_19),
            .ltout(),
            .carryin(\ADC_VDC.n19382 ),
            .carryout(\ADC_VDC.n19383 ),
            .clk(N__32896),
            .ce(N__29191),
            .sr(N__29104));
    defparam \ADC_VDC.cmd_rdadcbuf_i20_LC_9_7_4 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i20_LC_9_7_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i20_LC_9_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i20_LC_9_7_4  (
            .in0(_gnd_net_),
            .in1(N__26658),
            .in2(N__26769),
            .in3(N__25468),
            .lcout(cmd_rdadcbuf_20),
            .ltout(),
            .carryin(\ADC_VDC.n19383 ),
            .carryout(\ADC_VDC.n19384 ),
            .clk(N__32896),
            .ce(N__29191),
            .sr(N__29104));
    defparam \ADC_VDC.cmd_rdadcbuf_i21_LC_9_7_5 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i21_LC_9_7_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i21_LC_9_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i21_LC_9_7_5  (
            .in0(_gnd_net_),
            .in1(N__25443),
            .in2(N__25465),
            .in3(N__25432),
            .lcout(cmd_rdadcbuf_21),
            .ltout(),
            .carryin(\ADC_VDC.n19384 ),
            .carryout(\ADC_VDC.n19385 ),
            .clk(N__32896),
            .ce(N__29191),
            .sr(N__29104));
    defparam \ADC_VDC.cmd_rdadcbuf_i22_LC_9_7_6 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i22_LC_9_7_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i22_LC_9_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i22_LC_9_7_6  (
            .in0(_gnd_net_),
            .in1(N__26709),
            .in2(N__25428),
            .in3(N__25405),
            .lcout(cmd_rdadcbuf_22),
            .ltout(),
            .carryin(\ADC_VDC.n19385 ),
            .carryout(\ADC_VDC.n19386 ),
            .clk(N__32896),
            .ce(N__29191),
            .sr(N__29104));
    defparam \ADC_VDC.cmd_rdadcbuf_i23_LC_9_7_7 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i23_LC_9_7_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i23_LC_9_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i23_LC_9_7_7  (
            .in0(_gnd_net_),
            .in1(N__26745),
            .in2(N__25402),
            .in3(N__25381),
            .lcout(cmd_rdadcbuf_23),
            .ltout(),
            .carryin(\ADC_VDC.n19386 ),
            .carryout(\ADC_VDC.n19387 ),
            .clk(N__32896),
            .ce(N__29191),
            .sr(N__29104));
    defparam \ADC_VDC.cmd_rdadcbuf_i24_LC_9_8_0 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i24_LC_9_8_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i24_LC_9_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i24_LC_9_8_0  (
            .in0(_gnd_net_),
            .in1(N__25377),
            .in2(_gnd_net_),
            .in3(N__25366),
            .lcout(cmd_rdadcbuf_24),
            .ltout(),
            .carryin(bfn_9_8_0_),
            .carryout(\ADC_VDC.n19388 ),
            .clk(N__32894),
            .ce(N__29186),
            .sr(N__29113));
    defparam \ADC_VDC.cmd_rdadcbuf_i25_LC_9_8_1 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i25_LC_9_8_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i25_LC_9_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i25_LC_9_8_1  (
            .in0(_gnd_net_),
            .in1(N__25362),
            .in2(_gnd_net_),
            .in3(N__25351),
            .lcout(cmd_rdadcbuf_25),
            .ltout(),
            .carryin(\ADC_VDC.n19388 ),
            .carryout(\ADC_VDC.n19389 ),
            .clk(N__32894),
            .ce(N__29186),
            .sr(N__29113));
    defparam \ADC_VDC.cmd_rdadcbuf_i26_LC_9_8_2 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i26_LC_9_8_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i26_LC_9_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i26_LC_9_8_2  (
            .in0(_gnd_net_),
            .in1(N__25347),
            .in2(_gnd_net_),
            .in3(N__25336),
            .lcout(cmd_rdadcbuf_26),
            .ltout(),
            .carryin(\ADC_VDC.n19389 ),
            .carryout(\ADC_VDC.n19390 ),
            .clk(N__32894),
            .ce(N__29186),
            .sr(N__29113));
    defparam \ADC_VDC.cmd_rdadcbuf_i27_LC_9_8_3 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i27_LC_9_8_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i27_LC_9_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i27_LC_9_8_3  (
            .in0(_gnd_net_),
            .in1(N__25332),
            .in2(_gnd_net_),
            .in3(N__25321),
            .lcout(cmd_rdadcbuf_27),
            .ltout(),
            .carryin(\ADC_VDC.n19390 ),
            .carryout(\ADC_VDC.n19391 ),
            .clk(N__32894),
            .ce(N__29186),
            .sr(N__29113));
    defparam \ADC_VDC.cmd_rdadcbuf_i28_LC_9_8_4 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i28_LC_9_8_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i28_LC_9_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i28_LC_9_8_4  (
            .in0(_gnd_net_),
            .in1(N__25578),
            .in2(_gnd_net_),
            .in3(N__25567),
            .lcout(cmd_rdadcbuf_28),
            .ltout(),
            .carryin(\ADC_VDC.n19391 ),
            .carryout(\ADC_VDC.n19392 ),
            .clk(N__32894),
            .ce(N__29186),
            .sr(N__29113));
    defparam \ADC_VDC.cmd_rdadcbuf_i29_LC_9_8_5 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i29_LC_9_8_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i29_LC_9_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i29_LC_9_8_5  (
            .in0(_gnd_net_),
            .in1(N__25563),
            .in2(_gnd_net_),
            .in3(N__25552),
            .lcout(cmd_rdadcbuf_29),
            .ltout(),
            .carryin(\ADC_VDC.n19392 ),
            .carryout(\ADC_VDC.n19393 ),
            .clk(N__32894),
            .ce(N__29186),
            .sr(N__29113));
    defparam \ADC_VDC.cmd_rdadcbuf_i30_LC_9_8_6 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i30_LC_9_8_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i30_LC_9_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i30_LC_9_8_6  (
            .in0(_gnd_net_),
            .in1(N__25548),
            .in2(_gnd_net_),
            .in3(N__25537),
            .lcout(cmd_rdadcbuf_30),
            .ltout(),
            .carryin(\ADC_VDC.n19393 ),
            .carryout(\ADC_VDC.n19394 ),
            .clk(N__32894),
            .ce(N__29186),
            .sr(N__29113));
    defparam \ADC_VDC.cmd_rdadcbuf_i31_LC_9_8_7 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i31_LC_9_8_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i31_LC_9_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i31_LC_9_8_7  (
            .in0(_gnd_net_),
            .in1(N__25533),
            .in2(_gnd_net_),
            .in3(N__25522),
            .lcout(cmd_rdadcbuf_31),
            .ltout(),
            .carryin(\ADC_VDC.n19394 ),
            .carryout(\ADC_VDC.n19395 ),
            .clk(N__32894),
            .ce(N__29186),
            .sr(N__29113));
    defparam \ADC_VDC.cmd_rdadcbuf_i32_LC_9_9_0 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i32_LC_9_9_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i32_LC_9_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i32_LC_9_9_0  (
            .in0(_gnd_net_),
            .in1(N__25518),
            .in2(_gnd_net_),
            .in3(N__25507),
            .lcout(cmd_rdadcbuf_32),
            .ltout(),
            .carryin(bfn_9_9_0_),
            .carryout(\ADC_VDC.n19396 ),
            .clk(N__32884),
            .ce(N__29190),
            .sr(N__29109));
    defparam \ADC_VDC.cmd_rdadcbuf_i33_LC_9_9_1 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i33_LC_9_9_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i33_LC_9_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i33_LC_9_9_1  (
            .in0(_gnd_net_),
            .in1(N__25503),
            .in2(_gnd_net_),
            .in3(N__25492),
            .lcout(cmd_rdadcbuf_33),
            .ltout(),
            .carryin(\ADC_VDC.n19396 ),
            .carryout(\ADC_VDC.n19397 ),
            .clk(N__32884),
            .ce(N__29190),
            .sr(N__29109));
    defparam \ADC_VDC.add_23_36_lut_LC_9_9_2 .C_ON=1'b0;
    defparam \ADC_VDC.add_23_36_lut_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.add_23_36_lut_LC_9_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.add_23_36_lut_LC_9_9_2  (
            .in0(_gnd_net_),
            .in1(N__27047),
            .in2(_gnd_net_),
            .in3(N__25489),
            .lcout(\ADC_VDC.cmd_rdadcbuf_35_N_1130_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n21943_bdd_4_lut_LC_9_10_0.C_ON=1'b0;
    defparam n21943_bdd_4_lut_LC_9_10_0.SEQ_MODE=4'b0000;
    defparam n21943_bdd_4_lut_LC_9_10_0.LUT_INIT=16'b1110111001010000;
    LogicCell40 n21943_bdd_4_lut_LC_9_10_0 (
            .in0(N__56272),
            .in1(N__25486),
            .in2(N__27940),
            .in3(N__25477),
            .lcout(),
            .ltout(n21946_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_0__i0_LC_9_10_1.C_ON=1'b0;
    defparam comm_buf_0__i0_LC_9_10_1.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i0_LC_9_10_1.LUT_INIT=16'b1111101001010000;
    LogicCell40 comm_buf_0__i0_LC_9_10_1 (
            .in0(N__54099),
            .in1(_gnd_net_),
            .in2(N__25471),
            .in3(N__36255),
            .lcout(comm_buf_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55104),
            .ce(N__27504),
            .sr(N__27453));
    defparam i15211_2_lut_3_lut_LC_9_10_2.C_ON=1'b0;
    defparam i15211_2_lut_3_lut_LC_9_10_2.SEQ_MODE=4'b0000;
    defparam i15211_2_lut_3_lut_LC_9_10_2.LUT_INIT=16'b0000000000100010;
    LogicCell40 i15211_2_lut_3_lut_LC_9_10_2 (
            .in0(N__43461),
            .in1(N__51219),
            .in2(_gnd_net_),
            .in3(N__54097),
            .lcout(n14_adj_1524),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15203_2_lut_3_lut_LC_9_10_4.C_ON=1'b0;
    defparam i15203_2_lut_3_lut_LC_9_10_4.SEQ_MODE=4'b0000;
    defparam i15203_2_lut_3_lut_LC_9_10_4.LUT_INIT=16'b0000000000100010;
    LogicCell40 i15203_2_lut_3_lut_LC_9_10_4 (
            .in0(N__38650),
            .in1(N__51218),
            .in2(_gnd_net_),
            .in3(N__54096),
            .lcout(n14_adj_1551),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15205_2_lut_3_lut_LC_9_10_6.C_ON=1'b0;
    defparam i15205_2_lut_3_lut_LC_9_10_6.SEQ_MODE=4'b0000;
    defparam i15205_2_lut_3_lut_LC_9_10_6.LUT_INIT=16'b0000000000100010;
    LogicCell40 i15205_2_lut_3_lut_LC_9_10_6 (
            .in0(N__42623),
            .in1(N__51220),
            .in2(_gnd_net_),
            .in3(N__54098),
            .lcout(n14_adj_1525),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_0__i7_LC_9_11_0.C_ON=1'b0;
    defparam comm_buf_0__i7_LC_9_11_0.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i7_LC_9_11_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_0__i7_LC_9_11_0 (
            .in0(N__54103),
            .in1(N__36896),
            .in2(_gnd_net_),
            .in3(N__25597),
            .lcout(comm_buf_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55115),
            .ce(N__27512),
            .sr(N__27465));
    defparam comm_buf_0__i6_LC_9_11_1.C_ON=1'b0;
    defparam comm_buf_0__i6_LC_9_11_1.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i6_LC_9_11_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_0__i6_LC_9_11_1 (
            .in0(N__35810),
            .in1(N__25588),
            .in2(_gnd_net_),
            .in3(N__54105),
            .lcout(comm_buf_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55115),
            .ce(N__27512),
            .sr(N__27465));
    defparam comm_buf_0__i4_LC_9_11_2.C_ON=1'b0;
    defparam comm_buf_0__i4_LC_9_11_2.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i4_LC_9_11_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_0__i4_LC_9_11_2 (
            .in0(N__54102),
            .in1(N__35668),
            .in2(_gnd_net_),
            .in3(N__25720),
            .lcout(comm_buf_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55115),
            .ce(N__27512),
            .sr(N__27465));
    defparam comm_buf_0__i3_LC_9_11_3.C_ON=1'b0;
    defparam comm_buf_0__i3_LC_9_11_3.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i3_LC_9_11_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 comm_buf_0__i3_LC_9_11_3 (
            .in0(N__35563),
            .in1(N__54104),
            .in2(_gnd_net_),
            .in3(N__41230),
            .lcout(comm_buf_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55115),
            .ce(N__27512),
            .sr(N__27465));
    defparam comm_cmd_0__bdd_4_lut_19413_LC_9_12_1.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19413_LC_9_12_1.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19413_LC_9_12_1.LUT_INIT=16'b1101100010101010;
    LogicCell40 comm_cmd_0__bdd_4_lut_19413_LC_9_12_1 (
            .in0(N__56562),
            .in1(N__38936),
            .in2(N__41656),
            .in3(N__57443),
            .lcout(),
            .ltout(n22015_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22015_bdd_4_lut_LC_9_12_2.C_ON=1'b0;
    defparam n22015_bdd_4_lut_LC_9_12_2.SEQ_MODE=4'b0000;
    defparam n22015_bdd_4_lut_LC_9_12_2.LUT_INIT=16'b1111001011000010;
    LogicCell40 n22015_bdd_4_lut_LC_9_12_2 (
            .in0(N__44031),
            .in1(N__57444),
            .in2(N__25582),
            .in3(N__36925),
            .lcout(n20871),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18223_3_lut_LC_9_12_3.C_ON=1'b0;
    defparam i18223_3_lut_LC_9_12_3.SEQ_MODE=4'b0000;
    defparam i18223_3_lut_LC_9_12_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 i18223_3_lut_LC_9_12_3 (
            .in0(N__56563),
            .in1(N__31198),
            .in2(_gnd_net_),
            .in3(N__47311),
            .lcout(),
            .ltout(n20818_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18225_4_lut_LC_9_12_4.C_ON=1'b0;
    defparam i18225_4_lut_LC_9_12_4.SEQ_MODE=4'b0000;
    defparam i18225_4_lut_LC_9_12_4.LUT_INIT=16'b1111110010111000;
    LogicCell40 i18225_4_lut_LC_9_12_4 (
            .in0(N__25639),
            .in1(N__57445),
            .in2(N__25624),
            .in3(N__56567),
            .lcout(),
            .ltout(n20820_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_2__bdd_4_lut_19408_LC_9_12_5.C_ON=1'b0;
    defparam comm_cmd_2__bdd_4_lut_19408_LC_9_12_5.SEQ_MODE=4'b0000;
    defparam comm_cmd_2__bdd_4_lut_19408_LC_9_12_5.LUT_INIT=16'b1111010110001000;
    LogicCell40 comm_cmd_2__bdd_4_lut_19408_LC_9_12_5 (
            .in0(N__56344),
            .in1(N__25621),
            .in2(N__25615),
            .in3(N__47746),
            .lcout(n21967),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_0__i1_LC_9_12_6.C_ON=1'b0;
    defparam comm_buf_0__i1_LC_9_12_6.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i1_LC_9_12_6.LUT_INIT=16'b1011101110001000;
    LogicCell40 comm_buf_0__i1_LC_9_12_6 (
            .in0(N__35995),
            .in1(N__54106),
            .in2(_gnd_net_),
            .in3(N__25606),
            .lcout(comm_buf_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55124),
            .ce(N__27517),
            .sr(N__27469));
    defparam i36_4_lut_4_lut_LC_9_12_7.C_ON=1'b0;
    defparam i36_4_lut_4_lut_LC_9_12_7.SEQ_MODE=4'b0000;
    defparam i36_4_lut_4_lut_LC_9_12_7.LUT_INIT=16'b0010010010101110;
    LogicCell40 i36_4_lut_4_lut_LC_9_12_7 (
            .in0(N__56343),
            .in1(N__57442),
            .in2(N__56699),
            .in3(N__47745),
            .lcout(n30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19398_LC_9_13_0.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19398_LC_9_13_0.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19398_LC_9_13_0.LUT_INIT=16'b1110010010101010;
    LogicCell40 comm_cmd_0__bdd_4_lut_19398_LC_9_13_0 (
            .in0(N__56635),
            .in1(N__26100),
            .in2(N__28134),
            .in3(N__57242),
            .lcout(),
            .ltout(n22003_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22003_bdd_4_lut_LC_9_13_1.C_ON=1'b0;
    defparam n22003_bdd_4_lut_LC_9_13_1.SEQ_MODE=4'b0000;
    defparam n22003_bdd_4_lut_LC_9_13_1.LUT_INIT=16'b1110001111100000;
    LogicCell40 n22003_bdd_4_lut_LC_9_13_1 (
            .in0(N__27587),
            .in1(N__57250),
            .in2(N__25600),
            .in3(N__33864),
            .lcout(n22006),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i24_LC_9_13_2 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i24_LC_9_13_2 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i24_LC_9_13_2 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i24_LC_9_13_2  (
            .in0(N__50512),
            .in1(N__25982),
            .in2(N__25873),
            .in3(N__50882),
            .lcout(cmd_rdadctmp_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55136),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i0_LC_9_13_3.C_ON=1'b0;
    defparam comm_cmd_i0_LC_9_13_3.SEQ_MODE=4'b1000;
    defparam comm_cmd_i0_LC_9_13_3.LUT_INIT=16'b1110010001000100;
    LogicCell40 comm_cmd_i0_LC_9_13_3 (
            .in0(N__30943),
            .in1(N__56637),
            .in2(N__30993),
            .in3(N__36259),
            .lcout(comm_cmd_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55136),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_4_lut_adj_101_LC_9_13_4.C_ON=1'b0;
    defparam i1_2_lut_4_lut_adj_101_LC_9_13_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_4_lut_adj_101_LC_9_13_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_2_lut_4_lut_adj_101_LC_9_13_4 (
            .in0(N__56636),
            .in1(N__57241),
            .in2(N__45381),
            .in3(N__47747),
            .lcout(n20624),
            .ltout(n20624_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_90_LC_9_13_5.C_ON=1'b0;
    defparam i1_4_lut_adj_90_LC_9_13_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_90_LC_9_13_5.LUT_INIT=16'b1100111101000101;
    LogicCell40 i1_4_lut_adj_90_LC_9_13_5 (
            .in0(N__52168),
            .in1(N__49239),
            .in2(N__25765),
            .in3(N__54722),
            .lcout(n11417),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19057_2_lut_LC_9_13_7.C_ON=1'b0;
    defparam i19057_2_lut_LC_9_13_7.SEQ_MODE=4'b0000;
    defparam i19057_2_lut_LC_9_13_7.LUT_INIT=16'b1010101000000000;
    LogicCell40 i19057_2_lut_LC_9_13_7 (
            .in0(N__31357),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56634),
            .lcout(n20936),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.i4_4_lut_LC_9_14_0 .C_ON=1'b0;
    defparam \SIG_DDS.i4_4_lut_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \SIG_DDS.i4_4_lut_LC_9_14_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \SIG_DDS.i4_4_lut_LC_9_14_0  (
            .in0(N__55695),
            .in1(N__25910),
            .in2(N__25937),
            .in3(N__43677),
            .lcout(),
            .ltout(\SIG_DDS.n10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.dds_state_i0_LC_9_14_1 .C_ON=1'b0;
    defparam \SIG_DDS.dds_state_i0_LC_9_14_1 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.dds_state_i0_LC_9_14_1 .LUT_INIT=16'b1000000010110011;
    LogicCell40 \SIG_DDS.dds_state_i0_LC_9_14_1  (
            .in0(N__25774),
            .in1(N__55655),
            .in2(N__25762),
            .in3(N__55696),
            .lcout(dds_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55149),
            .ce(N__45538),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_LC_9_14_2.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_LC_9_14_2.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_LC_9_14_2.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_0__bdd_4_lut_LC_9_14_2 (
            .in0(N__42045),
            .in1(N__57386),
            .in2(N__25759),
            .in3(N__56642),
            .lcout(n22207),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_2__bdd_4_lut_19428_LC_9_14_3.C_ON=1'b0;
    defparam comm_cmd_2__bdd_4_lut_19428_LC_9_14_3.SEQ_MODE=4'b0000;
    defparam comm_cmd_2__bdd_4_lut_19428_LC_9_14_3.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_cmd_2__bdd_4_lut_19428_LC_9_14_3 (
            .in0(N__56374),
            .in1(N__47752),
            .in2(N__28999),
            .in3(N__56336),
            .lcout(),
            .ltout(n22027_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22027_bdd_4_lut_LC_9_14_4.C_ON=1'b0;
    defparam n22027_bdd_4_lut_LC_9_14_4.SEQ_MODE=4'b0000;
    defparam n22027_bdd_4_lut_LC_9_14_4.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22027_bdd_4_lut_LC_9_14_4 (
            .in0(N__56337),
            .in1(N__25729),
            .in2(N__25723),
            .in3(N__25645),
            .lcout(n22030),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22207_bdd_4_lut_LC_9_14_5.C_ON=1'b0;
    defparam n22207_bdd_4_lut_LC_9_14_5.SEQ_MODE=4'b0000;
    defparam n22207_bdd_4_lut_LC_9_14_5.LUT_INIT=16'b1111101001000100;
    LogicCell40 n22207_bdd_4_lut_LC_9_14_5 (
            .in0(N__57387),
            .in1(N__25710),
            .in2(N__25675),
            .in3(N__25651),
            .lcout(n20801),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.bit_cnt_i3_LC_9_15_0 .C_ON=1'b0;
    defparam \SIG_DDS.bit_cnt_i3_LC_9_15_0 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.bit_cnt_i3_LC_9_15_0 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \SIG_DDS.bit_cnt_i3_LC_9_15_0  (
            .in0(N__43687),
            .in1(N__25912),
            .in2(N__25939),
            .in3(N__25786),
            .lcout(\SIG_DDS.bit_cnt_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55164),
            .ce(N__55672),
            .sr(N__43711));
    defparam \SIG_DDS.bit_cnt_i1_LC_9_15_1 .C_ON=1'b0;
    defparam \SIG_DDS.bit_cnt_i1_LC_9_15_1 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.bit_cnt_i1_LC_9_15_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \SIG_DDS.bit_cnt_i1_LC_9_15_1  (
            .in0(_gnd_net_),
            .in1(N__25930),
            .in2(_gnd_net_),
            .in3(N__43685),
            .lcout(\SIG_DDS.bit_cnt_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55164),
            .ce(N__55672),
            .sr(N__43711));
    defparam i18250_3_lut_LC_9_15_3.C_ON=1'b0;
    defparam i18250_3_lut_LC_9_15_3.SEQ_MODE=4'b0000;
    defparam i18250_3_lut_LC_9_15_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 i18250_3_lut_LC_9_15_3 (
            .in0(N__25968),
            .in1(N__31945),
            .in2(_gnd_net_),
            .in3(N__57391),
            .lcout(n20845),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.bit_cnt_i2_LC_9_15_4 .C_ON=1'b0;
    defparam \SIG_DDS.bit_cnt_i2_LC_9_15_4 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.bit_cnt_i2_LC_9_15_4 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \SIG_DDS.bit_cnt_i2_LC_9_15_4  (
            .in0(N__43686),
            .in1(_gnd_net_),
            .in2(N__25938),
            .in3(N__25911),
            .lcout(\SIG_DDS.bit_cnt_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55164),
            .ce(N__55672),
            .sr(N__43711));
    defparam mux_129_Mux_3_i16_3_lut_LC_9_15_6.C_ON=1'b0;
    defparam mux_129_Mux_3_i16_3_lut_LC_9_15_6.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_3_i16_3_lut_LC_9_15_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_129_Mux_3_i16_3_lut_LC_9_15_6 (
            .in0(N__56694),
            .in1(N__31827),
            .in2(_gnd_net_),
            .in3(N__36713),
            .lcout(n16_adj_1500),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_3_i19_3_lut_LC_9_15_7.C_ON=1'b0;
    defparam mux_129_Mux_3_i19_3_lut_LC_9_15_7.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_3_i19_3_lut_LC_9_15_7.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_129_Mux_3_i19_3_lut_LC_9_15_7 (
            .in0(N__26698),
            .in1(N__25889),
            .in2(_gnd_net_),
            .in3(N__56693),
            .lcout(n19_adj_1501),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i15_LC_9_16_0 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i15_LC_9_16_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i15_LC_9_16_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i15_LC_9_16_0  (
            .in0(N__48969),
            .in1(N__50801),
            .in2(N__25872),
            .in3(N__31979),
            .lcout(buf_adcdata_iac_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55179),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_4_lut_adj_261_LC_9_16_1.C_ON=1'b0;
    defparam i3_4_lut_adj_261_LC_9_16_1.SEQ_MODE=4'b0000;
    defparam i3_4_lut_adj_261_LC_9_16_1.LUT_INIT=16'b0000000000000010;
    LogicCell40 i3_4_lut_adj_261_LC_9_16_1 (
            .in0(N__54719),
            .in1(N__39187),
            .in2(N__25840),
            .in3(N__53536),
            .lcout(n10503),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22117_bdd_4_lut_LC_9_16_2.C_ON=1'b0;
    defparam n22117_bdd_4_lut_LC_9_16_2.SEQ_MODE=4'b0000;
    defparam n22117_bdd_4_lut_LC_9_16_2.LUT_INIT=16'b1100110011100010;
    LogicCell40 n22117_bdd_4_lut_LC_9_16_2 (
            .in0(N__28237),
            .in1(N__25831),
            .in2(N__25819),
            .in3(N__47824),
            .lcout(n22120),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.i18704_2_lut_LC_9_16_4 .C_ON=1'b0;
    defparam \SIG_DDS.i18704_2_lut_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \SIG_DDS.i18704_2_lut_LC_9_16_4 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \SIG_DDS.i18704_2_lut_LC_9_16_4  (
            .in0(N__25785),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55887),
            .lcout(\SIG_DDS.n21292 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i5_LC_9_16_5.C_ON=1'b0;
    defparam buf_device_acadc_i5_LC_9_16_5.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i5_LC_9_16_5.LUT_INIT=16'b1011101110001000;
    LogicCell40 buf_device_acadc_i5_LC_9_16_5 (
            .in0(N__42144),
            .in1(N__39236),
            .in2(_gnd_net_),
            .in3(N__26096),
            .lcout(VAC_OSR0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55179),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19467_LC_9_16_6.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19467_LC_9_16_6.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19467_LC_9_16_6.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_0__bdd_4_lut_19467_LC_9_16_6 (
            .in0(N__28085),
            .in1(N__57370),
            .in2(N__26070),
            .in3(N__56686),
            .lcout(n22075),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i17_LC_9_17_0 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i17_LC_9_17_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i17_LC_9_17_0 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \ADC_IAC.ADC_DATA_i17_LC_9_17_0  (
            .in0(N__26027),
            .in1(N__27777),
            .in2(N__50937),
            .in3(N__48960),
            .lcout(buf_adcdata_iac_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55194),
            .ce(),
            .sr(_gnd_net_));
    defparam trig_dds0_304_LC_9_17_1.C_ON=1'b0;
    defparam trig_dds0_304_LC_9_17_1.SEQ_MODE=4'b1000;
    defparam trig_dds0_304_LC_9_17_1.LUT_INIT=16'b0111010000110000;
    LogicCell40 trig_dds0_304_LC_9_17_1 (
            .in0(N__52111),
            .in1(N__26047),
            .in2(N__53005),
            .in3(N__54720),
            .lcout(trig_dds0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55194),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19556_LC_9_17_2.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19556_LC_9_17_2.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19556_LC_9_17_2.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_0__bdd_4_lut_19556_LC_9_17_2 (
            .in0(N__28050),
            .in1(N__57389),
            .in2(N__26031),
            .in3(N__56802),
            .lcout(),
            .ltout(n22201_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22201_bdd_4_lut_LC_9_17_3.C_ON=1'b0;
    defparam n22201_bdd_4_lut_LC_9_17_3.SEQ_MODE=4'b0000;
    defparam n22201_bdd_4_lut_LC_9_17_3.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22201_bdd_4_lut_LC_9_17_3 (
            .in0(N__57390),
            .in1(N__32336),
            .in2(N__26011),
            .in3(N__27571),
            .lcout(n20805),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_start_329_LC_9_17_5.C_ON=1'b0;
    defparam eis_start_329_LC_9_17_5.SEQ_MODE=4'b1000;
    defparam eis_start_329_LC_9_17_5.LUT_INIT=16'b1011101110001000;
    LogicCell40 eis_start_329_LC_9_17_5 (
            .in0(N__43474),
            .in1(N__29879),
            .in2(_gnd_net_),
            .in3(N__30442),
            .lcout(eis_start),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55194),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i16_LC_9_17_7 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i16_LC_9_17_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i16_LC_9_17_7 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_IAC.ADC_DATA_i16_LC_9_17_7  (
            .in0(N__48959),
            .in1(N__50884),
            .in2(N__27993),
            .in3(N__25992),
            .lcout(buf_adcdata_iac_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55194),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i25_LC_9_18_0 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i25_LC_9_18_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i25_LC_9_18_0 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i25_LC_9_18_0  (
            .in0(N__27773),
            .in1(N__50951),
            .in2(N__25993),
            .in3(N__50453),
            .lcout(cmd_rdadctmp_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55208),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19447_LC_9_18_2.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19447_LC_9_18_2.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19447_LC_9_18_2.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_0__bdd_4_lut_19447_LC_9_18_2 (
            .in0(N__26207),
            .in1(N__57484),
            .in2(N__26262),
            .in3(N__56801),
            .lcout(n22045),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i23_LC_9_18_3 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i23_LC_9_18_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i23_LC_9_18_3 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i23_LC_9_18_3  (
            .in0(N__50949),
            .in1(N__48911),
            .in2(N__26293),
            .in3(N__26258),
            .lcout(buf_adcdata_iac_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55208),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_rst_I_0_1_lut_LC_9_18_4.C_ON=1'b0;
    defparam acadc_rst_I_0_1_lut_LC_9_18_4.SEQ_MODE=4'b0000;
    defparam acadc_rst_I_0_1_lut_LC_9_18_4.LUT_INIT=16'b0101010101010101;
    LogicCell40 acadc_rst_I_0_1_lut_LC_9_18_4 (
            .in0(N__32101),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(AC_ADC_SYNC),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i8_LC_9_18_5.C_ON=1'b0;
    defparam buf_device_acadc_i8_LC_9_18_5.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i8_LC_9_18_5.LUT_INIT=16'b1011101110001000;
    LogicCell40 buf_device_acadc_i8_LC_9_18_5 (
            .in0(N__45765),
            .in1(N__39237),
            .in2(_gnd_net_),
            .in3(N__26208),
            .lcout(VAC_FLT1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55208),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i18_LC_9_18_6 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i18_LC_9_18_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i18_LC_9_18_6 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i18_LC_9_18_6  (
            .in0(N__48910),
            .in1(N__50950),
            .in2(N__27756),
            .in3(N__27800),
            .lcout(buf_adcdata_iac_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55208),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.SCLK_35_LC_9_19_7 .C_ON=1'b0;
    defparam \ADC_IAC.SCLK_35_LC_9_19_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.SCLK_35_LC_9_19_7 .LUT_INIT=16'b1101000011100100;
    LogicCell40 \ADC_IAC.SCLK_35_LC_9_19_7  (
            .in0(N__50723),
            .in1(N__30021),
            .in2(N__26184),
            .in3(N__29950),
            .lcout(IAC_SCLK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55220),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i11_3_lut_LC_10_3_0 .C_ON=1'b0;
    defparam \ADC_VDC.i11_3_lut_LC_10_3_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i11_3_lut_LC_10_3_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \ADC_VDC.i11_3_lut_LC_10_3_0  (
            .in0(N__27013),
            .in1(N__28276),
            .in2(_gnd_net_),
            .in3(N__27022),
            .lcout(\ADC_VDC.n18394 ),
            .ltout(\ADC_VDC.n18394_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i15984_3_lut_LC_10_3_1 .C_ON=1'b0;
    defparam \ADC_VDC.i15984_3_lut_LC_10_3_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i15984_3_lut_LC_10_3_1 .LUT_INIT=16'b0011001111111100;
    LogicCell40 \ADC_VDC.i15984_3_lut_LC_10_3_1  (
            .in0(_gnd_net_),
            .in1(N__34773),
            .in2(N__26167),
            .in3(N__34114),
            .lcout(\ADC_VDC.n18397 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam EIS_SYNCCLK_I_0_1_lut_LC_10_3_6.C_ON=1'b0;
    defparam EIS_SYNCCLK_I_0_1_lut_LC_10_3_6.SEQ_MODE=4'b0000;
    defparam EIS_SYNCCLK_I_0_1_lut_LC_10_3_6.LUT_INIT=16'b0000000011111111;
    LogicCell40 EIS_SYNCCLK_I_0_1_lut_LC_10_3_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26164),
            .lcout(IAC_CLK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i37_4_lut_LC_10_4_0 .C_ON=1'b0;
    defparam \ADC_VDC.i37_4_lut_LC_10_4_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i37_4_lut_LC_10_4_0 .LUT_INIT=16'b1110011001000110;
    LogicCell40 \ADC_VDC.i37_4_lut_LC_10_4_0  (
            .in0(N__34770),
            .in1(N__34876),
            .in2(N__34148),
            .in3(N__30679),
            .lcout(),
            .ltout(\ADC_VDC.n31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_4_lut_adj_36_LC_10_4_1 .C_ON=1'b0;
    defparam \ADC_VDC.i1_4_lut_adj_36_LC_10_4_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_4_lut_adj_36_LC_10_4_1 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \ADC_VDC.i1_4_lut_adj_36_LC_10_4_1  (
            .in0(N__28285),
            .in1(N__34589),
            .in2(N__26335),
            .in3(N__34299),
            .lcout(\ADC_VDC.n20514 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.adc_state_1__bdd_4_lut_4_lut_LC_10_4_2 .C_ON=1'b0;
    defparam \ADC_VDC.adc_state_1__bdd_4_lut_4_lut_LC_10_4_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.adc_state_1__bdd_4_lut_4_lut_LC_10_4_2 .LUT_INIT=16'b0010110001101100;
    LogicCell40 \ADC_VDC.adc_state_1__bdd_4_lut_4_lut_LC_10_4_2  (
            .in0(N__34771),
            .in1(N__34120),
            .in2(N__34630),
            .in3(N__26307),
            .lcout(),
            .ltout(\ADC_VDC.n21925_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.n21925_bdd_4_lut_4_lut_LC_10_4_3 .C_ON=1'b0;
    defparam \ADC_VDC.n21925_bdd_4_lut_4_lut_LC_10_4_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.n21925_bdd_4_lut_4_lut_LC_10_4_3 .LUT_INIT=16'b1010010011110100;
    LogicCell40 \ADC_VDC.n21925_bdd_4_lut_4_lut_LC_10_4_3  (
            .in0(N__34593),
            .in1(N__30649),
            .in2(N__26332),
            .in3(N__34772),
            .lcout(),
            .ltout(\ADC_VDC.n21928_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.adc_state_i1_LC_10_4_4 .C_ON=1'b0;
    defparam \ADC_VDC.adc_state_i1_LC_10_4_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.adc_state_i1_LC_10_4_4 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \ADC_VDC.adc_state_i1_LC_10_4_4  (
            .in0(N__26329),
            .in1(N__34594),
            .in2(N__26323),
            .in3(N__34355),
            .lcout(\ADC_VDC.adc_state_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32846),
            .ce(N__26320),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_2_lut_3_lut_LC_10_4_5 .C_ON=1'b0;
    defparam \ADC_VDC.i1_2_lut_3_lut_LC_10_4_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_2_lut_3_lut_LC_10_4_5 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \ADC_VDC.i1_2_lut_3_lut_LC_10_4_5  (
            .in0(N__32515),
            .in1(N__32551),
            .in2(_gnd_net_),
            .in3(N__30667),
            .lcout(),
            .ltout(\ADC_VDC.n6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i4_4_lut_LC_10_4_6 .C_ON=1'b0;
    defparam \ADC_VDC.i4_4_lut_LC_10_4_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i4_4_lut_LC_10_4_6 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \ADC_VDC.i4_4_lut_LC_10_4_6  (
            .in0(N__32470),
            .in1(N__32641),
            .in2(N__26311),
            .in3(N__32599),
            .lcout(\ADC_VDC.n10519 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i3_LC_10_5_0 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i3_LC_10_5_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i3_LC_10_5_0 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i3_LC_10_5_0  (
            .in0(N__34259),
            .in1(N__26798),
            .in2(N__26389),
            .in3(N__26586),
            .lcout(cmd_rdadctmp_3_adj_1469),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32880),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_3_lut_4_lut_adj_40_LC_10_5_1 .C_ON=1'b0;
    defparam \ADC_VDC.i1_3_lut_4_lut_adj_40_LC_10_5_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_3_lut_4_lut_adj_40_LC_10_5_1 .LUT_INIT=16'b1101110000000000;
    LogicCell40 \ADC_VDC.i1_3_lut_4_lut_adj_40_LC_10_5_1  (
            .in0(N__34096),
            .in1(N__34257),
            .in2(N__34751),
            .in3(N__34503),
            .lcout(n12853),
            .ltout(n12853_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i1_LC_10_5_2 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i1_LC_10_5_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i1_LC_10_5_2 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i1_LC_10_5_2  (
            .in0(N__34258),
            .in1(N__26610),
            .in2(N__26296),
            .in3(N__26408),
            .lcout(cmd_rdadctmp_1_adj_1471),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32880),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i0_LC_10_5_3 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i0_LC_10_5_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i0_LC_10_5_3 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i0_LC_10_5_3  (
            .in0(N__26797),
            .in1(N__26609),
            .in2(N__34879),
            .in3(N__34260),
            .lcout(cmd_rdadctmp_0_adj_1472),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32880),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_4_lut_4_lut_4_lut_LC_10_5_4 .C_ON=1'b0;
    defparam \ADC_VDC.i1_4_lut_4_lut_4_lut_LC_10_5_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_4_lut_4_lut_4_lut_LC_10_5_4 .LUT_INIT=16'b1110001010100000;
    LogicCell40 \ADC_VDC.i1_4_lut_4_lut_4_lut_LC_10_5_4  (
            .in0(N__34255),
            .in1(N__34723),
            .in2(N__34564),
            .in3(N__34094),
            .lcout(\ADC_VDC.n13060 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i4_LC_10_5_5 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i4_LC_10_5_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i4_LC_10_5_5 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i4_LC_10_5_5  (
            .in0(N__26585),
            .in1(N__26564),
            .in2(N__26836),
            .in3(N__34261),
            .lcout(cmd_rdadctmp_4_adj_1468),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32880),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_4_lut_adj_43_LC_10_5_6 .C_ON=1'b0;
    defparam \ADC_VDC.i1_4_lut_adj_43_LC_10_5_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_4_lut_adj_43_LC_10_5_6 .LUT_INIT=16'b1011000011100000;
    LogicCell40 \ADC_VDC.i1_4_lut_adj_43_LC_10_5_6  (
            .in0(N__34256),
            .in1(N__34724),
            .in2(N__34565),
            .in3(N__34095),
            .lcout(\ADC_VDC.n12885 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i8_LC_10_5_7 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i8_LC_10_5_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i8_LC_10_5_7 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i8_LC_10_5_7  (
            .in0(N__26504),
            .in1(N__26532),
            .in2(N__26837),
            .in3(N__34262),
            .lcout(cmd_rdadctmp_8_adj_1464),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32880),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i17_LC_10_6_0 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i17_LC_10_6_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i17_LC_10_6_0 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i17_LC_10_6_0  (
            .in0(N__34303),
            .in1(N__26427),
            .in2(N__26879),
            .in3(N__26480),
            .lcout(cmd_rdadctmp_17_adj_1455),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32912),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i16_LC_10_6_1 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i16_LC_10_6_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i16_LC_10_6_1 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i16_LC_10_6_1  (
            .in0(N__26426),
            .in1(N__34306),
            .in2(N__26458),
            .in3(N__26842),
            .lcout(cmd_rdadctmp_16_adj_1456),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32912),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i2_LC_10_6_2 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i2_LC_10_6_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i2_LC_10_6_2 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i2_LC_10_6_2  (
            .in0(N__34304),
            .in1(N__26387),
            .in2(N__26880),
            .in3(N__26409),
            .lcout(cmd_rdadctmp_2_adj_1470),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32912),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i12_LC_10_6_3 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i12_LC_10_6_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i12_LC_10_6_3 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i12_LC_10_6_3  (
            .in0(N__26958),
            .in1(N__34305),
            .in2(N__26364),
            .in3(N__26841),
            .lcout(cmd_rdadctmp_12_adj_1460),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32912),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i11_LC_10_6_4 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i11_LC_10_6_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i11_LC_10_6_4 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i11_LC_10_6_4  (
            .in0(N__34302),
            .in1(N__26957),
            .in2(N__26878),
            .in3(N__26989),
            .lcout(cmd_rdadctmp_11_adj_1461),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32912),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i19078_2_lut_LC_10_6_5 .C_ON=1'b0;
    defparam \ADC_VDC.i19078_2_lut_LC_10_6_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i19078_2_lut_LC_10_6_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ADC_VDC.i19078_2_lut_LC_10_6_5  (
            .in0(_gnd_net_),
            .in1(N__34584),
            .in2(_gnd_net_),
            .in3(N__34301),
            .lcout(),
            .ltout(\ADC_VDC.n21673_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.SCLK_46_LC_10_6_6 .C_ON=1'b0;
    defparam \ADC_VDC.SCLK_46_LC_10_6_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.SCLK_46_LC_10_6_6 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \ADC_VDC.SCLK_46_LC_10_6_6  (
            .in0(N__26931),
            .in1(N__30613),
            .in2(N__26941),
            .in3(N__34141),
            .lcout(VDC_SCLK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32912),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i20_LC_10_6_7 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i20_LC_10_6_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i20_LC_10_6_7 .LUT_INIT=16'b0000110010101010;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i20_LC_10_6_7  (
            .in0(N__26768),
            .in1(N__26920),
            .in2(N__34393),
            .in3(N__26846),
            .lcout(cmd_rdadctmp_20_adj_1452),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32912),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i12_LC_10_7_0 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i12_LC_10_7_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i12_LC_10_7_0 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \ADC_VDC.ADC_DATA_i12_LC_10_7_0  (
            .in0(N__34567),
            .in1(N__28369),
            .in2(N__26727),
            .in3(N__26746),
            .lcout(buf_adcdata_vdc_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32871),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i11_LC_10_7_1 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i11_LC_10_7_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i11_LC_10_7_1 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i11_LC_10_7_1  (
            .in0(N__28365),
            .in1(N__34571),
            .in2(N__26691),
            .in3(N__26710),
            .lcout(buf_adcdata_vdc_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32871),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i4_LC_10_7_2 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i4_LC_10_7_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i4_LC_10_7_2 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \ADC_VDC.ADC_DATA_i4_LC_10_7_2  (
            .in0(N__34568),
            .in1(N__28370),
            .in2(N__26674),
            .in3(N__51342),
            .lcout(buf_adcdata_vdc_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32871),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i9_LC_10_7_3 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i9_LC_10_7_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i9_LC_10_7_3 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i9_LC_10_7_3  (
            .in0(N__28368),
            .in1(N__34573),
            .in2(N__35301),
            .in3(N__26659),
            .lcout(buf_adcdata_vdc_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32871),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i8_LC_10_7_4 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i8_LC_10_7_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i8_LC_10_7_4 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \ADC_VDC.ADC_DATA_i8_LC_10_7_4  (
            .in0(N__34570),
            .in1(N__28371),
            .in2(N__26628),
            .in3(N__26647),
            .lcout(buf_adcdata_vdc_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32871),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i7_LC_10_7_5 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i7_LC_10_7_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i7_LC_10_7_5 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i7_LC_10_7_5  (
            .in0(N__28367),
            .in1(N__34572),
            .in2(N__47898),
            .in3(N__27115),
            .lcout(buf_adcdata_vdc_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32871),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i6_LC_10_7_6 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i6_LC_10_7_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i6_LC_10_7_6 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \ADC_VDC.ADC_DATA_i6_LC_10_7_6  (
            .in0(N__34569),
            .in1(N__27103),
            .in2(N__40881),
            .in3(N__28372),
            .lcout(buf_adcdata_vdc_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32871),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i5_LC_10_7_7 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i5_LC_10_7_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i5_LC_10_7_7 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \ADC_VDC.ADC_DATA_i5_LC_10_7_7  (
            .in0(N__28366),
            .in1(N__34574),
            .in2(N__27091),
            .in3(N__38319),
            .lcout(buf_adcdata_vdc_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32871),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_3_lut_4_lut_4_lut_LC_10_8_1 .C_ON=1'b0;
    defparam \ADC_VDC.i1_3_lut_4_lut_4_lut_LC_10_8_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_3_lut_4_lut_4_lut_LC_10_8_1 .LUT_INIT=16'b1110001010100010;
    LogicCell40 \ADC_VDC.i1_3_lut_4_lut_4_lut_LC_10_8_1  (
            .in0(N__34385),
            .in1(N__34774),
            .in2(N__34642),
            .in3(N__34149),
            .lcout(\ADC_VDC.n13020 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i18765_3_lut_LC_10_8_2 .C_ON=1'b0;
    defparam \ADC_VDC.i18765_3_lut_LC_10_8_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i18765_3_lut_LC_10_8_2 .LUT_INIT=16'b0010001000010001;
    LogicCell40 \ADC_VDC.i18765_3_lut_LC_10_8_2  (
            .in0(N__27048),
            .in1(N__34624),
            .in2(_gnd_net_),
            .in3(N__27076),
            .lcout(),
            .ltout(\ADC_VDC.n21106_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadcbuf_i34_LC_10_8_3 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadcbuf_i34_LC_10_8_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i34_LC_10_8_3 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i34_LC_10_8_3  (
            .in0(N__34386),
            .in1(N__27067),
            .in2(N__27058),
            .in3(N__34150),
            .lcout(cmd_rdadcbuf_34),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32913),
            .ce(N__27031),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i9_4_lut_LC_10_8_5 .C_ON=1'b0;
    defparam \ADC_VDC.i9_4_lut_LC_10_8_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i9_4_lut_LC_10_8_5 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \ADC_VDC.i9_4_lut_LC_10_8_5  (
            .in0(N__29202),
            .in1(N__28497),
            .in2(N__28516),
            .in3(N__28434),
            .lcout(\ADC_VDC.n21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i7_4_lut_LC_10_8_6 .C_ON=1'b0;
    defparam \ADC_VDC.i7_4_lut_LC_10_8_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i7_4_lut_LC_10_8_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.i7_4_lut_LC_10_8_6  (
            .in0(N__29235),
            .in1(N__28530),
            .in2(N__29257),
            .in3(N__29220),
            .lcout(\ADC_VDC.n19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_3__i0_LC_10_9_0.C_ON=1'b0;
    defparam comm_buf_3__i0_LC_10_9_0.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i0_LC_10_9_0.LUT_INIT=16'b1110111000100010;
    LogicCell40 comm_buf_3__i0_LC_10_9_0 (
            .in0(N__27004),
            .in1(N__54086),
            .in2(_gnd_net_),
            .in3(N__36242),
            .lcout(comm_buf_3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55088),
            .ce(N__27259),
            .sr(N__27250));
    defparam comm_buf_3__i7_LC_10_9_1.C_ON=1'b0;
    defparam comm_buf_3__i7_LC_10_9_1.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i7_LC_10_9_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_3__i7_LC_10_9_1 (
            .in0(N__54085),
            .in1(N__36898),
            .in2(_gnd_net_),
            .in3(N__27226),
            .lcout(comm_buf_3_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55088),
            .ce(N__27259),
            .sr(N__27250));
    defparam comm_buf_3__i6_LC_10_9_2.C_ON=1'b0;
    defparam comm_buf_3__i6_LC_10_9_2.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i6_LC_10_9_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 comm_buf_3__i6_LC_10_9_2 (
            .in0(N__35798),
            .in1(N__54089),
            .in2(_gnd_net_),
            .in3(N__27208),
            .lcout(comm_buf_3_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55088),
            .ce(N__27259),
            .sr(N__27250));
    defparam comm_buf_3__i5_LC_10_9_3.C_ON=1'b0;
    defparam comm_buf_3__i5_LC_10_9_3.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i5_LC_10_9_3.LUT_INIT=16'b1111101001010000;
    LogicCell40 comm_buf_3__i5_LC_10_9_3 (
            .in0(N__54084),
            .in1(_gnd_net_),
            .in2(N__27190),
            .in3(N__37995),
            .lcout(comm_buf_3_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55088),
            .ce(N__27259),
            .sr(N__27250));
    defparam comm_buf_3__i4_LC_10_9_4.C_ON=1'b0;
    defparam comm_buf_3__i4_LC_10_9_4.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i4_LC_10_9_4.LUT_INIT=16'b1011101110001000;
    LogicCell40 comm_buf_3__i4_LC_10_9_4 (
            .in0(N__35640),
            .in1(N__54088),
            .in2(_gnd_net_),
            .in3(N__27175),
            .lcout(comm_buf_3_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55088),
            .ce(N__27259),
            .sr(N__27250));
    defparam comm_buf_3__i3_LC_10_9_5.C_ON=1'b0;
    defparam comm_buf_3__i3_LC_10_9_5.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i3_LC_10_9_5.LUT_INIT=16'b1110111001000100;
    LogicCell40 comm_buf_3__i3_LC_10_9_5 (
            .in0(N__54083),
            .in1(N__27157),
            .in2(_gnd_net_),
            .in3(N__35558),
            .lcout(comm_buf_3_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55088),
            .ce(N__27259),
            .sr(N__27250));
    defparam comm_buf_3__i2_LC_10_9_6.C_ON=1'b0;
    defparam comm_buf_3__i2_LC_10_9_6.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i2_LC_10_9_6.LUT_INIT=16'b1011101110001000;
    LogicCell40 comm_buf_3__i2_LC_10_9_6 (
            .in0(N__35441),
            .in1(N__54087),
            .in2(_gnd_net_),
            .in3(N__27148),
            .lcout(comm_buf_3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55088),
            .ce(N__27259),
            .sr(N__27250));
    defparam comm_buf_3__i1_LC_10_9_7.C_ON=1'b0;
    defparam comm_buf_3__i1_LC_10_9_7.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i1_LC_10_9_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_3__i1_LC_10_9_7 (
            .in0(N__54082),
            .in1(N__35977),
            .in2(_gnd_net_),
            .in3(N__27133),
            .lcout(comm_buf_3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55088),
            .ce(N__27259),
            .sr(N__27250));
    defparam i18988_2_lut_4_lut_LC_10_10_0.C_ON=1'b0;
    defparam i18988_2_lut_4_lut_LC_10_10_0.SEQ_MODE=4'b0000;
    defparam i18988_2_lut_4_lut_LC_10_10_0.LUT_INIT=16'b0000000001000000;
    LogicCell40 i18988_2_lut_4_lut_LC_10_10_0 (
            .in0(N__50096),
            .in1(N__49539),
            .in2(N__49957),
            .in3(N__53530),
            .lcout(),
            .ltout(n21143_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19_4_lut_adj_293_LC_10_10_1.C_ON=1'b0;
    defparam i19_4_lut_adj_293_LC_10_10_1.SEQ_MODE=4'b0000;
    defparam i19_4_lut_adj_293_LC_10_10_1.LUT_INIT=16'b1000000011010101;
    LogicCell40 i19_4_lut_adj_293_LC_10_10_1 (
            .in0(N__54079),
            .in1(N__51643),
            .in2(N__27118),
            .in3(N__51685),
            .lcout(),
            .ltout(n12_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_294_LC_10_10_2.C_ON=1'b0;
    defparam i1_3_lut_adj_294_LC_10_10_2.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_294_LC_10_10_2.LUT_INIT=16'b1111110000000000;
    LogicCell40 i1_3_lut_adj_294_LC_10_10_2 (
            .in0(_gnd_net_),
            .in1(N__49914),
            .in2(N__27262),
            .in3(N__49869),
            .lcout(n12116),
            .ltout(n12116_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12359_2_lut_LC_10_10_3.C_ON=1'b0;
    defparam i12359_2_lut_LC_10_10_3.SEQ_MODE=4'b0000;
    defparam i12359_2_lut_LC_10_10_3.LUT_INIT=16'b1111000000000000;
    LogicCell40 i12359_2_lut_LC_10_10_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27253),
            .in3(N__54701),
            .lcout(n14756),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_279_LC_10_10_4.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_279_LC_10_10_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_279_LC_10_10_4.LUT_INIT=16'b0001000100000000;
    LogicCell40 i1_2_lut_3_lut_adj_279_LC_10_10_4 (
            .in0(N__50095),
            .in1(N__53529),
            .in2(_gnd_net_),
            .in3(N__49947),
            .lcout(),
            .ltout(n25_adj_1592_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_288_LC_10_10_5.C_ON=1'b0;
    defparam i1_4_lut_adj_288_LC_10_10_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_288_LC_10_10_5.LUT_INIT=16'b1100110011011100;
    LogicCell40 i1_4_lut_adj_288_LC_10_10_5 (
            .in0(N__49538),
            .in1(N__46077),
            .in2(N__27238),
            .in3(N__51642),
            .lcout(),
            .ltout(n11944_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_289_LC_10_10_6.C_ON=1'b0;
    defparam i1_4_lut_adj_289_LC_10_10_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_289_LC_10_10_6.LUT_INIT=16'b1100000010000000;
    LogicCell40 i1_4_lut_adj_289_LC_10_10_6 (
            .in0(N__46429),
            .in1(N__49870),
            .in2(N__27235),
            .in3(N__37515),
            .lcout(n11941),
            .ltout(n11941_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12338_2_lut_LC_10_10_7.C_ON=1'b0;
    defparam i12338_2_lut_LC_10_10_7.SEQ_MODE=4'b0000;
    defparam i12338_2_lut_LC_10_10_7.LUT_INIT=16'b1111000000000000;
    LogicCell40 i12338_2_lut_LC_10_10_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27232),
            .in3(N__54700),
            .lcout(n14735),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19331_LC_10_11_0.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19331_LC_10_11_0.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19331_LC_10_11_0.LUT_INIT=16'b1110110001100100;
    LogicCell40 comm_cmd_0__bdd_4_lut_19331_LC_10_11_0 (
            .in0(N__57408),
            .in1(N__56797),
            .in2(N__41926),
            .in3(N__32100),
            .lcout(),
            .ltout(n21919_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n21919_bdd_4_lut_LC_10_11_1.C_ON=1'b0;
    defparam n21919_bdd_4_lut_LC_10_11_1.SEQ_MODE=4'b0000;
    defparam n21919_bdd_4_lut_LC_10_11_1.LUT_INIT=16'b1111001011000010;
    LogicCell40 n21919_bdd_4_lut_LC_10_11_1 (
            .in0(N__38175),
            .in1(N__57409),
            .in2(N__27229),
            .in3(N__38623),
            .lcout(n21922),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18199_3_lut_LC_10_11_2.C_ON=1'b0;
    defparam i18199_3_lut_LC_10_11_2.SEQ_MODE=4'b0000;
    defparam i18199_3_lut_LC_10_11_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 i18199_3_lut_LC_10_11_2 (
            .in0(N__31176),
            .in1(N__56798),
            .in2(_gnd_net_),
            .in3(N__47274),
            .lcout(),
            .ltout(n20794_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18201_4_lut_LC_10_11_3.C_ON=1'b0;
    defparam i18201_4_lut_LC_10_11_3.SEQ_MODE=4'b0000;
    defparam i18201_4_lut_LC_10_11_3.LUT_INIT=16'b1110111011110000;
    LogicCell40 i18201_4_lut_LC_10_11_3 (
            .in0(N__56800),
            .in1(N__27373),
            .in2(N__27358),
            .in3(N__57410),
            .lcout(),
            .ltout(n20796_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_2__bdd_4_lut_LC_10_11_4.C_ON=1'b0;
    defparam comm_cmd_2__bdd_4_lut_LC_10_11_4.SEQ_MODE=4'b0000;
    defparam comm_cmd_2__bdd_4_lut_LC_10_11_4.LUT_INIT=16'b1111010110001000;
    LogicCell40 comm_cmd_2__bdd_4_lut_LC_10_11_4 (
            .in0(N__56308),
            .in1(N__27355),
            .in2(N__27349),
            .in3(N__47694),
            .lcout(),
            .ltout(n22213_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22213_bdd_4_lut_LC_10_11_5.C_ON=1'b0;
    defparam n22213_bdd_4_lut_LC_10_11_5.SEQ_MODE=4'b0000;
    defparam n22213_bdd_4_lut_LC_10_11_5.LUT_INIT=16'b1111000010101100;
    LogicCell40 n22213_bdd_4_lut_LC_10_11_5 (
            .in0(N__27346),
            .in1(N__30157),
            .in2(N__27334),
            .in3(N__56309),
            .lcout(),
            .ltout(n22216_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_0__i2_LC_10_11_6.C_ON=1'b0;
    defparam comm_buf_0__i2_LC_10_11_6.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i2_LC_10_11_6.LUT_INIT=16'b1111110000110000;
    LogicCell40 comm_buf_0__i2_LC_10_11_6 (
            .in0(_gnd_net_),
            .in1(N__54101),
            .in2(N__27331),
            .in3(N__35450),
            .lcout(comm_buf_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55105),
            .ce(N__27505),
            .sr(N__27454));
    defparam i19000_4_lut_4_lut_LC_10_11_7.C_ON=1'b0;
    defparam i19000_4_lut_4_lut_LC_10_11_7.SEQ_MODE=4'b0000;
    defparam i19000_4_lut_4_lut_LC_10_11_7.LUT_INIT=16'b1101101011101111;
    LogicCell40 i19000_4_lut_4_lut_LC_10_11_7 (
            .in0(N__56799),
            .in1(N__47508),
            .in2(N__56342),
            .in3(N__57407),
            .lcout(n21071),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19336_LC_10_12_1.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19336_LC_10_12_1.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19336_LC_10_12_1.LUT_INIT=16'b1011101111000000;
    LogicCell40 comm_cmd_1__bdd_4_lut_19336_LC_10_12_1 (
            .in0(N__27328),
            .in1(N__47578),
            .in2(N__27313),
            .in3(N__57462),
            .lcout(),
            .ltout(n21907_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n21907_bdd_4_lut_LC_10_12_2.C_ON=1'b0;
    defparam n21907_bdd_4_lut_LC_10_12_2.SEQ_MODE=4'b0000;
    defparam n21907_bdd_4_lut_LC_10_12_2.LUT_INIT=16'b1111010010100100;
    LogicCell40 n21907_bdd_4_lut_LC_10_12_2 (
            .in0(N__47579),
            .in1(N__28174),
            .in2(N__27304),
            .in3(N__45067),
            .lcout(n21910),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19418_LC_10_12_3.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19418_LC_10_12_3.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19418_LC_10_12_3.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_0__bdd_4_lut_19418_LC_10_12_3 (
            .in0(N__29715),
            .in1(N__57463),
            .in2(N__27300),
            .in3(N__56638),
            .lcout(),
            .ltout(n22033_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22033_bdd_4_lut_LC_10_12_4.C_ON=1'b0;
    defparam n22033_bdd_4_lut_LC_10_12_4.SEQ_MODE=4'b0000;
    defparam n22033_bdd_4_lut_LC_10_12_4.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22033_bdd_4_lut_LC_10_12_4 (
            .in0(N__57464),
            .in1(N__32310),
            .in2(N__27265),
            .in3(N__29393),
            .lcout(),
            .ltout(n22036_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18228_3_lut_LC_10_12_5.C_ON=1'b0;
    defparam i18228_3_lut_LC_10_12_5.SEQ_MODE=4'b0000;
    defparam i18228_3_lut_LC_10_12_5.LUT_INIT=16'b1111110000110000;
    LogicCell40 i18228_3_lut_LC_10_12_5 (
            .in0(_gnd_net_),
            .in1(N__47580),
            .in2(N__27544),
            .in3(N__27541),
            .lcout(),
            .ltout(n20823_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1537450_i1_3_lut_LC_10_12_6.C_ON=1'b0;
    defparam i1537450_i1_3_lut_LC_10_12_6.SEQ_MODE=4'b0000;
    defparam i1537450_i1_3_lut_LC_10_12_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 i1537450_i1_3_lut_LC_10_12_6 (
            .in0(_gnd_net_),
            .in1(N__27529),
            .in2(N__27523),
            .in3(N__56274),
            .lcout(),
            .ltout(n30_adj_1514_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_0__i5_LC_10_12_7.C_ON=1'b0;
    defparam comm_buf_0__i5_LC_10_12_7.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i5_LC_10_12_7.LUT_INIT=16'b1010101011110000;
    LogicCell40 comm_buf_0__i5_LC_10_12_7 (
            .in0(N__38022),
            .in1(_gnd_net_),
            .in2(N__27520),
            .in3(N__54100),
            .lcout(comm_buf_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55116),
            .ce(N__27513),
            .sr(N__27464));
    defparam \CLK_DDS.tmp_buf_i10_LC_10_13_0 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i10_LC_10_13_0 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i10_LC_10_13_0 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \CLK_DDS.tmp_buf_i10_LC_10_13_0  (
            .in0(N__28795),
            .in1(N__28947),
            .in2(N__27628),
            .in3(N__30187),
            .lcout(\CLK_DDS.tmp_buf_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55125),
            .ce(N__28551),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i11_LC_10_13_1 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i11_LC_10_13_1 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i11_LC_10_13_1 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \CLK_DDS.tmp_buf_i11_LC_10_13_1  (
            .in0(N__29556),
            .in1(N__28954),
            .in2(N__27418),
            .in3(N__28799),
            .lcout(\CLK_DDS.tmp_buf_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55125),
            .ce(N__28551),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i12_LC_10_13_2 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i12_LC_10_13_2 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i12_LC_10_13_2 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \CLK_DDS.tmp_buf_i12_LC_10_13_2  (
            .in0(N__28796),
            .in1(N__27588),
            .in2(N__27409),
            .in3(N__28950),
            .lcout(\CLK_DDS.tmp_buf_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55125),
            .ce(N__28551),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i13_LC_10_13_3 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i13_LC_10_13_3 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i13_LC_10_13_3 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLK_DDS.tmp_buf_i13_LC_10_13_3  (
            .in0(N__28951),
            .in1(N__28800),
            .in2(N__27400),
            .in3(N__29401),
            .lcout(\CLK_DDS.tmp_buf_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55125),
            .ce(N__28551),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i14_LC_10_13_4 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i14_LC_10_13_4 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i14_LC_10_13_4 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \CLK_DDS.tmp_buf_i14_LC_10_13_4  (
            .in0(N__28797),
            .in1(N__28948),
            .in2(N__27391),
            .in3(N__27608),
            .lcout(\CLK_DDS.tmp_buf_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55125),
            .ce(N__28551),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i15_LC_10_13_5 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i15_LC_10_13_5 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i15_LC_10_13_5 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLK_DDS.tmp_buf_i15_LC_10_13_5  (
            .in0(N__28952),
            .in1(N__28801),
            .in2(N__27382),
            .in3(N__27920),
            .lcout(tmp_buf_15_adj_1448),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55125),
            .ce(N__28551),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i9_LC_10_13_6 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i9_LC_10_13_6 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i9_LC_10_13_6 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \CLK_DDS.tmp_buf_i9_LC_10_13_6  (
            .in0(N__28798),
            .in1(N__28949),
            .in2(N__27570),
            .in3(N__27619),
            .lcout(\CLK_DDS.tmp_buf_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55125),
            .ce(N__28551),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i8_LC_10_13_7 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i8_LC_10_13_7 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i8_LC_10_13_7 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLK_DDS.tmp_buf_i8_LC_10_13_7  (
            .in0(N__28953),
            .in1(N__28802),
            .in2(N__27640),
            .in3(N__27964),
            .lcout(\CLK_DDS.tmp_buf_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55125),
            .ce(N__28551),
            .sr(_gnd_net_));
    defparam buf_dds1_i14_LC_10_14_0.C_ON=1'b0;
    defparam buf_dds1_i14_LC_10_14_0.SEQ_MODE=4'b1000;
    defparam buf_dds1_i14_LC_10_14_0.LUT_INIT=16'b1000101010000000;
    LogicCell40 buf_dds1_i14_LC_10_14_0 (
            .in0(N__46017),
            .in1(N__40786),
            .in2(N__45914),
            .in3(N__27609),
            .lcout(buf_dds1_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55137),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i12_LC_10_14_1.C_ON=1'b0;
    defparam buf_dds1_i12_LC_10_14_1.SEQ_MODE=4'b1000;
    defparam buf_dds1_i12_LC_10_14_1.LUT_INIT=16'b1110001000000000;
    LogicCell40 buf_dds1_i12_LC_10_14_1 (
            .in0(N__27589),
            .in1(N__45901),
            .in2(N__46708),
            .in3(N__46016),
            .lcout(buf_dds1_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55137),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i15_LC_10_14_2.C_ON=1'b0;
    defparam buf_dds1_i15_LC_10_14_2.SEQ_MODE=4'b1000;
    defparam buf_dds1_i15_LC_10_14_2.LUT_INIT=16'b1000101010000000;
    LogicCell40 buf_dds1_i15_LC_10_14_2 (
            .in0(N__46018),
            .in1(N__30814),
            .in2(N__45915),
            .in3(N__27921),
            .lcout(buf_dds1_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55137),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i11_LC_10_14_3.C_ON=1'b0;
    defparam buf_dds1_i11_LC_10_14_3.SEQ_MODE=4'b1000;
    defparam buf_dds1_i11_LC_10_14_3.LUT_INIT=16'b1110001000000000;
    LogicCell40 buf_dds1_i11_LC_10_14_3 (
            .in0(N__29555),
            .in1(N__45900),
            .in2(N__43806),
            .in3(N__46015),
            .lcout(buf_dds1_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55137),
            .ce(),
            .sr(_gnd_net_));
    defparam trig_dds1_305_LC_10_14_4.C_ON=1'b0;
    defparam trig_dds1_305_LC_10_14_4.SEQ_MODE=4'b1000;
    defparam trig_dds1_305_LC_10_14_4.LUT_INIT=16'b0110000001100100;
    LogicCell40 trig_dds1_305_LC_10_14_4 (
            .in0(N__52169),
            .in1(N__54699),
            .in2(N__28654),
            .in3(N__45937),
            .lcout(trig_dds1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55137),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i9_LC_10_14_6.C_ON=1'b0;
    defparam buf_dds1_i9_LC_10_14_6.SEQ_MODE=4'b1000;
    defparam buf_dds1_i9_LC_10_14_6.LUT_INIT=16'b1000101010000000;
    LogicCell40 buf_dds1_i9_LC_10_14_6 (
            .in0(N__46019),
            .in1(N__44085),
            .in2(N__45916),
            .in3(N__27566),
            .lcout(buf_dds1_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55137),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_stop_328_LC_10_14_7.C_ON=1'b0;
    defparam eis_stop_328_LC_10_14_7.SEQ_MODE=4'b1000;
    defparam eis_stop_328_LC_10_14_7.LUT_INIT=16'b1011101110001000;
    LogicCell40 eis_stop_328_LC_10_14_7 (
            .in0(N__44084),
            .in1(N__29887),
            .in2(_gnd_net_),
            .in3(N__38935),
            .lcout(eis_stop),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55137),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i0_LC_10_15_0 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i0_LC_10_15_0 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i0_LC_10_15_0 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLK_DDS.tmp_buf_i0_LC_10_15_0  (
            .in0(N__28974),
            .in1(N__28804),
            .in2(N__27730),
            .in3(N__27826),
            .lcout(\CLK_DDS.tmp_buf_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55150),
            .ce(N__28555),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i1_LC_10_15_1 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i1_LC_10_15_1 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i1_LC_10_15_1 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \CLK_DDS.tmp_buf_i1_LC_10_15_1  (
            .in0(N__28803),
            .in1(N__28978),
            .in2(N__27706),
            .in3(N__31933),
            .lcout(\CLK_DDS.tmp_buf_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55150),
            .ce(N__28555),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i2_LC_10_15_2 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i2_LC_10_15_2 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i2_LC_10_15_2 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLK_DDS.tmp_buf_i2_LC_10_15_2  (
            .in0(N__28975),
            .in1(N__28805),
            .in2(N__27697),
            .in3(N__32017),
            .lcout(\CLK_DDS.tmp_buf_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55150),
            .ce(N__28555),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i3_LC_10_15_3 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i3_LC_10_15_3 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i3_LC_10_15_3 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \CLK_DDS.tmp_buf_i3_LC_10_15_3  (
            .in0(N__31828),
            .in1(N__28979),
            .in2(N__27688),
            .in3(N__28810),
            .lcout(\CLK_DDS.tmp_buf_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55150),
            .ce(N__28555),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i4_LC_10_15_4 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i4_LC_10_15_4 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i4_LC_10_15_4 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLK_DDS.tmp_buf_i4_LC_10_15_4  (
            .in0(N__28976),
            .in1(N__28806),
            .in2(N__27679),
            .in3(N__36143),
            .lcout(\CLK_DDS.tmp_buf_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55150),
            .ce(N__28555),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i5_LC_10_15_5 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i5_LC_10_15_5 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i5_LC_10_15_5 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLK_DDS.tmp_buf_i5_LC_10_15_5  (
            .in0(N__28980),
            .in1(N__28808),
            .in2(N__27667),
            .in3(N__29508),
            .lcout(\CLK_DDS.tmp_buf_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55150),
            .ce(N__28555),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i6_LC_10_15_6 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i6_LC_10_15_6 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i6_LC_10_15_6 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLK_DDS.tmp_buf_i6_LC_10_15_6  (
            .in0(N__28977),
            .in1(N__28807),
            .in2(N__27658),
            .in3(N__36115),
            .lcout(\CLK_DDS.tmp_buf_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55150),
            .ce(N__28555),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i7_LC_10_15_7 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i7_LC_10_15_7 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i7_LC_10_15_7 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLK_DDS.tmp_buf_i7_LC_10_15_7  (
            .in0(N__28981),
            .in1(N__28809),
            .in2(N__27649),
            .in3(N__42544),
            .lcout(\CLK_DDS.tmp_buf_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55150),
            .ce(N__28555),
            .sr(_gnd_net_));
    defparam buf_dds0_i3_LC_10_16_0.C_ON=1'b0;
    defparam buf_dds0_i3_LC_10_16_0.SEQ_MODE=4'b1000;
    defparam buf_dds0_i3_LC_10_16_0.LUT_INIT=16'b0101110100001000;
    LogicCell40 buf_dds0_i3_LC_10_16_0 (
            .in0(N__45692),
            .in1(N__36397),
            .in2(N__52172),
            .in3(N__36717),
            .lcout(buf_dds0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55165),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i14_LC_10_16_1.C_ON=1'b0;
    defparam buf_dds0_i14_LC_10_16_1.SEQ_MODE=4'b1000;
    defparam buf_dds0_i14_LC_10_16_1.LUT_INIT=16'b1111000010101010;
    LogicCell40 buf_dds0_i14_LC_10_16_1 (
            .in0(N__32258),
            .in1(_gnd_net_),
            .in2(N__41545),
            .in3(N__45691),
            .lcout(buf_dds0_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55165),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i0_LC_10_16_2.C_ON=1'b0;
    defparam acadc_skipCount_i0_LC_10_16_2.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i0_LC_10_16_2.LUT_INIT=16'b0101110100001000;
    LogicCell40 acadc_skipCount_i0_LC_10_16_2 (
            .in0(N__39330),
            .in1(N__41356),
            .in2(N__52171),
            .in3(N__35856),
            .lcout(acadc_skipCount_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55165),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i13_LC_10_16_3.C_ON=1'b0;
    defparam acadc_skipCount_i13_LC_10_16_3.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i13_LC_10_16_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 acadc_skipCount_i13_LC_10_16_3 (
            .in0(N__44846),
            .in1(N__39329),
            .in2(_gnd_net_),
            .in3(N__30205),
            .lcout(acadc_skipCount_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55165),
            .ce(),
            .sr(_gnd_net_));
    defparam n22045_bdd_4_lut_LC_10_16_4.C_ON=1'b0;
    defparam n22045_bdd_4_lut_LC_10_16_4.SEQ_MODE=4'b0000;
    defparam n22045_bdd_4_lut_LC_10_16_4.LUT_INIT=16'b1100110010111000;
    LogicCell40 n22045_bdd_4_lut_LC_10_16_4 (
            .in0(N__27922),
            .in1(N__27901),
            .in2(N__45595),
            .in3(N__57502),
            .lcout(n22048),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i7_LC_10_16_5.C_ON=1'b0;
    defparam buf_device_acadc_i7_LC_10_16_5.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i7_LC_10_16_5.LUT_INIT=16'b1011101110001000;
    LogicCell40 buf_device_acadc_i7_LC_10_16_5 (
            .in0(N__41544),
            .in1(N__39219),
            .in2(_gnd_net_),
            .in3(N__27857),
            .lcout(VAC_FLT0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55165),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_0_i16_3_lut_LC_10_16_6.C_ON=1'b0;
    defparam mux_129_Mux_0_i16_3_lut_LC_10_16_6.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_0_i16_3_lut_LC_10_16_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_129_Mux_0_i16_3_lut_LC_10_16_6 (
            .in0(N__27824),
            .in1(N__40374),
            .in2(_gnd_net_),
            .in3(N__56921),
            .lcout(n16_adj_1480),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i0_LC_10_16_7.C_ON=1'b0;
    defparam buf_dds1_i0_LC_10_16_7.SEQ_MODE=4'b1000;
    defparam buf_dds1_i0_LC_10_16_7.LUT_INIT=16'b1110010000000000;
    LogicCell40 buf_dds1_i0_LC_10_16_7 (
            .in0(N__45840),
            .in1(N__27825),
            .in2(N__41364),
            .in3(N__46020),
            .lcout(buf_dds1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55165),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i8_LC_10_17_1.C_ON=1'b0;
    defparam buf_dds1_i8_LC_10_17_1.SEQ_MODE=4'b1000;
    defparam buf_dds1_i8_LC_10_17_1.LUT_INIT=16'b1110001000000000;
    LogicCell40 buf_dds1_i8_LC_10_17_1 (
            .in0(N__27963),
            .in1(N__45911),
            .in2(N__43533),
            .in3(N__46021),
            .lcout(buf_dds1_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55180),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19511_LC_10_17_3.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19511_LC_10_17_3.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19511_LC_10_17_3.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_cmd_0__bdd_4_lut_19511_LC_10_17_3 (
            .in0(N__28013),
            .in1(N__56913),
            .in2(N__27801),
            .in3(N__57489),
            .lcout(n22147),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i26_LC_10_17_4 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i26_LC_10_17_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i26_LC_10_17_4 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i26_LC_10_17_4  (
            .in0(N__27746),
            .in1(N__50883),
            .in2(N__27778),
            .in3(N__50479),
            .lcout(cmd_rdadctmp_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55180),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i9_LC_10_17_6.C_ON=1'b0;
    defparam buf_dds0_i9_LC_10_17_6.SEQ_MODE=4'b1000;
    defparam buf_dds0_i9_LC_10_17_6.LUT_INIT=16'b0101000011001100;
    LogicCell40 buf_dds0_i9_LC_10_17_6 (
            .in0(N__52112),
            .in1(N__32337),
            .in2(N__44148),
            .in3(N__45673),
            .lcout(buf_dds0_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55180),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_5_i23_3_lut_LC_10_17_7.C_ON=1'b0;
    defparam mux_128_Mux_5_i23_3_lut_LC_10_17_7.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_5_i23_3_lut_LC_10_17_7.LUT_INIT=16'b1110111000100010;
    LogicCell40 mux_128_Mux_5_i23_3_lut_LC_10_17_7 (
            .in0(N__30045),
            .in1(N__56914),
            .in2(_gnd_net_),
            .in3(N__30204),
            .lcout(n23_adj_1513),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i20_LC_10_18_0 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i20_LC_10_18_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i20_LC_10_18_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i20_LC_10_18_0  (
            .in0(N__48953),
            .in1(N__50948),
            .in2(N__28162),
            .in3(N__28121),
            .lcout(buf_adcdata_iac_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55195),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i4_LC_10_18_1.C_ON=1'b0;
    defparam buf_device_acadc_i4_LC_10_18_1.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i4_LC_10_18_1.LUT_INIT=16'b0111010000110000;
    LogicCell40 buf_device_acadc_i4_LC_10_18_1 (
            .in0(N__52108),
            .in1(N__39240),
            .in2(N__28086),
            .in3(N__43817),
            .lcout(IAC_FLT1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55195),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i2_LC_10_18_2.C_ON=1'b0;
    defparam buf_device_acadc_i2_LC_10_18_2.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i2_LC_10_18_2.LUT_INIT=16'b0111010100100000;
    LogicCell40 buf_device_acadc_i2_LC_10_18_2 (
            .in0(N__39238),
            .in1(N__52109),
            .in2(N__44149),
            .in3(N__28046),
            .lcout(IAC_OSR1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55195),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i13_LC_10_18_3.C_ON=1'b0;
    defparam buf_dds0_i13_LC_10_18_3.SEQ_MODE=4'b1000;
    defparam buf_dds0_i13_LC_10_18_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 buf_dds0_i13_LC_10_18_3 (
            .in0(N__44850),
            .in1(N__32300),
            .in2(_gnd_net_),
            .in3(N__45677),
            .lcout(buf_dds0_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55195),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i3_LC_10_18_4.C_ON=1'b0;
    defparam buf_device_acadc_i3_LC_10_18_4.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i3_LC_10_18_4.LUT_INIT=16'b0111010100100000;
    LogicCell40 buf_device_acadc_i3_LC_10_18_4 (
            .in0(N__39239),
            .in1(N__52110),
            .in2(N__38733),
            .in3(N__28014),
            .lcout(IAC_FLT0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55195),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19551_LC_10_18_5.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19551_LC_10_18_5.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19551_LC_10_18_5.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_0__bdd_4_lut_19551_LC_10_18_5 (
            .in0(N__28211),
            .in1(N__57541),
            .in2(N__27992),
            .in3(N__56967),
            .lcout(),
            .ltout(n22189_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22189_bdd_4_lut_LC_10_18_6.C_ON=1'b0;
    defparam n22189_bdd_4_lut_LC_10_18_6.SEQ_MODE=4'b0000;
    defparam n22189_bdd_4_lut_LC_10_18_6.LUT_INIT=16'b1110010111100000;
    LogicCell40 n22189_bdd_4_lut_LC_10_18_6 (
            .in0(N__57542),
            .in1(N__27959),
            .in2(N__27943),
            .in3(N__43413),
            .lcout(n20769),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_5_i16_3_lut_LC_10_19_0.C_ON=1'b0;
    defparam mux_129_Mux_5_i16_3_lut_LC_10_19_0.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_5_i16_3_lut_LC_10_19_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_129_Mux_5_i16_3_lut_LC_10_19_0 (
            .in0(N__29509),
            .in1(N__43066),
            .in2(_gnd_net_),
            .in3(N__56968),
            .lcout(n16_adj_1489),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i1_LC_10_19_6.C_ON=1'b0;
    defparam buf_device_acadc_i1_LC_10_19_6.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i1_LC_10_19_6.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_device_acadc_i1_LC_10_19_6 (
            .in0(N__52162),
            .in1(N__39241),
            .in2(N__43534),
            .in3(N__28212),
            .lcout(IAC_OSR0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55209),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.t0off_i0_LC_11_3_0 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i0_LC_11_3_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i0_LC_11_3_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i0_LC_11_3_0  (
            .in0(_gnd_net_),
            .in1(N__30349),
            .in2(_gnd_net_),
            .in3(N__28195),
            .lcout(\ADC_VDC.genclk.t0off_0 ),
            .ltout(),
            .carryin(bfn_11_3_0_),
            .carryout(\ADC_VDC.genclk.n19410 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__30532),
            .sr(N__37444));
    defparam \ADC_VDC.genclk.t0off_i1_LC_11_3_1 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i1_LC_11_3_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i1_LC_11_3_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i1_LC_11_3_1  (
            .in0(_gnd_net_),
            .in1(N__30379),
            .in2(N__52809),
            .in3(N__28192),
            .lcout(\ADC_VDC.genclk.t0off_1 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19410 ),
            .carryout(\ADC_VDC.genclk.n19411 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__30532),
            .sr(N__37444));
    defparam \ADC_VDC.genclk.t0off_i2_LC_11_3_2 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i2_LC_11_3_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i2_LC_11_3_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i2_LC_11_3_2  (
            .in0(_gnd_net_),
            .in1(N__52754),
            .in2(N__30322),
            .in3(N__28189),
            .lcout(\ADC_VDC.genclk.t0off_2 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19411 ),
            .carryout(\ADC_VDC.genclk.n19412 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__30532),
            .sr(N__37444));
    defparam \ADC_VDC.genclk.t0off_i3_LC_11_3_3 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i3_LC_11_3_3 .SEQ_MODE=4'b1001;
    defparam \ADC_VDC.genclk.t0off_i3_LC_11_3_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i3_LC_11_3_3  (
            .in0(_gnd_net_),
            .in1(N__30232),
            .in2(N__52810),
            .in3(N__28186),
            .lcout(\ADC_VDC.genclk.t0off_3 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19412 ),
            .carryout(\ADC_VDC.genclk.n19413 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__30532),
            .sr(N__37444));
    defparam \ADC_VDC.genclk.t0off_i4_LC_11_3_4 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i4_LC_11_3_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i4_LC_11_3_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i4_LC_11_3_4  (
            .in0(_gnd_net_),
            .in1(N__52758),
            .in2(N__30367),
            .in3(N__28183),
            .lcout(\ADC_VDC.genclk.t0off_4 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19413 ),
            .carryout(\ADC_VDC.genclk.n19414 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__30532),
            .sr(N__37444));
    defparam \ADC_VDC.genclk.t0off_i5_LC_11_3_5 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i5_LC_11_3_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i5_LC_11_3_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i5_LC_11_3_5  (
            .in0(_gnd_net_),
            .in1(N__30246),
            .in2(N__52811),
            .in3(N__28180),
            .lcout(\ADC_VDC.genclk.t0off_5 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19414 ),
            .carryout(\ADC_VDC.genclk.n19415 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__30532),
            .sr(N__37444));
    defparam \ADC_VDC.genclk.t0off_i6_LC_11_3_6 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i6_LC_11_3_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i6_LC_11_3_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i6_LC_11_3_6  (
            .in0(_gnd_net_),
            .in1(N__52762),
            .in2(N__30394),
            .in3(N__28177),
            .lcout(\ADC_VDC.genclk.t0off_6 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19415 ),
            .carryout(\ADC_VDC.genclk.n19416 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__30532),
            .sr(N__37444));
    defparam \ADC_VDC.genclk.t0off_i7_LC_11_3_7 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i7_LC_11_3_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i7_LC_11_3_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i7_LC_11_3_7  (
            .in0(_gnd_net_),
            .in1(N__30306),
            .in2(N__52812),
            .in3(N__28264),
            .lcout(\ADC_VDC.genclk.t0off_7 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19416 ),
            .carryout(\ADC_VDC.genclk.n19417 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__30532),
            .sr(N__37444));
    defparam \ADC_VDC.genclk.t0off_i8_LC_11_4_0 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i8_LC_11_4_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i8_LC_11_4_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i8_LC_11_4_0  (
            .in0(_gnd_net_),
            .in1(N__30259),
            .in2(N__52750),
            .in3(N__28261),
            .lcout(\ADC_VDC.genclk.t0off_8 ),
            .ltout(),
            .carryin(bfn_11_4_0_),
            .carryout(\ADC_VDC.genclk.n19418 ),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__30528),
            .sr(N__37445));
    defparam \ADC_VDC.genclk.t0off_i9_LC_11_4_1 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i9_LC_11_4_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i9_LC_11_4_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i9_LC_11_4_1  (
            .in0(_gnd_net_),
            .in1(N__52667),
            .in2(N__30583),
            .in3(N__28258),
            .lcout(\ADC_VDC.genclk.t0off_9 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19418 ),
            .carryout(\ADC_VDC.genclk.n19419 ),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__30528),
            .sr(N__37445));
    defparam \ADC_VDC.genclk.t0off_i10_LC_11_4_2 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i10_LC_11_4_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i10_LC_11_4_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i10_LC_11_4_2  (
            .in0(_gnd_net_),
            .in1(N__30292),
            .in2(N__52747),
            .in3(N__28255),
            .lcout(\ADC_VDC.genclk.t0off_10 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19419 ),
            .carryout(\ADC_VDC.genclk.n19420 ),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__30528),
            .sr(N__37445));
    defparam \ADC_VDC.genclk.t0off_i11_LC_11_4_3 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i11_LC_11_4_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i11_LC_11_4_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i11_LC_11_4_3  (
            .in0(_gnd_net_),
            .in1(N__52655),
            .in2(N__30553),
            .in3(N__28252),
            .lcout(\ADC_VDC.genclk.t0off_11 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19420 ),
            .carryout(\ADC_VDC.genclk.n19421 ),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__30528),
            .sr(N__37445));
    defparam \ADC_VDC.genclk.t0off_i12_LC_11_4_4 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i12_LC_11_4_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i12_LC_11_4_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i12_LC_11_4_4  (
            .in0(_gnd_net_),
            .in1(N__30334),
            .in2(N__52748),
            .in3(N__28249),
            .lcout(\ADC_VDC.genclk.t0off_12 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19421 ),
            .carryout(\ADC_VDC.genclk.n19422 ),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__30528),
            .sr(N__37445));
    defparam \ADC_VDC.genclk.t0off_i13_LC_11_4_5 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i13_LC_11_4_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i13_LC_11_4_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i13_LC_11_4_5  (
            .in0(_gnd_net_),
            .in1(N__52659),
            .in2(N__30274),
            .in3(N__28246),
            .lcout(\ADC_VDC.genclk.t0off_13 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19422 ),
            .carryout(\ADC_VDC.genclk.n19423 ),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__30528),
            .sr(N__37445));
    defparam \ADC_VDC.genclk.t0off_i14_LC_11_4_6 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i14_LC_11_4_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i14_LC_11_4_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i14_LC_11_4_6  (
            .in0(_gnd_net_),
            .in1(N__30595),
            .in2(N__52749),
            .in3(N__28243),
            .lcout(\ADC_VDC.genclk.t0off_14 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19423 ),
            .carryout(\ADC_VDC.genclk.n19424 ),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__30528),
            .sr(N__37445));
    defparam \ADC_VDC.genclk.t0off_i15_LC_11_4_7 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.t0off_i15_LC_11_4_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i15_LC_11_4_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ADC_VDC.genclk.t0off_i15_LC_11_4_7  (
            .in0(N__30567),
            .in1(N__52663),
            .in2(_gnd_net_),
            .in3(N__28240),
            .lcout(\ADC_VDC.genclk.t0off_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__30528),
            .sr(N__37445));
    defparam \ADC_VDC.i1_3_lut_4_lut_LC_11_5_0 .C_ON=1'b0;
    defparam \ADC_VDC.i1_3_lut_4_lut_LC_11_5_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_3_lut_4_lut_LC_11_5_0 .LUT_INIT=16'b1010101000001000;
    LogicCell40 \ADC_VDC.i1_3_lut_4_lut_LC_11_5_0  (
            .in0(N__34290),
            .in1(N__34742),
            .in2(N__34147),
            .in3(N__34490),
            .lcout(n13073),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.adc_state_i3_LC_11_5_1 .C_ON=1'b0;
    defparam \ADC_VDC.adc_state_i3_LC_11_5_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.adc_state_i3_LC_11_5_1 .LUT_INIT=16'b0010010000001100;
    LogicCell40 \ADC_VDC.adc_state_i3_LC_11_5_1  (
            .in0(N__34113),
            .in1(N__34292),
            .in2(N__34562),
            .in3(N__34745),
            .lcout(adc_state_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32861),
            .ce(N__30508),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i12542_2_lut_LC_11_5_3 .C_ON=1'b0;
    defparam \ADC_VDC.i12542_2_lut_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i12542_2_lut_LC_11_5_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ADC_VDC.i12542_2_lut_LC_11_5_3  (
            .in0(_gnd_net_),
            .in1(N__29134),
            .in2(_gnd_net_),
            .in3(N__34289),
            .lcout(\ADC_VDC.n14900 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_2_lut_adj_31_LC_11_5_4 .C_ON=1'b0;
    defparam \ADC_VDC.i1_2_lut_adj_31_LC_11_5_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_2_lut_adj_31_LC_11_5_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \ADC_VDC.i1_2_lut_adj_31_LC_11_5_4  (
            .in0(N__34291),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34489),
            .lcout(),
            .ltout(\ADC_VDC.n20618_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_4_lut_adj_38_LC_11_5_5 .C_ON=1'b0;
    defparam \ADC_VDC.i1_4_lut_adj_38_LC_11_5_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_4_lut_adj_38_LC_11_5_5 .LUT_INIT=16'b1100010011001100;
    LogicCell40 \ADC_VDC.i1_4_lut_adj_38_LC_11_5_5  (
            .in0(N__34112),
            .in1(N__30475),
            .in2(N__28300),
            .in3(N__30469),
            .lcout(\ADC_VDC.n47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.adc_state_i0_LC_11_6_1 .C_ON=1'b0;
    defparam \ADC_VDC.adc_state_i0_LC_11_6_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.adc_state_i0_LC_11_6_1 .LUT_INIT=16'b0000000001011110;
    LogicCell40 \ADC_VDC.adc_state_i0_LC_11_6_1  (
            .in0(N__34300),
            .in1(N__34844),
            .in2(N__34563),
            .in3(N__34716),
            .lcout(\ADC_VDC.adc_state_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32873),
            .ce(N__28297),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i15997_3_lut_LC_11_6_2 .C_ON=1'b0;
    defparam \ADC_VDC.i15997_3_lut_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i15997_3_lut_LC_11_6_2 .LUT_INIT=16'b1111101001011010;
    LogicCell40 \ADC_VDC.i15997_3_lut_LC_11_6_2  (
            .in0(N__34845),
            .in1(_gnd_net_),
            .in2(N__34746),
            .in3(N__34151),
            .lcout(\ADC_VDC.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_2_lut_adj_30_LC_11_6_3 .C_ON=1'b0;
    defparam \ADC_VDC.i1_2_lut_adj_30_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_2_lut_adj_30_LC_11_6_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ADC_VDC.i1_2_lut_adj_30_LC_11_6_3  (
            .in0(_gnd_net_),
            .in1(N__34712),
            .in2(_gnd_net_),
            .in3(N__34122),
            .lcout(\ADC_VDC.n7_adj_1403 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i18107_2_lut_LC_11_6_4 .C_ON=1'b0;
    defparam \ADC_VDC.i18107_2_lut_LC_11_6_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i18107_2_lut_LC_11_6_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ADC_VDC.i18107_2_lut_LC_11_6_4  (
            .in0(N__34846),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34152),
            .lcout(\ADC_VDC.n20702 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i8_4_lut_LC_11_6_5 .C_ON=1'b0;
    defparam \ADC_VDC.i8_4_lut_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i8_4_lut_LC_11_6_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.i8_4_lut_LC_11_6_5  (
            .in0(N__28464),
            .in1(N__29271),
            .in2(N__28483),
            .in3(N__28449),
            .lcout(\ADC_VDC.n20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.i19065_4_lut_LC_11_6_6 .C_ON=1'b0;
    defparam \CLK_DDS.i19065_4_lut_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \CLK_DDS.i19065_4_lut_LC_11_6_6 .LUT_INIT=16'b1000100111001100;
    LogicCell40 \CLK_DDS.i19065_4_lut_LC_11_6_6  (
            .in0(N__28909),
            .in1(N__28774),
            .in2(N__28664),
            .in3(N__28621),
            .lcout(\CLK_DDS.n12722 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.avg_cnt_i0_LC_11_7_0 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i0_LC_11_7_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i0_LC_11_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i0_LC_11_7_0  (
            .in0(_gnd_net_),
            .in1(N__28531),
            .in2(_gnd_net_),
            .in3(N__28519),
            .lcout(\ADC_VDC.avg_cnt_0 ),
            .ltout(),
            .carryin(bfn_11_7_0_),
            .carryout(\ADC_VDC.n19399 ),
            .clk(N__32895),
            .ce(N__29178),
            .sr(N__29095));
    defparam \ADC_VDC.avg_cnt_i1_LC_11_7_1 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i1_LC_11_7_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i1_LC_11_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i1_LC_11_7_1  (
            .in0(_gnd_net_),
            .in1(N__28515),
            .in2(_gnd_net_),
            .in3(N__28501),
            .lcout(\ADC_VDC.avg_cnt_1 ),
            .ltout(),
            .carryin(\ADC_VDC.n19399 ),
            .carryout(\ADC_VDC.n19400 ),
            .clk(N__32895),
            .ce(N__29178),
            .sr(N__29095));
    defparam \ADC_VDC.avg_cnt_i2_LC_11_7_2 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i2_LC_11_7_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i2_LC_11_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i2_LC_11_7_2  (
            .in0(_gnd_net_),
            .in1(N__28498),
            .in2(_gnd_net_),
            .in3(N__28486),
            .lcout(\ADC_VDC.avg_cnt_2 ),
            .ltout(),
            .carryin(\ADC_VDC.n19400 ),
            .carryout(\ADC_VDC.n19401 ),
            .clk(N__32895),
            .ce(N__29178),
            .sr(N__29095));
    defparam \ADC_VDC.avg_cnt_i3_LC_11_7_3 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i3_LC_11_7_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i3_LC_11_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i3_LC_11_7_3  (
            .in0(_gnd_net_),
            .in1(N__28482),
            .in2(_gnd_net_),
            .in3(N__28468),
            .lcout(\ADC_VDC.avg_cnt_3 ),
            .ltout(),
            .carryin(\ADC_VDC.n19401 ),
            .carryout(\ADC_VDC.n19402 ),
            .clk(N__32895),
            .ce(N__29178),
            .sr(N__29095));
    defparam \ADC_VDC.avg_cnt_i4_LC_11_7_4 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i4_LC_11_7_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i4_LC_11_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i4_LC_11_7_4  (
            .in0(_gnd_net_),
            .in1(N__28465),
            .in2(_gnd_net_),
            .in3(N__28453),
            .lcout(\ADC_VDC.avg_cnt_4 ),
            .ltout(),
            .carryin(\ADC_VDC.n19402 ),
            .carryout(\ADC_VDC.n19403 ),
            .clk(N__32895),
            .ce(N__29178),
            .sr(N__29095));
    defparam \ADC_VDC.avg_cnt_i5_LC_11_7_5 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i5_LC_11_7_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i5_LC_11_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i5_LC_11_7_5  (
            .in0(_gnd_net_),
            .in1(N__28450),
            .in2(_gnd_net_),
            .in3(N__28438),
            .lcout(\ADC_VDC.avg_cnt_5 ),
            .ltout(),
            .carryin(\ADC_VDC.n19403 ),
            .carryout(\ADC_VDC.n19404 ),
            .clk(N__32895),
            .ce(N__29178),
            .sr(N__29095));
    defparam \ADC_VDC.avg_cnt_i6_LC_11_7_6 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i6_LC_11_7_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i6_LC_11_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i6_LC_11_7_6  (
            .in0(_gnd_net_),
            .in1(N__28435),
            .in2(_gnd_net_),
            .in3(N__28423),
            .lcout(\ADC_VDC.avg_cnt_6 ),
            .ltout(),
            .carryin(\ADC_VDC.n19404 ),
            .carryout(\ADC_VDC.n19405 ),
            .clk(N__32895),
            .ce(N__29178),
            .sr(N__29095));
    defparam \ADC_VDC.avg_cnt_i7_LC_11_7_7 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i7_LC_11_7_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i7_LC_11_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i7_LC_11_7_7  (
            .in0(_gnd_net_),
            .in1(N__29272),
            .in2(_gnd_net_),
            .in3(N__29260),
            .lcout(\ADC_VDC.avg_cnt_7 ),
            .ltout(),
            .carryin(\ADC_VDC.n19405 ),
            .carryout(\ADC_VDC.n19406 ),
            .clk(N__32895),
            .ce(N__29178),
            .sr(N__29095));
    defparam \ADC_VDC.avg_cnt_i8_LC_11_8_0 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i8_LC_11_8_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i8_LC_11_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i8_LC_11_8_0  (
            .in0(_gnd_net_),
            .in1(N__29253),
            .in2(_gnd_net_),
            .in3(N__29239),
            .lcout(\ADC_VDC.avg_cnt_8 ),
            .ltout(),
            .carryin(bfn_11_8_0_),
            .carryout(\ADC_VDC.n19407 ),
            .clk(N__32893),
            .ce(N__29177),
            .sr(N__29099));
    defparam \ADC_VDC.avg_cnt_i9_LC_11_8_1 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i9_LC_11_8_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i9_LC_11_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i9_LC_11_8_1  (
            .in0(_gnd_net_),
            .in1(N__29236),
            .in2(_gnd_net_),
            .in3(N__29224),
            .lcout(\ADC_VDC.avg_cnt_9 ),
            .ltout(),
            .carryin(\ADC_VDC.n19407 ),
            .carryout(\ADC_VDC.n19408 ),
            .clk(N__32893),
            .ce(N__29177),
            .sr(N__29099));
    defparam \ADC_VDC.avg_cnt_i10_LC_11_8_2 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i10_LC_11_8_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i10_LC_11_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i10_LC_11_8_2  (
            .in0(_gnd_net_),
            .in1(N__29221),
            .in2(_gnd_net_),
            .in3(N__29209),
            .lcout(\ADC_VDC.avg_cnt_10 ),
            .ltout(),
            .carryin(\ADC_VDC.n19408 ),
            .carryout(\ADC_VDC.n19409 ),
            .clk(N__32893),
            .ce(N__29177),
            .sr(N__29099));
    defparam \ADC_VDC.avg_cnt_i11_LC_11_8_3 .C_ON=1'b0;
    defparam \ADC_VDC.avg_cnt_i11_LC_11_8_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i11_LC_11_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i11_LC_11_8_3  (
            .in0(_gnd_net_),
            .in1(N__29203),
            .in2(_gnd_net_),
            .in3(N__29206),
            .lcout(\ADC_VDC.avg_cnt_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32893),
            .ce(N__29177),
            .sr(N__29099));
    defparam mux_128_Mux_7_i23_3_lut_LC_11_9_0.C_ON=1'b0;
    defparam mux_128_Mux_7_i23_3_lut_LC_11_9_0.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_7_i23_3_lut_LC_11_9_0.LUT_INIT=16'b1110111000100010;
    LogicCell40 mux_128_Mux_7_i23_3_lut_LC_11_9_0 (
            .in0(N__29356),
            .in1(N__56956),
            .in2(_gnd_net_),
            .in3(N__36598),
            .lcout(),
            .ltout(n23_adj_1510_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18238_4_lut_LC_11_9_1.C_ON=1'b0;
    defparam i18238_4_lut_LC_11_9_1.SEQ_MODE=4'b0000;
    defparam i18238_4_lut_LC_11_9_1.LUT_INIT=16'b0111010000110000;
    LogicCell40 i18238_4_lut_LC_11_9_1 (
            .in0(N__56957),
            .in1(N__57393),
            .in2(N__29035),
            .in3(N__41692),
            .lcout(n20833),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18215_4_lut_LC_11_9_2.C_ON=1'b0;
    defparam i18215_4_lut_LC_11_9_2.SEQ_MODE=4'b0000;
    defparam i18215_4_lut_LC_11_9_2.LUT_INIT=16'b1111101010001000;
    LogicCell40 i18215_4_lut_LC_11_9_2 (
            .in0(N__57392),
            .in1(N__29017),
            .in2(N__31150),
            .in3(N__56958),
            .lcout(n20810),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i7_LC_11_9_3.C_ON=1'b0;
    defparam buf_control_i7_LC_11_9_3.SEQ_MODE=4'b1000;
    defparam buf_control_i7_LC_11_9_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 buf_control_i7_LC_11_9_3 (
            .in0(N__29377),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(buf_control_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55084),
            .ce(N__29344),
            .sr(N__40641));
    defparam i18851_2_lut_LC_11_9_4.C_ON=1'b0;
    defparam i18851_2_lut_LC_11_9_4.SEQ_MODE=4'b0000;
    defparam i18851_2_lut_LC_11_9_4.LUT_INIT=16'b1010101000000000;
    LogicCell40 i18851_2_lut_LC_11_9_4 (
            .in0(N__57394),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51286),
            .lcout(),
            .ltout(n21050_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18824_4_lut_LC_11_9_5.C_ON=1'b0;
    defparam i18824_4_lut_LC_11_9_5.SEQ_MODE=4'b0000;
    defparam i18824_4_lut_LC_11_9_5.LUT_INIT=16'b0100000000000000;
    LogicCell40 i18824_4_lut_LC_11_9_5 (
            .in0(N__54674),
            .in1(N__47696),
            .in2(N__29347),
            .in3(N__56169),
            .lcout(n21049),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_81_LC_11_9_6.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_81_LC_11_9_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_81_LC_11_9_6.LUT_INIT=16'b1010101010001000;
    LogicCell40 i1_2_lut_3_lut_adj_81_LC_11_9_6 (
            .in0(N__54672),
            .in1(N__51285),
            .in2(_gnd_net_),
            .in3(N__54080),
            .lcout(n20081),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_287_LC_11_9_7.C_ON=1'b0;
    defparam i1_4_lut_adj_287_LC_11_9_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_287_LC_11_9_7.LUT_INIT=16'b1100110000001000;
    LogicCell40 i1_4_lut_adj_287_LC_11_9_7 (
            .in0(N__54081),
            .in1(N__49236),
            .in2(N__40621),
            .in3(N__54673),
            .lcout(n11905),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_150_LC_11_10_0.C_ON=1'b0;
    defparam i1_2_lut_adj_150_LC_11_10_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_150_LC_11_10_0.LUT_INIT=16'b0100010001000100;
    LogicCell40 i1_2_lut_adj_150_LC_11_10_0 (
            .in0(N__53509),
            .in1(N__44400),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n10508),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i6_LC_11_10_1.C_ON=1'b0;
    defparam buf_cfgRTD_i6_LC_11_10_1.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i6_LC_11_10_1.LUT_INIT=16'b1011101110001000;
    LogicCell40 buf_cfgRTD_i6_LC_11_10_1 (
            .in0(N__41527),
            .in1(N__45310),
            .in2(_gnd_net_),
            .in3(N__29296),
            .lcout(buf_cfgRTD_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55089),
            .ce(),
            .sr(_gnd_net_));
    defparam i15009_2_lut_3_lut_LC_11_10_3.C_ON=1'b0;
    defparam i15009_2_lut_3_lut_LC_11_10_3.SEQ_MODE=4'b0000;
    defparam i15009_2_lut_3_lut_LC_11_10_3.LUT_INIT=16'b0000010100000000;
    LogicCell40 i15009_2_lut_3_lut_LC_11_10_3 (
            .in0(N__29421),
            .in1(_gnd_net_),
            .in2(N__29437),
            .in3(N__29448),
            .lcout(comm_state_3_N_428_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_245_LC_11_10_4.C_ON=1'b0;
    defparam i1_4_lut_adj_245_LC_11_10_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_245_LC_11_10_4.LUT_INIT=16'b1000110010001000;
    LogicCell40 i1_4_lut_adj_245_LC_11_10_4 (
            .in0(N__54656),
            .in1(N__49237),
            .in2(N__51297),
            .in3(N__44356),
            .lcout(n11882),
            .ltout(n11882_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i4_LC_11_10_5.C_ON=1'b0;
    defparam comm_cmd_i4_LC_11_10_5.SEQ_MODE=4'b1000;
    defparam comm_cmd_i4_LC_11_10_5.LUT_INIT=16'b1000111110000000;
    LogicCell40 comm_cmd_i4_LC_11_10_5 (
            .in0(N__35662),
            .in1(N__30989),
            .in2(N__29275),
            .in3(N__29449),
            .lcout(comm_cmd_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55089),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_302_LC_11_10_6.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_302_LC_11_10_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_302_LC_11_10_6.LUT_INIT=16'b1111111111011101;
    LogicCell40 i1_2_lut_3_lut_adj_302_LC_11_10_6 (
            .in0(N__29447),
            .in1(N__29420),
            .in2(_gnd_net_),
            .in3(N__29432),
            .lcout(n20602),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i6_LC_11_10_7.C_ON=1'b0;
    defparam comm_cmd_i6_LC_11_10_7.SEQ_MODE=4'b1000;
    defparam comm_cmd_i6_LC_11_10_7.LUT_INIT=16'b1100000010101010;
    LogicCell40 comm_cmd_i6_LC_11_10_7 (
            .in0(N__29436),
            .in1(N__30990),
            .in2(N__35811),
            .in3(N__30928),
            .lcout(comm_cmd_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55089),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i2_LC_11_11_0.C_ON=1'b0;
    defparam comm_cmd_i2_LC_11_11_0.SEQ_MODE=4'b1000;
    defparam comm_cmd_i2_LC_11_11_0.LUT_INIT=16'b1011100000110000;
    LogicCell40 comm_cmd_i2_LC_11_11_0 (
            .in0(N__30999),
            .in1(N__30929),
            .in2(N__47701),
            .in3(N__35449),
            .lcout(comm_cmd_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55097),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i5_LC_11_11_1.C_ON=1'b0;
    defparam comm_cmd_i5_LC_11_11_1.SEQ_MODE=4'b1000;
    defparam comm_cmd_i5_LC_11_11_1.LUT_INIT=16'b1101010110000000;
    LogicCell40 comm_cmd_i5_LC_11_11_1 (
            .in0(N__30930),
            .in1(N__31000),
            .in2(N__38023),
            .in3(N__29422),
            .lcout(comm_cmd_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55097),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_3_lut_LC_11_11_2.C_ON=1'b0;
    defparam i3_3_lut_LC_11_11_2.SEQ_MODE=4'b0000;
    defparam i3_3_lut_LC_11_11_2.LUT_INIT=16'b0000110000000000;
    LogicCell40 i3_3_lut_LC_11_11_2 (
            .in0(_gnd_net_),
            .in1(N__51293),
            .in2(N__53531),
            .in3(N__46588),
            .lcout(),
            .ltout(n8_adj_1522_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_237_LC_11_11_3.C_ON=1'b0;
    defparam i1_4_lut_adj_237_LC_11_11_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_237_LC_11_11_3.LUT_INIT=16'b1100110010000000;
    LogicCell40 i1_4_lut_adj_237_LC_11_11_3 (
            .in0(N__29482),
            .in1(N__49238),
            .in2(N__29407),
            .in3(N__54657),
            .lcout(n12214),
            .ltout(n12214_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i2_LC_11_11_4.C_ON=1'b0;
    defparam comm_buf_6__i2_LC_11_11_4.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i2_LC_11_11_4.LUT_INIT=16'b0100111101000000;
    LogicCell40 comm_buf_6__i2_LC_11_11_4 (
            .in0(N__54659),
            .in1(N__35448),
            .in2(N__29404),
            .in3(N__35082),
            .lcout(comm_buf_6_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55097),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i3_LC_11_11_5.C_ON=1'b0;
    defparam comm_buf_6__i3_LC_11_11_5.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i3_LC_11_11_5.LUT_INIT=16'b0011000010101010;
    LogicCell40 comm_buf_6__i3_LC_11_11_5 (
            .in0(N__33075),
            .in1(N__54661),
            .in2(N__35568),
            .in3(N__29471),
            .lcout(comm_buf_6_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55097),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i13_LC_11_11_6.C_ON=1'b0;
    defparam buf_dds1_i13_LC_11_11_6.SEQ_MODE=4'b1000;
    defparam buf_dds1_i13_LC_11_11_6.LUT_INIT=16'b1111010111001100;
    LogicCell40 buf_dds1_i13_LC_11_11_6 (
            .in0(N__54658),
            .in1(N__29397),
            .in2(N__44851),
            .in3(N__45912),
            .lcout(buf_dds1_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55097),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i1_LC_11_11_7.C_ON=1'b0;
    defparam comm_buf_6__i1_LC_11_11_7.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i1_LC_11_11_7.LUT_INIT=16'b0011000010101010;
    LogicCell40 comm_buf_6__i1_LC_11_11_7 (
            .in0(N__47172),
            .in1(N__54660),
            .in2(N__35978),
            .in3(N__29470),
            .lcout(comm_buf_6_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55097),
            .ce(),
            .sr(_gnd_net_));
    defparam n22075_bdd_4_lut_LC_11_12_0.C_ON=1'b0;
    defparam n22075_bdd_4_lut_LC_11_12_0.SEQ_MODE=4'b0000;
    defparam n22075_bdd_4_lut_LC_11_12_0.LUT_INIT=16'b1100110010111000;
    LogicCell40 n22075_bdd_4_lut_LC_11_12_0 (
            .in0(N__29557),
            .in1(N__29536),
            .in2(N__43104),
            .in3(N__57441),
            .lcout(n22078),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i5_LC_11_12_1.C_ON=1'b0;
    defparam buf_dds1_i5_LC_11_12_1.SEQ_MODE=4'b1000;
    defparam buf_dds1_i5_LC_11_12_1.LUT_INIT=16'b1111001110101010;
    LogicCell40 buf_dds1_i5_LC_11_12_1 (
            .in0(N__29498),
            .in1(N__54665),
            .in2(N__50137),
            .in3(N__45891),
            .lcout(buf_dds1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55106),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i0_LC_11_12_2.C_ON=1'b0;
    defparam comm_buf_6__i0_LC_11_12_2.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i0_LC_11_12_2.LUT_INIT=16'b0100010011110000;
    LogicCell40 comm_buf_6__i0_LC_11_12_2 (
            .in0(N__54662),
            .in1(N__36254),
            .in2(N__38076),
            .in3(N__29472),
            .lcout(comm_buf_6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55106),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_adj_236_LC_11_12_3.C_ON=1'b0;
    defparam i2_2_lut_adj_236_LC_11_12_3.SEQ_MODE=4'b0000;
    defparam i2_2_lut_adj_236_LC_11_12_3.LUT_INIT=16'b1100110000000000;
    LogicCell40 i2_2_lut_adj_236_LC_11_12_3 (
            .in0(_gnd_net_),
            .in1(N__50097),
            .in2(_gnd_net_),
            .in3(N__54094),
            .lcout(n7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i7_LC_11_12_4.C_ON=1'b0;
    defparam comm_buf_6__i7_LC_11_12_4.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i7_LC_11_12_4.LUT_INIT=16'b0100010011110000;
    LogicCell40 comm_buf_6__i7_LC_11_12_4 (
            .in0(N__54664),
            .in1(N__36895),
            .in2(N__33960),
            .in3(N__29476),
            .lcout(comm_buf_6_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55106),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i6_LC_11_12_5.C_ON=1'b0;
    defparam comm_buf_6__i6_LC_11_12_5.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i6_LC_11_12_5.LUT_INIT=16'b0111001001010000;
    LogicCell40 comm_buf_6__i6_LC_11_12_5 (
            .in0(N__29475),
            .in1(N__54667),
            .in2(N__33166),
            .in3(N__35806),
            .lcout(comm_buf_6_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55106),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i5_LC_11_12_6.C_ON=1'b0;
    defparam comm_buf_6__i5_LC_11_12_6.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i5_LC_11_12_6.LUT_INIT=16'b0101000011001100;
    LogicCell40 comm_buf_6__i5_LC_11_12_6 (
            .in0(N__54663),
            .in1(N__38259),
            .in2(N__38016),
            .in3(N__29474),
            .lcout(comm_buf_6_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55106),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i4_LC_11_12_7.C_ON=1'b0;
    defparam comm_buf_6__i4_LC_11_12_7.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i4_LC_11_12_7.LUT_INIT=16'b0100010011100100;
    LogicCell40 comm_buf_6__i4_LC_11_12_7 (
            .in0(N__29473),
            .in1(N__46734),
            .in2(N__35663),
            .in3(N__54666),
            .lcout(comm_buf_6_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55106),
            .ce(),
            .sr(_gnd_net_));
    defparam i14137_4_lut_LC_11_13_0.C_ON=1'b0;
    defparam i14137_4_lut_LC_11_13_0.SEQ_MODE=4'b0000;
    defparam i14137_4_lut_LC_11_13_0.LUT_INIT=16'b1101111100010011;
    LogicCell40 i14137_4_lut_LC_11_13_0 (
            .in0(N__31489),
            .in1(N__32155),
            .in2(N__30462),
            .in3(N__38899),
            .lcout(),
            .ltout(n16539_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_state_i0_LC_11_13_1.C_ON=1'b0;
    defparam eis_state_i0_LC_11_13_1.SEQ_MODE=4'b1010;
    defparam eis_state_i0_LC_11_13_1.LUT_INIT=16'b1111101000010001;
    LogicCell40 eis_state_i0_LC_11_13_1 (
            .in0(N__37582),
            .in1(N__32159),
            .in2(N__29650),
            .in3(N__31837),
            .lcout(eis_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVeis_state_i0C_net),
            .ce(N__30406),
            .sr(N__32099));
    defparam i24_4_lut_LC_11_13_3.C_ON=1'b0;
    defparam i24_4_lut_LC_11_13_3.SEQ_MODE=4'b0000;
    defparam i24_4_lut_LC_11_13_3.LUT_INIT=16'b0110111001100010;
    LogicCell40 i24_4_lut_LC_11_13_3 (
            .in0(N__37581),
            .in1(N__32158),
            .in2(N__39122),
            .in3(N__46976),
            .lcout(),
            .ltout(n17_adj_1601_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_state_i1_LC_11_13_4.C_ON=1'b0;
    defparam eis_state_i1_LC_11_13_4.SEQ_MODE=4'b1010;
    defparam eis_state_i1_LC_11_13_4.LUT_INIT=16'b1111000011110010;
    LogicCell40 eis_state_i1_LC_11_13_4 (
            .in0(N__39106),
            .in1(N__37583),
            .in2(N__29647),
            .in3(N__29644),
            .lcout(eis_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVeis_state_i0C_net),
            .ce(N__30406),
            .sr(N__32099));
    defparam i1_2_lut_adj_211_LC_11_13_5.C_ON=1'b0;
    defparam i1_2_lut_adj_211_LC_11_13_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_211_LC_11_13_5.LUT_INIT=16'b1111111100110011;
    LogicCell40 i1_2_lut_adj_211_LC_11_13_5 (
            .in0(_gnd_net_),
            .in1(N__30454),
            .in2(_gnd_net_),
            .in3(N__31488),
            .lcout(n16547),
            .ltout(n16547_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i34_3_lut_LC_11_13_6.C_ON=1'b0;
    defparam i34_3_lut_LC_11_13_6.SEQ_MODE=4'b0000;
    defparam i34_3_lut_LC_11_13_6.LUT_INIT=16'b1010101011110000;
    LogicCell40 i34_3_lut_LC_11_13_6 (
            .in0(N__46975),
            .in1(_gnd_net_),
            .in2(N__29638),
            .in3(N__37580),
            .lcout(),
            .ltout(n13_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_state_i2_LC_11_13_7.C_ON=1'b0;
    defparam eis_state_i2_LC_11_13_7.SEQ_MODE=4'b1010;
    defparam eis_state_i2_LC_11_13_7.LUT_INIT=16'b1110110001100100;
    LogicCell40 eis_state_i2_LC_11_13_7 (
            .in0(N__39105),
            .in1(N__32160),
            .in2(N__29635),
            .in3(N__37528),
            .lcout(eis_end_N_716),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVeis_state_i0C_net),
            .ce(N__30406),
            .sr(N__32099));
    defparam mux_129_Mux_6_i26_3_lut_LC_11_14_0.C_ON=1'b0;
    defparam mux_129_Mux_6_i26_3_lut_LC_11_14_0.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_6_i26_3_lut_LC_11_14_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_129_Mux_6_i26_3_lut_LC_11_14_0 (
            .in0(N__56887),
            .in1(N__31222),
            .in2(_gnd_net_),
            .in3(N__47413),
            .lcout(n26_adj_1495),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19345_LC_11_14_3.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19345_LC_11_14_3.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19345_LC_11_14_3.LUT_INIT=16'b1110010010101010;
    LogicCell40 comm_cmd_1__bdd_4_lut_19345_LC_11_14_3 (
            .in0(N__57522),
            .in1(N__29632),
            .in2(N__29620),
            .in3(N__47699),
            .lcout(),
            .ltout(n21937_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n21937_bdd_4_lut_LC_11_14_4.C_ON=1'b0;
    defparam n21937_bdd_4_lut_LC_11_14_4.SEQ_MODE=4'b0000;
    defparam n21937_bdd_4_lut_LC_11_14_4.LUT_INIT=16'b1111010010100100;
    LogicCell40 n21937_bdd_4_lut_LC_11_14_4 (
            .in0(N__47700),
            .in1(N__36088),
            .in2(N__29590),
            .in3(N__29587),
            .lcout(),
            .ltout(n21940_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1542274_i1_3_lut_LC_11_14_5.C_ON=1'b0;
    defparam i1542274_i1_3_lut_LC_11_14_5.SEQ_MODE=4'b0000;
    defparam i1542274_i1_3_lut_LC_11_14_5.LUT_INIT=16'b1111110000110000;
    LogicCell40 i1542274_i1_3_lut_LC_11_14_5 (
            .in0(_gnd_net_),
            .in1(N__56273),
            .in2(N__29686),
            .in3(N__29656),
            .lcout(),
            .ltout(n30_adj_1490_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i6_LC_11_14_6.C_ON=1'b0;
    defparam comm_buf_1__i6_LC_11_14_6.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i6_LC_11_14_6.LUT_INIT=16'b1101100011011000;
    LogicCell40 comm_buf_1__i6_LC_11_14_6 (
            .in0(N__54051),
            .in1(N__35812),
            .in2(N__29683),
            .in3(_gnd_net_),
            .lcout(comm_buf_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55126),
            .ce(N__38557),
            .sr(N__36791));
    defparam buf_dds1_i4_LC_11_15_0.C_ON=1'b0;
    defparam buf_dds1_i4_LC_11_15_0.SEQ_MODE=4'b1000;
    defparam buf_dds1_i4_LC_11_15_0.LUT_INIT=16'b1000101010000000;
    LogicCell40 buf_dds1_i4_LC_11_15_0 (
            .in0(N__46006),
            .in1(N__46666),
            .in2(N__45913),
            .in3(N__36144),
            .lcout(buf_dds1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55138),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i12_LC_11_15_2.C_ON=1'b0;
    defparam buf_dds0_i12_LC_11_15_2.SEQ_MODE=4'b1000;
    defparam buf_dds0_i12_LC_11_15_2.LUT_INIT=16'b1100110010101010;
    LogicCell40 buf_dds0_i12_LC_11_15_2 (
            .in0(N__33857),
            .in1(N__42143),
            .in2(_gnd_net_),
            .in3(N__45657),
            .lcout(buf_dds0_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55138),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i10_LC_11_15_3.C_ON=1'b0;
    defparam buf_dds1_i10_LC_11_15_3.SEQ_MODE=4'b1000;
    defparam buf_dds1_i10_LC_11_15_3.LUT_INIT=16'b1110001000000000;
    LogicCell40 buf_dds1_i10_LC_11_15_3 (
            .in0(N__30185),
            .in1(N__45896),
            .in2(N__38731),
            .in3(N__46005),
            .lcout(buf_dds1_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55138),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i8_LC_11_15_4.C_ON=1'b0;
    defparam acadc_skipCount_i8_LC_11_15_4.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i8_LC_11_15_4.LUT_INIT=16'b0101110100001000;
    LogicCell40 acadc_skipCount_i8_LC_11_15_4 (
            .in0(N__39328),
            .in1(N__43520),
            .in2(N__52193),
            .in3(N__31533),
            .lcout(acadc_skipCount_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55138),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19482_LC_11_15_5.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19482_LC_11_15_5.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19482_LC_11_15_5.LUT_INIT=16'b1110010010101010;
    LogicCell40 comm_cmd_1__bdd_4_lut_19482_LC_11_15_5 (
            .in0(N__57521),
            .in1(N__29680),
            .in2(N__29674),
            .in3(N__47697),
            .lcout(),
            .ltout(n22111_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22111_bdd_4_lut_LC_11_15_6.C_ON=1'b0;
    defparam n22111_bdd_4_lut_LC_11_15_6.SEQ_MODE=4'b0000;
    defparam n22111_bdd_4_lut_LC_11_15_6.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22111_bdd_4_lut_LC_11_15_6 (
            .in0(N__47698),
            .in1(N__31905),
            .in2(N__29659),
            .in3(N__41722),
            .lcout(n22114),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i6_LC_11_15_7.C_ON=1'b0;
    defparam acadc_skipCount_i6_LC_11_15_7.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i6_LC_11_15_7.LUT_INIT=16'b0011000010101010;
    LogicCell40 acadc_skipCount_i6_LC_11_15_7 (
            .in0(N__31906),
            .in1(N__52177),
            .in2(N__51429),
            .in3(N__39327),
            .lcout(acadc_skipCount_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55138),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_4_lut_LC_11_16_0.C_ON=1'b0;
    defparam i1_3_lut_4_lut_LC_11_16_0.SEQ_MODE=4'b0000;
    defparam i1_3_lut_4_lut_LC_11_16_0.LUT_INIT=16'b0000000000100011;
    LogicCell40 i1_3_lut_4_lut_LC_11_16_0 (
            .in0(N__37593),
            .in1(N__32156),
            .in2(N__39151),
            .in3(N__32067),
            .lcout(n13443),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6372_3_lut_LC_11_16_1.C_ON=1'b0;
    defparam i6372_3_lut_LC_11_16_1.SEQ_MODE=4'b0000;
    defparam i6372_3_lut_LC_11_16_1.LUT_INIT=16'b1100110010101010;
    LogicCell40 i6372_3_lut_LC_11_16_1 (
            .in0(N__42596),
            .in1(N__42459),
            .in2(_gnd_net_),
            .in3(N__43295),
            .lcout(n8_adj_1536),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i5_LC_11_16_2.C_ON=1'b0;
    defparam buf_control_i5_LC_11_16_2.SEQ_MODE=4'b1000;
    defparam buf_control_i5_LC_11_16_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 buf_control_i5_LC_11_16_2 (
            .in0(N__44847),
            .in1(N__43871),
            .in2(_gnd_net_),
            .in3(N__30041),
            .lcout(AMPV_POW),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55151),
            .ce(),
            .sr(_gnd_net_));
    defparam i19145_2_lut_3_lut_LC_11_16_3.C_ON=1'b0;
    defparam i19145_2_lut_3_lut_LC_11_16_3.SEQ_MODE=4'b0000;
    defparam i19145_2_lut_3_lut_LC_11_16_3.LUT_INIT=16'b0000000000010001;
    LogicCell40 i19145_2_lut_3_lut_LC_11_16_3 (
            .in0(N__32068),
            .in1(N__39141),
            .in2(_gnd_net_),
            .in3(N__32180),
            .lcout(n20757),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.DTRIG_39_LC_11_16_4 .C_ON=1'b0;
    defparam \ADC_IAC.DTRIG_39_LC_11_16_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.DTRIG_39_LC_11_16_4 .LUT_INIT=16'b1111111000001000;
    LogicCell40 \ADC_IAC.DTRIG_39_LC_11_16_4  (
            .in0(N__30022),
            .in1(N__29949),
            .in2(N__50952),
            .in3(N__31861),
            .lcout(acadc_dtrig_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55151),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_rst_327_LC_11_16_5.C_ON=1'b0;
    defparam acadc_rst_327_LC_11_16_5.SEQ_MODE=4'b1000;
    defparam acadc_rst_327_LC_11_16_5.LUT_INIT=16'b1111000010101010;
    LogicCell40 acadc_rst_327_LC_11_16_5 (
            .in0(N__32069),
            .in1(_gnd_net_),
            .in2(N__38730),
            .in3(N__29886),
            .lcout(acadc_rst),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55151),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.DTRIG_39_LC_11_16_6 .C_ON=1'b0;
    defparam \ADC_VAC.DTRIG_39_LC_11_16_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.DTRIG_39_LC_11_16_6 .LUT_INIT=16'b1111111000001000;
    LogicCell40 \ADC_VAC.DTRIG_39_LC_11_16_6  (
            .in0(N__29863),
            .in1(N__29794),
            .in2(N__48335),
            .in3(N__31885),
            .lcout(acadc_dtrig_v),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55151),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i6_LC_11_16_7.C_ON=1'b0;
    defparam buf_device_acadc_i6_LC_11_16_7.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i6_LC_11_16_7.LUT_INIT=16'b1011101110001000;
    LogicCell40 buf_device_acadc_i6_LC_11_16_7 (
            .in0(N__44848),
            .in1(N__39205),
            .in2(_gnd_net_),
            .in3(N__29705),
            .lcout(VAC_OSR1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55151),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_126_LC_11_17_0.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_126_LC_11_17_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_126_LC_11_17_0.LUT_INIT=16'b0001000100000000;
    LogicCell40 i1_2_lut_3_lut_adj_126_LC_11_17_0 (
            .in0(N__31884),
            .in1(N__31859),
            .in2(_gnd_net_),
            .in3(N__38898),
            .lcout(),
            .ltout(n4_adj_1473_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19069_4_lut_LC_11_17_1.C_ON=1'b0;
    defparam i19069_4_lut_LC_11_17_1.SEQ_MODE=4'b0000;
    defparam i19069_4_lut_LC_11_17_1.LUT_INIT=16'b0100000001110111;
    LogicCell40 i19069_4_lut_LC_11_17_1 (
            .in0(N__37595),
            .in1(N__39108),
            .in2(N__30208),
            .in3(N__32157),
            .lcout(n20529),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i14975_2_lut_LC_11_17_2.C_ON=1'b0;
    defparam i14975_2_lut_LC_11_17_2.SEQ_MODE=4'b0000;
    defparam i14975_2_lut_LC_11_17_2.LUT_INIT=16'b1111111111001100;
    LogicCell40 i14975_2_lut_LC_11_17_2 (
            .in0(_gnd_net_),
            .in1(N__31882),
            .in2(_gnd_net_),
            .in3(N__31858),
            .lcout(n17357),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_269_LC_11_17_3.C_ON=1'b0;
    defparam i1_2_lut_adj_269_LC_11_17_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_269_LC_11_17_3.LUT_INIT=16'b1010101000000000;
    LogicCell40 i1_2_lut_adj_269_LC_11_17_3 (
            .in0(N__37594),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39107),
            .lcout(n35),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i10_LC_11_17_4.C_ON=1'b0;
    defparam buf_dds0_i10_LC_11_17_4.SEQ_MODE=4'b1000;
    defparam buf_dds0_i10_LC_11_17_4.LUT_INIT=16'b0101000011001100;
    LogicCell40 buf_dds0_i10_LC_11_17_4 (
            .in0(N__52176),
            .in1(N__32366),
            .in2(N__38732),
            .in3(N__45656),
            .lcout(buf_dds0_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55166),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_61_i14_2_lut_LC_11_17_5.C_ON=1'b0;
    defparam equal_61_i14_2_lut_LC_11_17_5.SEQ_MODE=4'b0000;
    defparam equal_61_i14_2_lut_LC_11_17_5.LUT_INIT=16'b0011001111001100;
    LogicCell40 equal_61_i14_2_lut_LC_11_17_5 (
            .in0(_gnd_net_),
            .in1(N__33700),
            .in2(_gnd_net_),
            .in3(N__30203),
            .lcout(n14_adj_1498),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_LC_11_17_6.C_ON=1'b0;
    defparam i2_4_lut_LC_11_17_6.SEQ_MODE=4'b0000;
    defparam i2_4_lut_LC_11_17_6.LUT_INIT=16'b0111110110111110;
    LogicCell40 i2_4_lut_LC_11_17_6 (
            .in0(N__33676),
            .in1(N__36948),
            .in2(N__33634),
            .in3(N__36563),
            .lcout(n18_adj_1587),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22147_bdd_4_lut_LC_11_17_7.C_ON=1'b0;
    defparam n22147_bdd_4_lut_LC_11_17_7.SEQ_MODE=4'b0000;
    defparam n22147_bdd_4_lut_LC_11_17_7.LUT_INIT=16'b1100110010111000;
    LogicCell40 n22147_bdd_4_lut_LC_11_17_7 (
            .in0(N__30186),
            .in1(N__30163),
            .in2(N__32370),
            .in3(N__57531),
            .lcout(n22150),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18095_4_lut_LC_11_18_0.C_ON=1'b0;
    defparam i18095_4_lut_LC_11_18_0.SEQ_MODE=4'b0000;
    defparam i18095_4_lut_LC_11_18_0.LUT_INIT=16'b1111111010101110;
    LogicCell40 i18095_4_lut_LC_11_18_0 (
            .in0(N__32094),
            .in1(N__32161),
            .in2(N__39157),
            .in3(N__37603),
            .lcout(),
            .ltout(n20690_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_trig_300_LC_11_18_1.C_ON=1'b0;
    defparam acadc_trig_300_LC_11_18_1.SEQ_MODE=4'b1000;
    defparam acadc_trig_300_LC_11_18_1.LUT_INIT=16'b1111010000000100;
    LogicCell40 acadc_trig_300_LC_11_18_1 (
            .in0(N__32163),
            .in1(N__39156),
            .in2(N__30145),
            .in3(N__30133),
            .lcout(acadc_trig),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVacadc_trig_300C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_end_299_LC_11_18_5.C_ON=1'b0;
    defparam eis_end_299_LC_11_18_5.SEQ_MODE=4'b1000;
    defparam eis_end_299_LC_11_18_5.LUT_INIT=16'b1110001011110000;
    LogicCell40 eis_end_299_LC_11_18_5 (
            .in0(N__32164),
            .in1(N__32095),
            .in2(N__30099),
            .in3(N__30106),
            .lcout(eis_end),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVacadc_trig_300C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_4_lut_adj_234_LC_11_18_6.C_ON=1'b0;
    defparam i24_4_lut_adj_234_LC_11_18_6.SEQ_MODE=4'b0000;
    defparam i24_4_lut_adj_234_LC_11_18_6.LUT_INIT=16'b1111110010101100;
    LogicCell40 i24_4_lut_adj_234_LC_11_18_6 (
            .in0(N__30461),
            .in1(N__30415),
            .in2(N__37605),
            .in3(N__38941),
            .lcout(),
            .ltout(n11_adj_1620_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19112_3_lut_LC_11_18_7.C_ON=1'b0;
    defparam i19112_3_lut_LC_11_18_7.SEQ_MODE=4'b0000;
    defparam i19112_3_lut_LC_11_18_7.LUT_INIT=16'b0101111111111111;
    LogicCell40 i19112_3_lut_LC_11_18_7 (
            .in0(N__32162),
            .in1(_gnd_net_),
            .in2(N__30409),
            .in3(N__39152),
            .lcout(n11730),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_187_i9_2_lut_3_lut_LC_11_19_7.C_ON=1'b0;
    defparam equal_187_i9_2_lut_3_lut_LC_11_19_7.SEQ_MODE=4'b0000;
    defparam equal_187_i9_2_lut_3_lut_LC_11_19_7.LUT_INIT=16'b1111111110111011;
    LogicCell40 equal_187_i9_2_lut_3_lut_LC_11_19_7 (
            .in0(N__57540),
            .in1(N__56965),
            .in2(_gnd_net_),
            .in3(N__47695),
            .lcout(n9_adj_1407),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i19095_2_lut_LC_12_3_4 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i19095_2_lut_LC_12_3_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i19095_2_lut_LC_12_3_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \ADC_VDC.genclk.i19095_2_lut_LC_12_3_4  (
            .in0(_gnd_net_),
            .in1(N__34962),
            .in2(_gnd_net_),
            .in3(N__34930),
            .lcout(\ADC_VDC.genclk.n14695 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i19040_4_lut_LC_12_4_0 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i19040_4_lut_LC_12_4_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i19040_4_lut_LC_12_4_0 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \ADC_VDC.genclk.i19040_4_lut_LC_12_4_0  (
            .in0(N__30390),
            .in1(N__30378),
            .in2(N__30366),
            .in3(N__30348),
            .lcout(),
            .ltout(\ADC_VDC.genclk.n21169_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i18722_4_lut_LC_12_4_1 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i18722_4_lut_LC_12_4_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i18722_4_lut_LC_12_4_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i18722_4_lut_LC_12_4_1  (
            .in0(N__30538),
            .in1(N__30220),
            .in2(N__30337),
            .in3(N__30280),
            .lcout(\ADC_VDC.genclk.n21167 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i11_4_lut_LC_12_4_2 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i11_4_lut_LC_12_4_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i11_4_lut_LC_12_4_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i11_4_lut_LC_12_4_2  (
            .in0(N__30333),
            .in1(N__30318),
            .in2(N__30307),
            .in3(N__30291),
            .lcout(\ADC_VDC.genclk.n27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i10_4_lut_LC_12_4_3 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i10_4_lut_LC_12_4_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i10_4_lut_LC_12_4_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i10_4_lut_LC_12_4_3  (
            .in0(N__30270),
            .in1(N__30258),
            .in2(N__30247),
            .in3(N__30231),
            .lcout(\ADC_VDC.genclk.n26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i12_4_lut_LC_12_4_4 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i12_4_lut_LC_12_4_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i12_4_lut_LC_12_4_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i12_4_lut_LC_12_4_4  (
            .in0(N__30594),
            .in1(N__30579),
            .in2(N__30568),
            .in3(N__30549),
            .lcout(\ADC_VDC.genclk.n28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i19072_2_lut_LC_12_4_5 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i19072_2_lut_LC_12_4_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i19072_2_lut_LC_12_4_5 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \ADC_VDC.genclk.i19072_2_lut_LC_12_4_5  (
            .in0(N__34935),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34963),
            .lcout(\ADC_VDC.genclk.n11721 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i19088_4_lut_LC_12_5_0 .C_ON=1'b0;
    defparam \ADC_VDC.i19088_4_lut_LC_12_5_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i19088_4_lut_LC_12_5_0 .LUT_INIT=16'b1000101010101010;
    LogicCell40 \ADC_VDC.i19088_4_lut_LC_12_5_0  (
            .in0(N__34294),
            .in1(N__34485),
            .in2(N__34877),
            .in3(N__30637),
            .lcout(\ADC_VDC.n4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i19137_4_lut_LC_12_5_2 .C_ON=1'b0;
    defparam \ADC_VDC.i19137_4_lut_LC_12_5_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i19137_4_lut_LC_12_5_2 .LUT_INIT=16'b1101110011011111;
    LogicCell40 \ADC_VDC.i19137_4_lut_LC_12_5_2  (
            .in0(N__30624),
            .in1(N__34487),
            .in2(N__34356),
            .in3(N__30754),
            .lcout(\ADC_VDC.n17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i7713_3_lut_4_lut_LC_12_5_4 .C_ON=1'b0;
    defparam \ADC_VDC.i7713_3_lut_4_lut_LC_12_5_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i7713_3_lut_4_lut_LC_12_5_4 .LUT_INIT=16'b0101001011011010;
    LogicCell40 \ADC_VDC.i7713_3_lut_4_lut_LC_12_5_4  (
            .in0(N__34743),
            .in1(N__34158),
            .in2(N__34878),
            .in3(N__30772),
            .lcout(),
            .ltout(\ADC_VDC.n10112_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_4_lut_4_lut_LC_12_5_5 .C_ON=1'b0;
    defparam \ADC_VDC.i1_4_lut_4_lut_LC_12_5_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_4_lut_4_lut_LC_12_5_5 .LUT_INIT=16'b1011101011111110;
    LogicCell40 \ADC_VDC.i1_4_lut_4_lut_LC_12_5_5  (
            .in0(N__34486),
            .in1(N__34295),
            .in2(N__30511),
            .in3(N__30625),
            .lcout(\ADC_VDC.n12793 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.adc_state_i2_LC_12_5_6 .C_ON=1'b0;
    defparam \ADC_VDC.adc_state_i2_LC_12_5_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.adc_state_i2_LC_12_5_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ADC_VDC.adc_state_i2_LC_12_5_6  (
            .in0(N__34744),
            .in1(N__34488),
            .in2(_gnd_net_),
            .in3(N__34159),
            .lcout(adc_state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32778),
            .ce(N__30499),
            .sr(N__30493));
    defparam \ADC_VDC.i1_4_lut_adj_37_LC_12_5_7 .C_ON=1'b0;
    defparam \ADC_VDC.i1_4_lut_adj_37_LC_12_5_7 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_4_lut_adj_37_LC_12_5_7 .LUT_INIT=16'b1111001011111110;
    LogicCell40 \ADC_VDC.i1_4_lut_adj_37_LC_12_5_7  (
            .in0(N__30481),
            .in1(N__34293),
            .in2(N__34561),
            .in3(N__30623),
            .lcout(\ADC_VDC.n72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i18115_2_lut_LC_12_6_0 .C_ON=1'b0;
    defparam \ADC_VDC.i18115_2_lut_LC_12_6_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i18115_2_lut_LC_12_6_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ADC_VDC.i18115_2_lut_LC_12_6_0  (
            .in0(_gnd_net_),
            .in1(N__34741),
            .in2(_gnd_net_),
            .in3(N__30770),
            .lcout(\ADC_VDC.n20710 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i2_3_lut_LC_12_6_1 .C_ON=1'b0;
    defparam \ADC_VDC.i2_3_lut_LC_12_6_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i2_3_lut_LC_12_6_1 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \ADC_VDC.i2_3_lut_LC_12_6_1  (
            .in0(N__32435),
            .in1(N__32930),
            .in2(_gnd_net_),
            .in3(N__32951),
            .lcout(\ADC_VDC.n20490 ),
            .ltout(\ADC_VDC.n20490_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_2_lut_adj_32_LC_12_6_2 .C_ON=1'b0;
    defparam \ADC_VDC.i1_2_lut_adj_32_LC_12_6_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_2_lut_adj_32_LC_12_6_2 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \ADC_VDC.i1_2_lut_adj_32_LC_12_6_2  (
            .in0(N__32509),
            .in1(_gnd_net_),
            .in2(N__30688),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\ADC_VDC.n11251_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i4_4_lut_adj_34_LC_12_6_3 .C_ON=1'b0;
    defparam \ADC_VDC.i4_4_lut_adj_34_LC_12_6_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i4_4_lut_adj_34_LC_12_6_3 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \ADC_VDC.i4_4_lut_adj_34_LC_12_6_3  (
            .in0(N__32463),
            .in1(N__32566),
            .in2(N__30685),
            .in3(N__32546),
            .lcout(\ADC_VDC.n15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i5_3_lut_LC_12_6_4 .C_ON=1'b0;
    defparam \ADC_VDC.i5_3_lut_LC_12_6_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i5_3_lut_LC_12_6_4 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \ADC_VDC.i5_3_lut_LC_12_6_4  (
            .in0(N__32952),
            .in1(N__32931),
            .in2(_gnd_net_),
            .in3(N__30778),
            .lcout(),
            .ltout(\ADC_VDC.n20523_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i18909_4_lut_LC_12_6_5 .C_ON=1'b0;
    defparam \ADC_VDC.i18909_4_lut_LC_12_6_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i18909_4_lut_LC_12_6_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \ADC_VDC.i18909_4_lut_LC_12_6_5  (
            .in0(N__32464),
            .in1(N__34307),
            .in2(N__30682),
            .in3(N__32632),
            .lcout(\ADC_VDC.n21178 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i18807_4_lut_LC_12_6_6 .C_ON=1'b0;
    defparam \ADC_VDC.i18807_4_lut_LC_12_6_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i18807_4_lut_LC_12_6_6 .LUT_INIT=16'b1111000010000000;
    LogicCell40 \ADC_VDC.i18807_4_lut_LC_12_6_6  (
            .in0(N__30601),
            .in1(N__32465),
            .in2(N__34768),
            .in3(N__30663),
            .lcout(\ADC_VDC.n21025 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i18117_2_lut_LC_12_6_7 .C_ON=1'b0;
    defparam \ADC_VDC.i18117_2_lut_LC_12_6_7 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i18117_2_lut_LC_12_6_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ADC_VDC.i18117_2_lut_LC_12_6_7  (
            .in0(_gnd_net_),
            .in1(N__34865),
            .in2(_gnd_net_),
            .in3(N__30636),
            .lcout(\ADC_VDC.n20712 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i19071_4_lut_4_lut_LC_12_7_0 .C_ON=1'b0;
    defparam \ADC_VDC.i19071_4_lut_4_lut_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i19071_4_lut_4_lut_LC_12_7_0 .LUT_INIT=16'b1111110011101101;
    LogicCell40 \ADC_VDC.i19071_4_lut_4_lut_LC_12_7_0  (
            .in0(N__34740),
            .in1(N__34368),
            .in2(N__34620),
            .in3(N__34157),
            .lcout(\ADC_VDC.n11662 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i18962_4_lut_LC_12_7_1 .C_ON=1'b0;
    defparam \ADC_VDC.i18962_4_lut_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i18962_4_lut_LC_12_7_1 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \ADC_VDC.i18962_4_lut_LC_12_7_1  (
            .in0(N__32590),
            .in1(N__32542),
            .in2(N__32640),
            .in3(N__32505),
            .lcout(\ADC_VDC.n21028 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_12_7_2.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_12_7_2.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_12_7_2.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_12_7_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_137_Mux_7_i1_3_lut_LC_12_7_3.C_ON=1'b0;
    defparam mux_137_Mux_7_i1_3_lut_LC_12_7_3.SEQ_MODE=4'b0000;
    defparam mux_137_Mux_7_i1_3_lut_LC_12_7_3.LUT_INIT=16'b1100110010101010;
    LogicCell40 mux_137_Mux_7_i1_3_lut_LC_12_7_3 (
            .in0(N__30810),
            .in1(N__42624),
            .in2(_gnd_net_),
            .in3(N__51632),
            .lcout(n1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i4_4_lut_adj_35_LC_12_7_4 .C_ON=1'b0;
    defparam \ADC_VDC.i4_4_lut_adj_35_LC_12_7_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i4_4_lut_adj_35_LC_12_7_4 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \ADC_VDC.i4_4_lut_adj_35_LC_12_7_4  (
            .in0(N__32541),
            .in1(N__32589),
            .in2(N__32511),
            .in3(N__32436),
            .lcout(\ADC_VDC.n10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i40_3_lut_4_lut_LC_12_7_6 .C_ON=1'b0;
    defparam \ADC_VDC.i40_3_lut_4_lut_LC_12_7_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i40_3_lut_4_lut_LC_12_7_6 .LUT_INIT=16'b1010110100100101;
    LogicCell40 \ADC_VDC.i40_3_lut_4_lut_LC_12_7_6  (
            .in0(N__34739),
            .in1(N__34156),
            .in2(N__34864),
            .in3(N__30771),
            .lcout(\ADC_VDC.n19_adj_1405 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam wdtick_cnt_3763_3764__i1_LC_12_8_0.C_ON=1'b0;
    defparam wdtick_cnt_3763_3764__i1_LC_12_8_0.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3763_3764__i1_LC_12_8_0.LUT_INIT=16'b0011001100010001;
    LogicCell40 wdtick_cnt_3763_3764__i1_LC_12_8_0 (
            .in0(N__30701),
            .in1(N__30740),
            .in2(_gnd_net_),
            .in3(N__30721),
            .lcout(wdtick_cnt_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40928),
            .ce(N__33040),
            .sr(N__40683));
    defparam wdtick_cnt_3763_3764__i3_LC_12_8_1.C_ON=1'b0;
    defparam wdtick_cnt_3763_3764__i3_LC_12_8_1.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3763_3764__i3_LC_12_8_1.LUT_INIT=16'b0101101010100000;
    LogicCell40 wdtick_cnt_3763_3764__i3_LC_12_8_1 (
            .in0(N__30723),
            .in1(_gnd_net_),
            .in2(N__30745),
            .in3(N__30702),
            .lcout(wdtick_cnt_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40928),
            .ce(N__33040),
            .sr(N__40683));
    defparam wdtick_cnt_3763_3764__i2_LC_12_8_2.C_ON=1'b0;
    defparam wdtick_cnt_3763_3764__i2_LC_12_8_2.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3763_3764__i2_LC_12_8_2.LUT_INIT=16'b0011001111001100;
    LogicCell40 wdtick_cnt_3763_3764__i2_LC_12_8_2 (
            .in0(_gnd_net_),
            .in1(N__30739),
            .in2(_gnd_net_),
            .in3(N__30722),
            .lcout(wdtick_cnt_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40928),
            .ce(N__33040),
            .sr(N__40683));
    defparam wdtick_flag_289_LC_12_9_0.C_ON=1'b0;
    defparam wdtick_flag_289_LC_12_9_0.SEQ_MODE=4'b1010;
    defparam wdtick_flag_289_LC_12_9_0.LUT_INIT=16'b1111111100010000;
    LogicCell40 wdtick_flag_289_LC_12_9_0 (
            .in0(N__30744),
            .in1(N__30724),
            .in2(N__30706),
            .in3(N__50256),
            .lcout(wdtick_flag),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40938),
            .ce(),
            .sr(N__40684));
    defparam i1_2_lut_LC_12_10_0.C_ON=1'b0;
    defparam i1_2_lut_LC_12_10_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_LC_12_10_0.LUT_INIT=16'b1111111110101010;
    LogicCell40 i1_2_lut_LC_12_10_0 (
            .in0(N__51209),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54563),
            .lcout(n12205),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18699_2_lut_LC_12_10_1.C_ON=1'b0;
    defparam i18699_2_lut_LC_12_10_1.SEQ_MODE=4'b0000;
    defparam i18699_2_lut_LC_12_10_1.LUT_INIT=16'b1111111110101010;
    LogicCell40 i18699_2_lut_LC_12_10_1 (
            .in0(N__38202),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53462),
            .lcout(n20931),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i7_LC_12_10_2.C_ON=1'b0;
    defparam comm_cmd_i7_LC_12_10_2.SEQ_MODE=4'b1000;
    defparam comm_cmd_i7_LC_12_10_2.LUT_INIT=16'b1101010110000000;
    LogicCell40 comm_cmd_i7_LC_12_10_2 (
            .in0(N__30932),
            .in1(N__30992),
            .in2(N__36897),
            .in3(N__49288),
            .lcout(comm_cmd_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55081),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i3_LC_12_10_3.C_ON=1'b0;
    defparam comm_cmd_i3_LC_12_10_3.SEQ_MODE=4'b1000;
    defparam comm_cmd_i3_LC_12_10_3.LUT_INIT=16'b1100000010101010;
    LogicCell40 comm_cmd_i3_LC_12_10_3 (
            .in0(N__56146),
            .in1(N__30991),
            .in2(N__35567),
            .in3(N__30931),
            .lcout(comm_cmd_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55081),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_278_LC_12_10_4.C_ON=1'b0;
    defparam i1_3_lut_adj_278_LC_12_10_4.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_278_LC_12_10_4.LUT_INIT=16'b1111111111101110;
    LogicCell40 i1_3_lut_adj_278_LC_12_10_4 (
            .in0(N__53461),
            .in1(N__56144),
            .in2(_gnd_net_),
            .in3(N__38201),
            .lcout(n20622),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_0_i30_3_lut_LC_12_10_6.C_ON=1'b0;
    defparam mux_130_Mux_0_i30_3_lut_LC_12_10_6.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_0_i30_3_lut_LC_12_10_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_130_Mux_0_i30_3_lut_LC_12_10_6 (
            .in0(N__30898),
            .in1(N__30883),
            .in2(_gnd_net_),
            .in3(N__56145),
            .lcout(n30_adj_1475),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_120_LC_12_10_7.C_ON=1'b0;
    defparam i1_2_lut_adj_120_LC_12_10_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_120_LC_12_10_7.LUT_INIT=16'b1010101011111111;
    LogicCell40 i1_2_lut_adj_120_LC_12_10_7 (
            .in0(N__54562),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51208),
            .lcout(n20627),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_4__i0_LC_12_11_0.C_ON=1'b0;
    defparam comm_buf_4__i0_LC_12_11_0.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i0_LC_12_11_0.LUT_INIT=16'b1110111000100010;
    LogicCell40 comm_buf_4__i0_LC_12_11_0 (
            .in0(N__30871),
            .in1(N__53979),
            .in2(_gnd_net_),
            .in3(N__36252),
            .lcout(comm_buf_4_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55086),
            .ce(N__49825),
            .sr(N__33106));
    defparam comm_buf_4__i7_LC_12_11_1.C_ON=1'b0;
    defparam comm_buf_4__i7_LC_12_11_1.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i7_LC_12_11_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_4__i7_LC_12_11_1 (
            .in0(N__53978),
            .in1(N__36881),
            .in2(_gnd_net_),
            .in3(N__30850),
            .lcout(comm_buf_4_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55086),
            .ce(N__49825),
            .sr(N__33106));
    defparam comm_buf_4__i6_LC_12_11_2.C_ON=1'b0;
    defparam comm_buf_4__i6_LC_12_11_2.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i6_LC_12_11_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_4__i6_LC_12_11_2 (
            .in0(N__35802),
            .in1(N__30832),
            .in2(_gnd_net_),
            .in3(N__53982),
            .lcout(comm_buf_4_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55086),
            .ce(N__49825),
            .sr(N__33106));
    defparam comm_buf_4__i5_LC_12_11_3.C_ON=1'b0;
    defparam comm_buf_4__i5_LC_12_11_3.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i5_LC_12_11_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_4__i5_LC_12_11_3 (
            .in0(N__53977),
            .in1(N__38017),
            .in2(_gnd_net_),
            .in3(N__31123),
            .lcout(comm_buf_4_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55086),
            .ce(N__49825),
            .sr(N__33106));
    defparam comm_buf_4__i4_LC_12_11_4.C_ON=1'b0;
    defparam comm_buf_4__i4_LC_12_11_4.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i4_LC_12_11_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_4__i4_LC_12_11_4 (
            .in0(N__35664),
            .in1(N__31105),
            .in2(_gnd_net_),
            .in3(N__53981),
            .lcout(comm_buf_4_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55086),
            .ce(N__49825),
            .sr(N__33106));
    defparam comm_buf_4__i3_LC_12_11_5.C_ON=1'b0;
    defparam comm_buf_4__i3_LC_12_11_5.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i3_LC_12_11_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_4__i3_LC_12_11_5 (
            .in0(N__53976),
            .in1(N__35559),
            .in2(_gnd_net_),
            .in3(N__31087),
            .lcout(comm_buf_4_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55086),
            .ce(N__49825),
            .sr(N__33106));
    defparam comm_buf_4__i2_LC_12_11_6.C_ON=1'b0;
    defparam comm_buf_4__i2_LC_12_11_6.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i2_LC_12_11_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_4__i2_LC_12_11_6 (
            .in0(N__35451),
            .in1(N__31069),
            .in2(_gnd_net_),
            .in3(N__53980),
            .lcout(comm_buf_4_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55086),
            .ce(N__49825),
            .sr(N__33106));
    defparam comm_buf_4__i1_LC_12_11_7.C_ON=1'b0;
    defparam comm_buf_4__i1_LC_12_11_7.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i1_LC_12_11_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_4__i1_LC_12_11_7 (
            .in0(N__53975),
            .in1(N__35967),
            .in2(_gnd_net_),
            .in3(N__31048),
            .lcout(comm_buf_4_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55086),
            .ce(N__49825),
            .sr(N__33106));
    defparam data_idxvec_i0_LC_12_12_0.C_ON=1'b1;
    defparam data_idxvec_i0_LC_12_12_0.SEQ_MODE=4'b1000;
    defparam data_idxvec_i0_LC_12_12_0.LUT_INIT=16'b1010001110101100;
    LogicCell40 data_idxvec_i0_LC_12_12_0 (
            .in0(N__31027),
            .in1(N__35895),
            .in2(N__54711),
            .in3(N__31012),
            .lcout(data_idxvec_0),
            .ltout(),
            .carryin(bfn_12_12_0_),
            .carryout(n19335),
            .clk(N__55094),
            .ce(N__38581),
            .sr(_gnd_net_));
    defparam data_idxvec_i1_LC_12_12_1.C_ON=1'b1;
    defparam data_idxvec_i1_LC_12_12_1.SEQ_MODE=4'b1000;
    defparam data_idxvec_i1_LC_12_12_1.LUT_INIT=16'b1010001110101100;
    LogicCell40 data_idxvec_i1_LC_12_12_1 (
            .in0(N__38443),
            .in1(N__36039),
            .in2(N__54713),
            .in3(N__31009),
            .lcout(data_idxvec_1),
            .ltout(),
            .carryin(n19335),
            .carryout(n19336),
            .clk(N__55094),
            .ce(N__38581),
            .sr(_gnd_net_));
    defparam data_idxvec_i2_LC_12_12_2.C_ON=1'b1;
    defparam data_idxvec_i2_LC_12_12_2.SEQ_MODE=4'b1000;
    defparam data_idxvec_i2_LC_12_12_2.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i2_LC_12_12_2 (
            .in0(N__41283),
            .in1(N__54645),
            .in2(N__33340),
            .in3(N__31006),
            .lcout(data_idxvec_2),
            .ltout(),
            .carryin(n19336),
            .carryout(n19337),
            .clk(N__55094),
            .ce(N__38581),
            .sr(_gnd_net_));
    defparam data_idxvec_i3_LC_12_12_3.C_ON=1'b1;
    defparam data_idxvec_i3_LC_12_12_3.SEQ_MODE=4'b1000;
    defparam data_idxvec_i3_LC_12_12_3.LUT_INIT=16'b1010001110101100;
    LogicCell40 data_idxvec_i3_LC_12_12_3 (
            .in0(N__38855),
            .in1(N__33390),
            .in2(N__54714),
            .in3(N__31003),
            .lcout(data_idxvec_3),
            .ltout(),
            .carryin(n19337),
            .carryout(n19338),
            .clk(N__55094),
            .ce(N__38581),
            .sr(_gnd_net_));
    defparam data_idxvec_i4_LC_12_12_4.C_ON=1'b1;
    defparam data_idxvec_i4_LC_12_12_4.SEQ_MODE=4'b1000;
    defparam data_idxvec_i4_LC_12_12_4.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i4_LC_12_12_4 (
            .in0(N__38470),
            .in1(N__54649),
            .in2(N__33439),
            .in3(N__31228),
            .lcout(data_idxvec_4),
            .ltout(),
            .carryin(n19338),
            .carryout(n19339),
            .clk(N__55094),
            .ce(N__38581),
            .sr(_gnd_net_));
    defparam data_idxvec_i5_LC_12_12_5.C_ON=1'b1;
    defparam data_idxvec_i5_LC_12_12_5.SEQ_MODE=4'b1000;
    defparam data_idxvec_i5_LC_12_12_5.LUT_INIT=16'b1010001110101100;
    LogicCell40 data_idxvec_i5_LC_12_12_5 (
            .in0(N__50132),
            .in1(N__31287),
            .in2(N__54715),
            .in3(N__31225),
            .lcout(data_idxvec_5),
            .ltout(),
            .carryin(n19339),
            .carryout(n19340),
            .clk(N__55094),
            .ce(N__38581),
            .sr(_gnd_net_));
    defparam data_idxvec_i6_LC_12_12_6.C_ON=1'b1;
    defparam data_idxvec_i6_LC_12_12_6.SEQ_MODE=4'b1000;
    defparam data_idxvec_i6_LC_12_12_6.LUT_INIT=16'b1010001110101100;
    LogicCell40 data_idxvec_i6_LC_12_12_6 (
            .in0(N__51375),
            .in1(N__31221),
            .in2(N__54712),
            .in3(N__31207),
            .lcout(data_idxvec_6),
            .ltout(),
            .carryin(n19340),
            .carryout(n19341),
            .clk(N__55094),
            .ce(N__38581),
            .sr(_gnd_net_));
    defparam data_idxvec_i7_LC_12_12_7.C_ON=1'b1;
    defparam data_idxvec_i7_LC_12_12_7.SEQ_MODE=4'b1000;
    defparam data_idxvec_i7_LC_12_12_7.LUT_INIT=16'b1010001110101100;
    LogicCell40 data_idxvec_i7_LC_12_12_7 (
            .in0(N__41259),
            .in1(N__36678),
            .in2(N__54716),
            .in3(N__31204),
            .lcout(data_idxvec_7),
            .ltout(),
            .carryin(n19341),
            .carryout(n19342),
            .clk(N__55094),
            .ce(N__38581),
            .sr(_gnd_net_));
    defparam data_idxvec_i8_LC_12_13_0.C_ON=1'b1;
    defparam data_idxvec_i8_LC_12_13_0.SEQ_MODE=4'b1000;
    defparam data_idxvec_i8_LC_12_13_0.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i8_LC_12_13_0 (
            .in0(N__41781),
            .in1(N__54576),
            .in2(N__41470),
            .in3(N__31201),
            .lcout(data_idxvec_8),
            .ltout(),
            .carryin(bfn_12_13_0_),
            .carryout(n19343),
            .clk(N__55103),
            .ce(N__38580),
            .sr(_gnd_net_));
    defparam data_idxvec_i9_LC_12_13_1.C_ON=1'b1;
    defparam data_idxvec_i9_LC_12_13_1.SEQ_MODE=4'b1000;
    defparam data_idxvec_i9_LC_12_13_1.LUT_INIT=16'b1010001110101100;
    LogicCell40 data_idxvec_i9_LC_12_13_1 (
            .in0(N__38143),
            .in1(N__31194),
            .in2(N__54693),
            .in3(N__31180),
            .lcout(data_idxvec_9),
            .ltout(),
            .carryin(n19343),
            .carryout(n19344),
            .clk(N__55103),
            .ce(N__38580),
            .sr(_gnd_net_));
    defparam data_idxvec_i10_LC_12_13_2.C_ON=1'b1;
    defparam data_idxvec_i10_LC_12_13_2.SEQ_MODE=4'b1000;
    defparam data_idxvec_i10_LC_12_13_2.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i10_LC_12_13_2 (
            .in0(N__41943),
            .in1(N__54580),
            .in2(N__31177),
            .in3(N__31156),
            .lcout(data_idxvec_10),
            .ltout(),
            .carryin(n19344),
            .carryout(n19345),
            .clk(N__55103),
            .ce(N__38580),
            .sr(_gnd_net_));
    defparam data_idxvec_i11_LC_12_13_3.C_ON=1'b1;
    defparam data_idxvec_i11_LC_12_13_3.SEQ_MODE=4'b1000;
    defparam data_idxvec_i11_LC_12_13_3.LUT_INIT=16'b1010001110101100;
    LogicCell40 data_idxvec_i11_LC_12_13_3 (
            .in0(N__38590),
            .in1(N__44988),
            .in2(N__54694),
            .in3(N__31153),
            .lcout(data_idxvec_11),
            .ltout(),
            .carryin(n19345),
            .carryout(n19346),
            .clk(N__55103),
            .ce(N__38580),
            .sr(_gnd_net_));
    defparam data_idxvec_i12_LC_12_13_4.C_ON=1'b1;
    defparam data_idxvec_i12_LC_12_13_4.SEQ_MODE=4'b1000;
    defparam data_idxvec_i12_LC_12_13_4.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i12_LC_12_13_4 (
            .in0(N__42126),
            .in1(N__54584),
            .in2(N__31146),
            .in3(N__31126),
            .lcout(data_idxvec_12),
            .ltout(),
            .carryin(n19346),
            .carryout(n19347),
            .clk(N__55103),
            .ce(N__38580),
            .sr(_gnd_net_));
    defparam data_idxvec_i13_LC_12_13_5.C_ON=1'b1;
    defparam data_idxvec_i13_LC_12_13_5.SEQ_MODE=4'b1000;
    defparam data_idxvec_i13_LC_12_13_5.LUT_INIT=16'b1010001110101100;
    LogicCell40 data_idxvec_i13_LC_12_13_5 (
            .in0(N__44849),
            .in1(N__31356),
            .in2(N__54695),
            .in3(N__31342),
            .lcout(data_idxvec_13),
            .ltout(),
            .carryin(n19347),
            .carryout(n19348),
            .clk(N__55103),
            .ce(N__38580),
            .sr(_gnd_net_));
    defparam data_idxvec_i14_LC_12_13_6.C_ON=1'b1;
    defparam data_idxvec_i14_LC_12_13_6.SEQ_MODE=4'b1000;
    defparam data_idxvec_i14_LC_12_13_6.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i14_LC_12_13_6 (
            .in0(N__41526),
            .in1(N__54588),
            .in2(N__31332),
            .in3(N__31312),
            .lcout(data_idxvec_14),
            .ltout(),
            .carryin(n19348),
            .carryout(n19349),
            .clk(N__55103),
            .ce(N__38580),
            .sr(_gnd_net_));
    defparam data_idxvec_i15_LC_12_13_7.C_ON=1'b0;
    defparam data_idxvec_i15_LC_12_13_7.SEQ_MODE=4'b1000;
    defparam data_idxvec_i15_LC_12_13_7.LUT_INIT=16'b1011000111100100;
    LogicCell40 data_idxvec_i15_LC_12_13_7 (
            .in0(N__54589),
            .in1(N__31302),
            .in2(N__45772),
            .in3(N__31309),
            .lcout(data_idxvec_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55103),
            .ce(N__38580),
            .sr(_gnd_net_));
    defparam mux_129_Mux_5_i26_3_lut_LC_12_14_2.C_ON=1'b0;
    defparam mux_129_Mux_5_i26_3_lut_LC_12_14_2.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_5_i26_3_lut_LC_12_14_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_129_Mux_5_i26_3_lut_LC_12_14_2 (
            .in0(N__56890),
            .in1(N__31288),
            .in2(_gnd_net_),
            .in3(N__46783),
            .lcout(),
            .ltout(n26_adj_1486_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19546_LC_12_14_3.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19546_LC_12_14_3.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19546_LC_12_14_3.LUT_INIT=16'b1101100010101010;
    LogicCell40 comm_cmd_1__bdd_4_lut_19546_LC_12_14_3 (
            .in0(N__57523),
            .in1(N__31234),
            .in2(N__31273),
            .in3(N__47786),
            .lcout(),
            .ltout(n22177_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22177_bdd_4_lut_LC_12_14_4.C_ON=1'b0;
    defparam n22177_bdd_4_lut_LC_12_14_4.SEQ_MODE=4'b0000;
    defparam n22177_bdd_4_lut_LC_12_14_4.LUT_INIT=16'b1110010111100000;
    LogicCell40 n22177_bdd_4_lut_LC_12_14_4 (
            .in0(N__47787),
            .in1(N__38422),
            .in2(N__31270),
            .in3(N__31376),
            .lcout(),
            .ltout(n22180_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1542877_i1_3_lut_LC_12_14_5.C_ON=1'b0;
    defparam i1542877_i1_3_lut_LC_12_14_5.SEQ_MODE=4'b0000;
    defparam i1542877_i1_3_lut_LC_12_14_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 i1542877_i1_3_lut_LC_12_14_5 (
            .in0(_gnd_net_),
            .in1(N__31267),
            .in2(N__31255),
            .in3(N__56257),
            .lcout(),
            .ltout(n30_adj_1485_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i5_LC_12_14_6.C_ON=1'b0;
    defparam comm_buf_1__i5_LC_12_14_6.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i5_LC_12_14_6.LUT_INIT=16'b1101100011011000;
    LogicCell40 comm_buf_1__i5_LC_12_14_6 (
            .in0(N__54095),
            .in1(N__38018),
            .in2(N__31252),
            .in3(_gnd_net_),
            .lcout(comm_buf_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55112),
            .ce(N__38546),
            .sr(N__36808));
    defparam i18810_2_lut_LC_12_14_7.C_ON=1'b0;
    defparam i18810_2_lut_LC_12_14_7.SEQ_MODE=4'b0000;
    defparam i18810_2_lut_LC_12_14_7.LUT_INIT=16'b1111111111001100;
    LogicCell40 i18810_2_lut_LC_12_14_7 (
            .in0(_gnd_net_),
            .in1(N__31249),
            .in2(_gnd_net_),
            .in3(N__56889),
            .lcout(n21036),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i3_LC_12_15_0.C_ON=1'b0;
    defparam data_index_i3_LC_12_15_0.SEQ_MODE=4'b1000;
    defparam data_index_i3_LC_12_15_0.LUT_INIT=16'b0010111000100010;
    LogicCell40 data_index_i3_LC_12_15_0 (
            .in0(N__41797),
            .in1(N__54591),
            .in2(N__52194),
            .in3(N__36346),
            .lcout(data_index_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55123),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_354_Mux_0_i15_4_lut_LC_12_15_1.C_ON=1'b0;
    defparam comm_state_3__I_0_354_Mux_0_i15_4_lut_LC_12_15_1.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_354_Mux_0_i15_4_lut_LC_12_15_1.LUT_INIT=16'b0100111001000100;
    LogicCell40 comm_state_3__I_0_354_Mux_0_i15_4_lut_LC_12_15_1 (
            .in0(N__54590),
            .in1(N__42874),
            .in2(N__52091),
            .in3(N__42859),
            .lcout(data_index_9_N_212_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4_4_lut_adj_316_LC_12_15_2.C_ON=1'b0;
    defparam i4_4_lut_adj_316_LC_12_15_2.SEQ_MODE=4'b0000;
    defparam i4_4_lut_adj_316_LC_12_15_2.LUT_INIT=16'b0111101111011110;
    LogicCell40 i4_4_lut_adj_316_LC_12_15_2 (
            .in0(N__33610),
            .in1(N__33655),
            .in2(N__31381),
            .in3(N__33353),
            .lcout(),
            .ltout(n20_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10_4_lut_LC_12_15_3.C_ON=1'b0;
    defparam i10_4_lut_LC_12_15_3.SEQ_MODE=4'b0000;
    defparam i10_4_lut_LC_12_15_3.LUT_INIT=16'b1111111111110110;
    LogicCell40 i10_4_lut_LC_12_15_3 (
            .in0(N__33733),
            .in1(N__31529),
            .in2(N__31513),
            .in3(N__31510),
            .lcout(),
            .ltout(n26_adj_1604_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15_4_lut_LC_12_15_4.C_ON=1'b0;
    defparam i15_4_lut_LC_12_15_4.SEQ_MODE=4'b0000;
    defparam i15_4_lut_LC_12_15_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i15_4_lut_LC_12_15_4 (
            .in0(N__31501),
            .in1(N__31891),
            .in2(N__31492),
            .in3(N__36271),
            .lcout(n31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_354_Mux_3_i15_4_lut_LC_12_15_5.C_ON=1'b0;
    defparam comm_state_3__I_0_354_Mux_3_i15_4_lut_LC_12_15_5.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_354_Mux_3_i15_4_lut_LC_12_15_5.LUT_INIT=16'b0011101100001000;
    LogicCell40 comm_state_3__I_0_354_Mux_3_i15_4_lut_LC_12_15_5 (
            .in0(N__36345),
            .in1(N__54592),
            .in2(N__52092),
            .in3(N__41796),
            .lcout(data_index_9_N_212_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i3_LC_12_15_6.C_ON=1'b0;
    defparam acadc_skipCount_i3_LC_12_15_6.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i3_LC_12_15_6.LUT_INIT=16'b0111001101000000;
    LogicCell40 acadc_skipCount_i3_LC_12_15_6 (
            .in0(N__52181),
            .in1(N__39323),
            .in2(N__36396),
            .in3(N__33354),
            .lcout(acadc_skipCount_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55123),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i5_LC_12_15_7.C_ON=1'b0;
    defparam acadc_skipCount_i5_LC_12_15_7.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i5_LC_12_15_7.LUT_INIT=16'b0000101011001010;
    LogicCell40 acadc_skipCount_i5_LC_12_15_7 (
            .in0(N__31377),
            .in1(N__50181),
            .in2(N__39331),
            .in3(N__52185),
            .lcout(acadc_skipCount_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55123),
            .ce(),
            .sr(_gnd_net_));
    defparam i19091_2_lut_LC_12_16_0.C_ON=1'b0;
    defparam i19091_2_lut_LC_12_16_0.SEQ_MODE=4'b0000;
    defparam i19091_2_lut_LC_12_16_0.LUT_INIT=16'b0000101000001010;
    LogicCell40 i19091_2_lut_LC_12_16_0 (
            .in0(N__33914),
            .in1(_gnd_net_),
            .in2(N__32185),
            .in3(_gnd_net_),
            .lcout(n14639),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_2_i16_3_lut_LC_12_16_1.C_ON=1'b0;
    defparam mux_129_Mux_2_i16_3_lut_LC_12_16_1.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_2_i16_3_lut_LC_12_16_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_129_Mux_2_i16_3_lut_LC_12_16_1 (
            .in0(N__32012),
            .in1(N__42753),
            .in2(_gnd_net_),
            .in3(N__56897),
            .lcout(n16_adj_1504),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i1_LC_12_16_2.C_ON=1'b0;
    defparam buf_dds1_i1_LC_12_16_2.SEQ_MODE=4'b1000;
    defparam buf_dds1_i1_LC_12_16_2.LUT_INIT=16'b1101100000000000;
    LogicCell40 buf_dds1_i1_LC_12_16_2 (
            .in0(N__45839),
            .in1(N__43382),
            .in2(N__31931),
            .in3(N__46013),
            .lcout(buf_dds1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55133),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_53_LC_12_16_3.C_ON=1'b0;
    defparam i1_4_lut_adj_53_LC_12_16_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_53_LC_12_16_3.LUT_INIT=16'b0111110110111110;
    LogicCell40 i1_4_lut_adj_53_LC_12_16_3 (
            .in0(N__33492),
            .in1(N__31904),
            .in2(N__33754),
            .in3(N__35855),
            .lcout(n17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i1_2_lut_LC_12_16_4 .C_ON=1'b0;
    defparam \ADC_VAC.i1_2_lut_LC_12_16_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i1_2_lut_LC_12_16_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ADC_VAC.i1_2_lut_LC_12_16_4  (
            .in0(_gnd_net_),
            .in1(N__31883),
            .in2(_gnd_net_),
            .in3(N__31860),
            .lcout(iac_raw_buf_N_728),
            .ltout(iac_raw_buf_N_728_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_state_1__bdd_4_lut_4_lut_LC_12_16_5.C_ON=1'b0;
    defparam eis_state_1__bdd_4_lut_4_lut_LC_12_16_5.SEQ_MODE=4'b0000;
    defparam eis_state_1__bdd_4_lut_4_lut_LC_12_16_5.LUT_INIT=16'b1000111010101010;
    LogicCell40 eis_state_1__bdd_4_lut_4_lut_LC_12_16_5 (
            .in0(N__39137),
            .in1(N__32181),
            .in2(N__31840),
            .in3(N__37604),
            .lcout(n21997),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i3_LC_12_16_6.C_ON=1'b0;
    defparam buf_dds1_i3_LC_12_16_6.SEQ_MODE=4'b1000;
    defparam buf_dds1_i3_LC_12_16_6.LUT_INIT=16'b1110010011101110;
    LogicCell40 buf_dds1_i3_LC_12_16_6 (
            .in0(N__45838),
            .in1(N__31820),
            .in2(N__38869),
            .in3(N__54710),
            .lcout(buf_dds1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55133),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_274_LC_12_17_1.C_ON=1'b0;
    defparam i1_3_lut_adj_274_LC_12_17_1.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_274_LC_12_17_1.LUT_INIT=16'b1101110100000000;
    LogicCell40 i1_3_lut_adj_274_LC_12_17_1 (
            .in0(N__31804),
            .in1(N__52173),
            .in2(_gnd_net_),
            .in3(N__54596),
            .lcout(n12353),
            .ltout(n12353_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i1_LC_12_17_2.C_ON=1'b0;
    defparam buf_dds0_i1_LC_12_17_2.SEQ_MODE=4'b1000;
    defparam buf_dds0_i1_LC_12_17_2.LUT_INIT=16'b0100111101000000;
    LogicCell40 buf_dds0_i1_LC_12_17_2 (
            .in0(N__52175),
            .in1(N__43390),
            .in2(N__31792),
            .in3(N__32231),
            .lcout(buf_dds0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55145),
            .ce(),
            .sr(_gnd_net_));
    defparam i3787_3_lut_4_lut_4_lut_LC_12_17_3.C_ON=1'b0;
    defparam i3787_3_lut_4_lut_4_lut_LC_12_17_3.SEQ_MODE=4'b0000;
    defparam i3787_3_lut_4_lut_4_lut_LC_12_17_3.LUT_INIT=16'b0001000000000000;
    LogicCell40 i3787_3_lut_4_lut_4_lut_LC_12_17_3 (
            .in0(N__32070),
            .in1(N__32179),
            .in2(N__31789),
            .in3(N__46968),
            .lcout(iac_raw_buf_N_726),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19122_4_lut_LC_12_17_4.C_ON=1'b0;
    defparam i19122_4_lut_LC_12_17_4.SEQ_MODE=4'b0000;
    defparam i19122_4_lut_LC_12_17_4.LUT_INIT=16'b0000000000000111;
    LogicCell40 i19122_4_lut_LC_12_17_4 (
            .in0(N__32178),
            .in1(N__37602),
            .in2(N__32087),
            .in3(N__39142),
            .lcout(n11538),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18710_2_lut_LC_12_17_5.C_ON=1'b0;
    defparam i18710_2_lut_LC_12_17_5.SEQ_MODE=4'b0000;
    defparam i18710_2_lut_LC_12_17_5.LUT_INIT=16'b0101010100000000;
    LogicCell40 i18710_2_lut_LC_12_17_5 (
            .in0(N__56888),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32032),
            .lcout(n20949),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i0_LC_12_17_6.C_ON=1'b0;
    defparam buf_dds0_i0_LC_12_17_6.SEQ_MODE=4'b1000;
    defparam buf_dds0_i0_LC_12_17_6.LUT_INIT=16'b0100010011110000;
    LogicCell40 buf_dds0_i0_LC_12_17_6 (
            .in0(N__52174),
            .in1(N__41355),
            .in2(N__40373),
            .in3(N__45655),
            .lcout(buf_dds0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55145),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i2_LC_12_17_7.C_ON=1'b0;
    defparam buf_dds1_i2_LC_12_17_7.SEQ_MODE=4'b1000;
    defparam buf_dds1_i2_LC_12_17_7.LUT_INIT=16'b1010000010001000;
    LogicCell40 buf_dds1_i2_LC_12_17_7 (
            .in0(N__46014),
            .in1(N__32016),
            .in2(N__42823),
            .in3(N__45895),
            .lcout(buf_dds1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55145),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i7_LC_12_18_0 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i7_LC_12_18_0 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i7_LC_12_18_0 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \SIG_DDS.tmp_buf_i7_LC_12_18_0  (
            .in0(N__39064),
            .in1(N__37138),
            .in2(N__55888),
            .in3(N__55622),
            .lcout(\SIG_DDS.tmp_buf_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55160),
            .ce(N__40330),
            .sr(_gnd_net_));
    defparam \SIG_DDS.i12468_3_lut_LC_12_18_1 .C_ON=1'b0;
    defparam \SIG_DDS.i12468_3_lut_LC_12_18_1 .SEQ_MODE=4'b0000;
    defparam \SIG_DDS.i12468_3_lut_LC_12_18_1 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \SIG_DDS.i12468_3_lut_LC_12_18_1  (
            .in0(N__55711),
            .in1(N__55873),
            .in2(_gnd_net_),
            .in3(N__55620),
            .lcout(n14869),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.i19105_4_lut_LC_12_18_3 .C_ON=1'b0;
    defparam \SIG_DDS.i19105_4_lut_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \SIG_DDS.i19105_4_lut_LC_12_18_3 .LUT_INIT=16'b1111111111011110;
    LogicCell40 \SIG_DDS.i19105_4_lut_LC_12_18_3  (
            .in0(N__55712),
            .in1(N__55874),
            .in2(N__53018),
            .in3(N__55621),
            .lcout(\SIG_DDS.n9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_7_i16_3_lut_LC_12_18_5.C_ON=1'b0;
    defparam mux_129_Mux_7_i16_3_lut_LC_12_18_5.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_7_i16_3_lut_LC_12_18_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_129_Mux_7_i16_3_lut_LC_12_18_5 (
            .in0(N__42543),
            .in1(N__39063),
            .in2(_gnd_net_),
            .in3(N__56964),
            .lcout(),
            .ltout(n16_adj_1621_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n21961_bdd_4_lut_LC_12_18_6.C_ON=1'b0;
    defparam n21961_bdd_4_lut_LC_12_18_6.SEQ_MODE=4'b0000;
    defparam n21961_bdd_4_lut_LC_12_18_6.LUT_INIT=16'b1100110010111000;
    LogicCell40 n21961_bdd_4_lut_LC_12_18_6 (
            .in0(N__31986),
            .in1(N__31960),
            .in2(N__31948),
            .in3(N__47834),
            .lcout(n21964),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i10_LC_12_19_0 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i10_LC_12_19_0 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i10_LC_12_19_0 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \SIG_DDS.tmp_buf_i10_LC_12_19_0  (
            .in0(N__55880),
            .in1(N__32371),
            .in2(N__32320),
            .in3(N__55662),
            .lcout(\SIG_DDS.tmp_buf_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55175),
            .ce(N__40329),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i11_LC_12_19_1 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i11_LC_12_19_1 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i11_LC_12_19_1 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \SIG_DDS.tmp_buf_i11_LC_12_19_1  (
            .in0(N__55663),
            .in1(N__55881),
            .in2(N__43108),
            .in3(N__32350),
            .lcout(\SIG_DDS.tmp_buf_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55175),
            .ce(N__40329),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i9_LC_12_19_2 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i9_LC_12_19_2 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i9_LC_12_19_2 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \SIG_DDS.tmp_buf_i9_LC_12_19_2  (
            .in0(N__55886),
            .in1(N__55668),
            .in2(N__32203),
            .in3(N__32344),
            .lcout(\SIG_DDS.tmp_buf_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55175),
            .ce(N__40329),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i13_LC_12_19_3 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i13_LC_12_19_3 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i13_LC_12_19_3 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \SIG_DDS.tmp_buf_i13_LC_12_19_3  (
            .in0(N__55664),
            .in1(N__55882),
            .in2(N__33838),
            .in3(N__32311),
            .lcout(\SIG_DDS.tmp_buf_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55175),
            .ce(N__40329),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i14_LC_12_19_4 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i14_LC_12_19_4 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i14_LC_12_19_4 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \SIG_DDS.tmp_buf_i14_LC_12_19_4  (
            .in0(N__55883),
            .in1(N__55665),
            .in2(N__32281),
            .in3(N__32271),
            .lcout(\SIG_DDS.tmp_buf_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55175),
            .ce(N__40329),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i1_LC_12_19_5 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i1_LC_12_19_5 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i1_LC_12_19_5 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \SIG_DDS.tmp_buf_i1_LC_12_19_5  (
            .in0(N__55666),
            .in1(N__55884),
            .in2(N__40342),
            .in3(N__32238),
            .lcout(\SIG_DDS.tmp_buf_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55175),
            .ce(N__40329),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i8_LC_12_19_7 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i8_LC_12_19_7 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i8_LC_12_19_7 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \SIG_DDS.tmp_buf_i8_LC_12_19_7  (
            .in0(N__55667),
            .in1(N__55885),
            .in2(N__32212),
            .in3(N__43417),
            .lcout(\SIG_DDS.tmp_buf_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55175),
            .ce(N__40329),
            .sr(_gnd_net_));
    defparam \comm_spi.i19174_4_lut_3_lut_LC_13_3_0 .C_ON=1'b0;
    defparam \comm_spi.i19174_4_lut_3_lut_LC_13_3_0 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19174_4_lut_3_lut_LC_13_3_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \comm_spi.i19174_4_lut_3_lut_LC_13_3_0  (
            .in0(N__32194),
            .in1(N__32409),
            .in2(_gnd_net_),
            .in3(N__55464),
            .lcout(\comm_spi.n22629 ),
            .ltout(\comm_spi.n22629_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i12199_3_lut_LC_13_3_1 .C_ON=1'b0;
    defparam \comm_spi.i12199_3_lut_LC_13_3_1 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i12199_3_lut_LC_13_3_1 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \comm_spi.i12199_3_lut_LC_13_3_1  (
            .in0(N__32401),
            .in1(_gnd_net_),
            .in2(N__32188),
            .in3(N__33802),
            .lcout(comm_rx_buf_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.t_clk_24_LC_13_3_2 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.t_clk_24_LC_13_3_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t_clk_24_LC_13_3_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ADC_VDC.genclk.t_clk_24_LC_13_3_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34931),
            .lcout(VDC_CLK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVADC_VDC.genclk.t_clk_24C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.div_state_i0_LC_13_3_3 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.div_state_i0_LC_13_3_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.div_state_i0_LC_13_3_3 .LUT_INIT=16'b1011111110110011;
    LogicCell40 \ADC_VDC.genclk.div_state_i0_LC_13_3_3  (
            .in0(N__32383),
            .in1(N__34970),
            .in2(N__34936),
            .in3(N__33781),
            .lcout(\ADC_VDC.genclk.div_state_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVADC_VDC.genclk.t_clk_24C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i19159_4_lut_3_lut_LC_13_3_4 .C_ON=1'b0;
    defparam \comm_spi.i19159_4_lut_3_lut_LC_13_3_4 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19159_4_lut_3_lut_LC_13_3_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.i19159_4_lut_3_lut_LC_13_3_4  (
            .in0(N__37346),
            .in1(N__33818),
            .in2(_gnd_net_),
            .in3(N__55463),
            .lcout(\comm_spi.n22632 ),
            .ltout(\comm_spi.n22632_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i12185_3_lut_LC_13_3_5 .C_ON=1'b0;
    defparam \comm_spi.i12185_3_lut_LC_13_3_5 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i12185_3_lut_LC_13_3_5 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \comm_spi.i12185_3_lut_LC_13_3_5  (
            .in0(N__34995),
            .in1(_gnd_net_),
            .in2(N__32416),
            .in3(N__37424),
            .lcout(\comm_spi.imosi ),
            .ltout(\comm_spi.imosi_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_86_2_lut_LC_13_3_6 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_86_2_lut_LC_13_3_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_86_2_lut_LC_13_3_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \comm_spi.RESET_I_0_86_2_lut_LC_13_3_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32413),
            .in3(N__55465),
            .lcout(\comm_spi.DOUT_7__N_738 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_87_2_lut_LC_13_3_7 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_87_2_lut_LC_13_3_7 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_87_2_lut_LC_13_3_7 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \comm_spi.RESET_I_0_87_2_lut_LC_13_3_7  (
            .in0(N__32410),
            .in1(_gnd_net_),
            .in2(N__55473),
            .in3(_gnd_net_),
            .lcout(\comm_spi.DOUT_7__N_739 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_rx_i0_12197_12198_set_LC_13_4_0 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i0_12197_12198_set_LC_13_4_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_rx_i0_12197_12198_set_LC_13_4_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.data_rx_i0_12197_12198_set_LC_13_4_0  (
            .in0(N__37426),
            .in1(N__34994),
            .in2(_gnd_net_),
            .in3(N__33820),
            .lcout(\comm_spi.n14599 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52364),
            .ce(),
            .sr(N__32395));
    defparam \ADC_VDC.genclk.div_state_1__I_0_1_lut_LC_13_5_0 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.div_state_1__I_0_1_lut_LC_13_5_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.div_state_1__I_0_1_lut_LC_13_5_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \ADC_VDC.genclk.div_state_1__I_0_1_lut_LC_13_5_0  (
            .in0(N__34913),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\ADC_VDC.genclk.div_state_1__N_1266 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i19148_2_lut_4_lut_LC_13_5_2 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i19148_2_lut_4_lut_LC_13_5_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i19148_2_lut_4_lut_LC_13_5_2 .LUT_INIT=16'b0001111110111111;
    LogicCell40 \ADC_VDC.genclk.i19148_2_lut_4_lut_LC_13_5_2  (
            .in0(N__34914),
            .in1(N__33780),
            .in2(N__34975),
            .in3(N__32382),
            .lcout(\ADC_VDC.genclk.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i19194_4_lut_3_lut_LC_13_5_3 .C_ON=1'b0;
    defparam \comm_spi.i19194_4_lut_3_lut_LC_13_5_3 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19194_4_lut_3_lut_LC_13_5_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.i19194_4_lut_3_lut_LC_13_5_3  (
            .in0(N__55458),
            .in1(N__48737),
            .in2(_gnd_net_),
            .in3(N__43562),
            .lcout(\comm_spi.n22635 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i24_4_lut_LC_13_5_5 .C_ON=1'b0;
    defparam \ADC_VDC.i24_4_lut_LC_13_5_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i24_4_lut_LC_13_5_5 .LUT_INIT=16'b1111001100001010;
    LogicCell40 \ADC_VDC.i24_4_lut_LC_13_5_5  (
            .in0(N__34648),
            .in1(N__34154),
            .in2(N__34384),
            .in3(N__34466),
            .lcout(),
            .ltout(\ADC_VDC.n11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_4_lut_LC_13_5_6 .C_ON=1'b0;
    defparam \ADC_VDC.i1_4_lut_LC_13_5_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_4_lut_LC_13_5_6 .LUT_INIT=16'b1110000011110000;
    LogicCell40 \ADC_VDC.i1_4_lut_LC_13_5_6  (
            .in0(N__34360),
            .in1(N__32557),
            .in2(N__32560),
            .in3(N__34769),
            .lcout(\ADC_VDC.n18381 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i14977_2_lut_LC_13_5_7 .C_ON=1'b0;
    defparam \ADC_VDC.i14977_2_lut_LC_13_5_7 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i14977_2_lut_LC_13_5_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ADC_VDC.i14977_2_lut_LC_13_5_7  (
            .in0(_gnd_net_),
            .in1(N__34465),
            .in2(_gnd_net_),
            .in3(N__34153),
            .lcout(\ADC_VDC.n17359 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.bit_cnt_3769__i0_LC_13_6_0 .C_ON=1'b1;
    defparam \ADC_VDC.bit_cnt_3769__i0_LC_13_6_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3769__i0_LC_13_6_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3769__i0_LC_13_6_0  (
            .in0(_gnd_net_),
            .in1(N__32547),
            .in2(_gnd_net_),
            .in3(N__32518),
            .lcout(\ADC_VDC.bit_cnt_0 ),
            .ltout(),
            .carryin(bfn_13_6_0_),
            .carryout(\ADC_VDC.n19469 ),
            .clk(N__32727),
            .ce(N__34012),
            .sr(N__32671));
    defparam \ADC_VDC.bit_cnt_3769__i1_LC_13_6_1 .C_ON=1'b1;
    defparam \ADC_VDC.bit_cnt_3769__i1_LC_13_6_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3769__i1_LC_13_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3769__i1_LC_13_6_1  (
            .in0(_gnd_net_),
            .in1(N__32510),
            .in2(_gnd_net_),
            .in3(N__32479),
            .lcout(\ADC_VDC.bit_cnt_1 ),
            .ltout(),
            .carryin(\ADC_VDC.n19469 ),
            .carryout(\ADC_VDC.n19470 ),
            .clk(N__32727),
            .ce(N__34012),
            .sr(N__32671));
    defparam \ADC_VDC.bit_cnt_3769__i2_LC_13_6_2 .C_ON=1'b1;
    defparam \ADC_VDC.bit_cnt_3769__i2_LC_13_6_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3769__i2_LC_13_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3769__i2_LC_13_6_2  (
            .in0(_gnd_net_),
            .in1(N__32595),
            .in2(_gnd_net_),
            .in3(N__32476),
            .lcout(\ADC_VDC.bit_cnt_2 ),
            .ltout(),
            .carryin(\ADC_VDC.n19470 ),
            .carryout(\ADC_VDC.n19471 ),
            .clk(N__32727),
            .ce(N__34012),
            .sr(N__32671));
    defparam \ADC_VDC.bit_cnt_3769__i3_LC_13_6_3 .C_ON=1'b1;
    defparam \ADC_VDC.bit_cnt_3769__i3_LC_13_6_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3769__i3_LC_13_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3769__i3_LC_13_6_3  (
            .in0(_gnd_net_),
            .in1(N__32633),
            .in2(_gnd_net_),
            .in3(N__32473),
            .lcout(\ADC_VDC.bit_cnt_3 ),
            .ltout(),
            .carryin(\ADC_VDC.n19471 ),
            .carryout(\ADC_VDC.n19472 ),
            .clk(N__32727),
            .ce(N__34012),
            .sr(N__32671));
    defparam \ADC_VDC.bit_cnt_3769__i4_LC_13_6_4 .C_ON=1'b1;
    defparam \ADC_VDC.bit_cnt_3769__i4_LC_13_6_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3769__i4_LC_13_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3769__i4_LC_13_6_4  (
            .in0(_gnd_net_),
            .in1(N__32466),
            .in2(_gnd_net_),
            .in3(N__32440),
            .lcout(\ADC_VDC.bit_cnt_4 ),
            .ltout(),
            .carryin(\ADC_VDC.n19472 ),
            .carryout(\ADC_VDC.n19473 ),
            .clk(N__32727),
            .ce(N__34012),
            .sr(N__32671));
    defparam \ADC_VDC.bit_cnt_3769__i5_LC_13_6_5 .C_ON=1'b1;
    defparam \ADC_VDC.bit_cnt_3769__i5_LC_13_6_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3769__i5_LC_13_6_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3769__i5_LC_13_6_5  (
            .in0(_gnd_net_),
            .in1(N__32437),
            .in2(_gnd_net_),
            .in3(N__32419),
            .lcout(\ADC_VDC.bit_cnt_5 ),
            .ltout(),
            .carryin(\ADC_VDC.n19473 ),
            .carryout(\ADC_VDC.n19474 ),
            .clk(N__32727),
            .ce(N__34012),
            .sr(N__32671));
    defparam \ADC_VDC.bit_cnt_3769__i6_LC_13_6_6 .C_ON=1'b1;
    defparam \ADC_VDC.bit_cnt_3769__i6_LC_13_6_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3769__i6_LC_13_6_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3769__i6_LC_13_6_6  (
            .in0(_gnd_net_),
            .in1(N__32953),
            .in2(_gnd_net_),
            .in3(N__32938),
            .lcout(\ADC_VDC.bit_cnt_6 ),
            .ltout(),
            .carryin(\ADC_VDC.n19474 ),
            .carryout(\ADC_VDC.n19475 ),
            .clk(N__32727),
            .ce(N__34012),
            .sr(N__32671));
    defparam \ADC_VDC.bit_cnt_3769__i7_LC_13_6_7 .C_ON=1'b0;
    defparam \ADC_VDC.bit_cnt_3769__i7_LC_13_6_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3769__i7_LC_13_6_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3769__i7_LC_13_6_7  (
            .in0(_gnd_net_),
            .in1(N__32932),
            .in2(_gnd_net_),
            .in3(N__32935),
            .lcout(\ADC_VDC.bit_cnt_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32727),
            .ce(N__34012),
            .sr(N__32671));
    defparam \comm_spi.imiso_83_12193_12194_set_LC_13_7_0 .C_ON=1'b0;
    defparam \comm_spi.imiso_83_12193_12194_set_LC_13_7_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.imiso_83_12193_12194_set_LC_13_7_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \comm_spi.imiso_83_12193_12194_set_LC_13_7_0  (
            .in0(N__40213),
            .in1(N__44272),
            .in2(_gnd_net_),
            .in3(N__40192),
            .lcout(\comm_spi.n14595 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.imiso_83_12193_12194_setC_net ),
            .ce(),
            .sr(N__40261));
    defparam mux_130_Mux_6_i30_3_lut_LC_13_7_4.C_ON=1'b0;
    defparam mux_130_Mux_6_i30_3_lut_LC_13_7_4.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_6_i30_3_lut_LC_13_7_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_130_Mux_6_i30_3_lut_LC_13_7_4 (
            .in0(N__32659),
            .in1(N__41215),
            .in2(_gnd_net_),
            .in3(N__56256),
            .lcout(n30_adj_1595),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_2_lut_adj_33_LC_13_7_5 .C_ON=1'b0;
    defparam \ADC_VDC.i1_2_lut_adj_33_LC_13_7_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_2_lut_adj_33_LC_13_7_5 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \ADC_VDC.i1_2_lut_adj_33_LC_13_7_5  (
            .in0(_gnd_net_),
            .in1(N__32625),
            .in2(_gnd_net_),
            .in3(N__32591),
            .lcout(\ADC_VDC.n6_adj_1404 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_104_2_lut_LC_13_7_6 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_104_2_lut_LC_13_7_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_104_2_lut_LC_13_7_6 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \comm_spi.RESET_I_0_104_2_lut_LC_13_7_6  (
            .in0(N__55461),
            .in1(N__37628),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\comm_spi.data_tx_7__N_778 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_96_2_lut_LC_13_7_7 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_96_2_lut_LC_13_7_7 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_96_2_lut_LC_13_7_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \comm_spi.RESET_I_0_96_2_lut_LC_13_7_7  (
            .in0(N__37629),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55462),
            .lcout(\comm_spi.data_tx_7__N_762 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i3_12209_12210_set_LC_13_8_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i3_12209_12210_set_LC_13_8_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i3_12209_12210_set_LC_13_8_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \comm_spi.data_tx_i3_12209_12210_set_LC_13_8_0  (
            .in0(N__37666),
            .in1(N__37726),
            .in2(_gnd_net_),
            .in3(N__37693),
            .lcout(\comm_spi.n14611 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52425),
            .ce(),
            .sr(N__33049));
    defparam i9327_1_lut_LC_13_8_2.C_ON=1'b0;
    defparam i9327_1_lut_LC_13_8_2.SEQ_MODE=4'b0000;
    defparam i9327_1_lut_LC_13_8_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 i9327_1_lut_LC_13_8_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50255),
            .lcout(n11727),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.bit_cnt_3767__i1_LC_13_9_2 .C_ON=1'b0;
    defparam \comm_spi.bit_cnt_3767__i1_LC_13_9_2 .SEQ_MODE=4'b1010;
    defparam \comm_spi.bit_cnt_3767__i1_LC_13_9_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \comm_spi.bit_cnt_3767__i1_LC_13_9_2  (
            .in0(N__33010),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33032),
            .lcout(\comm_spi.bit_cnt_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.bit_cnt_3767__i1C_net ),
            .ce(),
            .sr(N__55437));
    defparam \comm_spi.bit_cnt_3767__i0_LC_13_9_3 .C_ON=1'b0;
    defparam \comm_spi.bit_cnt_3767__i0_LC_13_9_3 .SEQ_MODE=4'b1010;
    defparam \comm_spi.bit_cnt_3767__i0_LC_13_9_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \comm_spi.bit_cnt_3767__i0_LC_13_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33009),
            .lcout(\comm_spi.bit_cnt_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.bit_cnt_3767__i1C_net ),
            .ce(),
            .sr(N__55437));
    defparam \comm_spi.bit_cnt_3767__i3_LC_13_9_6 .C_ON=1'b0;
    defparam \comm_spi.bit_cnt_3767__i3_LC_13_9_6 .SEQ_MODE=4'b1010;
    defparam \comm_spi.bit_cnt_3767__i3_LC_13_9_6 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \comm_spi.bit_cnt_3767__i3_LC_13_9_6  (
            .in0(N__32988),
            .in1(N__46377),
            .in2(N__33016),
            .in3(N__33034),
            .lcout(\comm_spi.bit_cnt_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.bit_cnt_3767__i1C_net ),
            .ce(),
            .sr(N__55437));
    defparam \comm_spi.bit_cnt_3767__i2_LC_13_9_7 .C_ON=1'b0;
    defparam \comm_spi.bit_cnt_3767__i2_LC_13_9_7 .SEQ_MODE=4'b1010;
    defparam \comm_spi.bit_cnt_3767__i2_LC_13_9_7 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \comm_spi.bit_cnt_3767__i2_LC_13_9_7  (
            .in0(N__33033),
            .in1(N__33011),
            .in2(_gnd_net_),
            .in3(N__32987),
            .lcout(\comm_spi.bit_cnt_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.bit_cnt_3767__i1C_net ),
            .ce(),
            .sr(N__55437));
    defparam i1_2_lut_3_lut_adj_275_LC_13_10_0.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_275_LC_13_10_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_275_LC_13_10_0.LUT_INIT=16'b1011101111111111;
    LogicCell40 i1_2_lut_3_lut_adj_275_LC_13_10_0 (
            .in0(N__54387),
            .in1(N__51210),
            .in2(_gnd_net_),
            .in3(N__53901),
            .lcout(n20653),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15208_2_lut_3_lut_LC_13_10_1.C_ON=1'b0;
    defparam i15208_2_lut_3_lut_LC_13_10_1.SEQ_MODE=4'b0000;
    defparam i15208_2_lut_3_lut_LC_13_10_1.LUT_INIT=16'b0000010000000100;
    LogicCell40 i15208_2_lut_3_lut_LC_13_10_1 (
            .in0(N__53903),
            .in1(N__42804),
            .in2(N__51261),
            .in3(_gnd_net_),
            .lcout(n14_adj_1528),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i2_3_lut_LC_13_10_2 .C_ON=1'b0;
    defparam \comm_spi.i2_3_lut_LC_13_10_2 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i2_3_lut_LC_13_10_2 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \comm_spi.i2_3_lut_LC_13_10_2  (
            .in0(N__33031),
            .in1(N__33015),
            .in2(_gnd_net_),
            .in3(N__32989),
            .lcout(\comm_spi.n16858 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_0__bdd_4_lut_LC_13_10_3.C_ON=1'b0;
    defparam comm_index_0__bdd_4_lut_LC_13_10_3.SEQ_MODE=4'b0000;
    defparam comm_index_0__bdd_4_lut_LC_13_10_3.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_index_0__bdd_4_lut_LC_13_10_3 (
            .in0(N__35149),
            .in1(N__49520),
            .in2(N__32971),
            .in3(N__51623),
            .lcout(),
            .ltout(n21991_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n21991_bdd_4_lut_LC_13_10_4.C_ON=1'b0;
    defparam n21991_bdd_4_lut_LC_13_10_4.SEQ_MODE=4'b0000;
    defparam n21991_bdd_4_lut_LC_13_10_4.LUT_INIT=16'b1110010111100000;
    LogicCell40 n21991_bdd_4_lut_LC_13_10_4 (
            .in0(N__49521),
            .in1(N__43383),
            .in2(N__32956),
            .in3(N__44112),
            .lcout(n21994),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12366_2_lut_LC_13_10_5.C_ON=1'b0;
    defparam i12366_2_lut_LC_13_10_5.SEQ_MODE=4'b0000;
    defparam i12366_2_lut_LC_13_10_5.LUT_INIT=16'b1100110000000000;
    LogicCell40 i12366_2_lut_LC_13_10_5 (
            .in0(_gnd_net_),
            .in1(N__54388),
            .in2(_gnd_net_),
            .in3(N__49821),
            .lcout(n14763),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15190_2_lut_3_lut_LC_13_10_6.C_ON=1'b0;
    defparam i15190_2_lut_3_lut_LC_13_10_6.SEQ_MODE=4'b0000;
    defparam i15190_2_lut_3_lut_LC_13_10_6.LUT_INIT=16'b0000000000100010;
    LogicCell40 i15190_2_lut_3_lut_LC_13_10_6 (
            .in0(N__36394),
            .in1(N__51217),
            .in2(_gnd_net_),
            .in3(N__53904),
            .lcout(n14_adj_1558),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15207_2_lut_3_lut_LC_13_10_7.C_ON=1'b0;
    defparam i15207_2_lut_3_lut_LC_13_10_7.SEQ_MODE=4'b0000;
    defparam i15207_2_lut_3_lut_LC_13_10_7.LUT_INIT=16'b0000010000000100;
    LogicCell40 i15207_2_lut_3_lut_LC_13_10_7 (
            .in0(N__53902),
            .in1(N__46646),
            .in2(N__51260),
            .in3(_gnd_net_),
            .lcout(n14_adj_1527),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_0__bdd_4_lut_19374_LC_13_11_0.C_ON=1'b0;
    defparam comm_index_0__bdd_4_lut_19374_LC_13_11_0.SEQ_MODE=4'b0000;
    defparam comm_index_0__bdd_4_lut_19374_LC_13_11_0.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_index_0__bdd_4_lut_19374_LC_13_11_0 (
            .in0(N__35191),
            .in1(N__49530),
            .in2(N__33100),
            .in3(N__51624),
            .lcout(),
            .ltout(n21979_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n21979_bdd_4_lut_LC_13_11_1.C_ON=1'b0;
    defparam n21979_bdd_4_lut_LC_13_11_1.SEQ_MODE=4'b0000;
    defparam n21979_bdd_4_lut_LC_13_11_1.LUT_INIT=16'b1111010010100100;
    LogicCell40 n21979_bdd_4_lut_LC_13_11_1 (
            .in0(N__49531),
            .in1(N__43768),
            .in2(N__33085),
            .in3(N__36395),
            .lcout(n21982),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_137_Mux_3_i4_3_lut_LC_13_11_2.C_ON=1'b0;
    defparam mux_137_Mux_3_i4_3_lut_LC_13_11_2.SEQ_MODE=4'b0000;
    defparam mux_137_Mux_3_i4_3_lut_LC_13_11_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_137_Mux_3_i4_3_lut_LC_13_11_2 (
            .in0(N__35461),
            .in1(N__33082),
            .in2(_gnd_net_),
            .in3(N__51625),
            .lcout(),
            .ltout(n4_adj_1567_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18188_4_lut_LC_13_11_3.C_ON=1'b0;
    defparam i18188_4_lut_LC_13_11_3.SEQ_MODE=4'b0000;
    defparam i18188_4_lut_LC_13_11_3.LUT_INIT=16'b0100010011110000;
    LogicCell40 i18188_4_lut_LC_13_11_3 (
            .in0(N__51626),
            .in1(N__33076),
            .in2(N__33061),
            .in3(N__49534),
            .lcout(),
            .ltout(n20783_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i3_LC_13_11_4.C_ON=1'b0;
    defparam comm_tx_buf_i3_LC_13_11_4.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i3_LC_13_11_4.LUT_INIT=16'b1111010110100000;
    LogicCell40 comm_tx_buf_i3_LC_13_11_4 (
            .in0(N__50069),
            .in1(_gnd_net_),
            .in2(N__33058),
            .in3(N__33055),
            .lcout(comm_tx_buf_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55098),
            .ce(N__47128),
            .sr(N__47061));
    defparam i14948_3_lut_LC_13_11_5.C_ON=1'b0;
    defparam i14948_3_lut_LC_13_11_5.SEQ_MODE=4'b0000;
    defparam i14948_3_lut_LC_13_11_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 i14948_3_lut_LC_13_11_5 (
            .in0(N__35674),
            .in1(N__50182),
            .in2(_gnd_net_),
            .in3(N__50067),
            .lcout(),
            .ltout(n17331_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18308_4_lut_LC_13_11_6.C_ON=1'b0;
    defparam i18308_4_lut_LC_13_11_6.SEQ_MODE=4'b0000;
    defparam i18308_4_lut_LC_13_11_6.LUT_INIT=16'b0100010011110000;
    LogicCell40 i18308_4_lut_LC_13_11_6 (
            .in0(N__50068),
            .in1(N__33190),
            .in2(N__33175),
            .in3(N__49532),
            .lcout(),
            .ltout(n20903_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i5_LC_13_11_7.C_ON=1'b0;
    defparam comm_tx_buf_i5_LC_13_11_7.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i5_LC_13_11_7.LUT_INIT=16'b1111010110100000;
    LogicCell40 comm_tx_buf_i5_LC_13_11_7 (
            .in0(N__51627),
            .in1(_gnd_net_),
            .in2(N__33172),
            .in3(N__38221),
            .lcout(comm_tx_buf_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55098),
            .ce(N__47128),
            .sr(N__47061));
    defparam mux_137_Mux_6_i1_3_lut_LC_13_12_0.C_ON=1'b0;
    defparam mux_137_Mux_6_i1_3_lut_LC_13_12_0.SEQ_MODE=4'b0000;
    defparam mux_137_Mux_6_i1_3_lut_LC_13_12_0.LUT_INIT=16'b1100110010101010;
    LogicCell40 mux_137_Mux_6_i1_3_lut_LC_13_12_0 (
            .in0(N__40785),
            .in1(N__51428),
            .in2(_gnd_net_),
            .in3(N__51631),
            .lcout(),
            .ltout(n1_adj_1561_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i6_LC_13_12_1.C_ON=1'b0;
    defparam comm_tx_buf_i6_LC_13_12_1.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i6_LC_13_12_1.LUT_INIT=16'b1010101011011000;
    LogicCell40 comm_tx_buf_i6_LC_13_12_1 (
            .in0(N__33112),
            .in1(N__33133),
            .in2(N__33169),
            .in3(N__50099),
            .lcout(comm_tx_buf_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55107),
            .ce(N__47140),
            .sr(N__47065));
    defparam i18895_2_lut_LC_13_12_2.C_ON=1'b0;
    defparam i18895_2_lut_LC_13_12_2.SEQ_MODE=4'b0000;
    defparam i18895_2_lut_LC_13_12_2.LUT_INIT=16'b0000000011001100;
    LogicCell40 i18895_2_lut_LC_13_12_2 (
            .in0(_gnd_net_),
            .in1(N__33162),
            .in2(_gnd_net_),
            .in3(N__51628),
            .lcout(n21051),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_137_Mux_6_i2_3_lut_LC_13_12_3.C_ON=1'b0;
    defparam mux_137_Mux_6_i2_3_lut_LC_13_12_3.SEQ_MODE=4'b0000;
    defparam mux_137_Mux_6_i2_3_lut_LC_13_12_3.LUT_INIT=16'b1111010110100000;
    LogicCell40 mux_137_Mux_6_i2_3_lut_LC_13_12_3 (
            .in0(N__51630),
            .in1(_gnd_net_),
            .in2(N__33148),
            .in3(N__35212),
            .lcout(n2_adj_1562),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_137_Mux_6_i4_3_lut_LC_13_12_4.C_ON=1'b0;
    defparam mux_137_Mux_6_i4_3_lut_LC_13_12_4.SEQ_MODE=4'b0000;
    defparam mux_137_Mux_6_i4_3_lut_LC_13_12_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_137_Mux_6_i4_3_lut_LC_13_12_4 (
            .in0(N__35701),
            .in1(N__33127),
            .in2(_gnd_net_),
            .in3(N__51629),
            .lcout(),
            .ltout(n4_adj_1563_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_1__bdd_4_lut_19472_LC_13_12_5.C_ON=1'b0;
    defparam comm_index_1__bdd_4_lut_19472_LC_13_12_5.SEQ_MODE=4'b0000;
    defparam comm_index_1__bdd_4_lut_19472_LC_13_12_5.LUT_INIT=16'b1101100010101010;
    LogicCell40 comm_index_1__bdd_4_lut_19472_LC_13_12_5 (
            .in0(N__49533),
            .in1(N__33121),
            .in2(N__33115),
            .in3(N__50098),
            .lcout(n22093),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_101_2_lut_LC_13_12_6 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_101_2_lut_LC_13_12_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_101_2_lut_LC_13_12_6 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \comm_spi.RESET_I_0_101_2_lut_LC_13_12_6  (
            .in0(N__55459),
            .in1(N__40274),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\comm_spi.data_tx_7__N_769 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_93_2_lut_LC_13_12_7 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_93_2_lut_LC_13_12_7 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_93_2_lut_LC_13_12_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \comm_spi.RESET_I_0_93_2_lut_LC_13_12_7  (
            .in0(N__40275),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55460),
            .lcout(\comm_spi.data_tx_7__N_759 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_2_i26_3_lut_LC_13_13_0.C_ON=1'b0;
    defparam mux_129_Mux_2_i26_3_lut_LC_13_13_0.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_2_i26_3_lut_LC_13_13_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_129_Mux_2_i26_3_lut_LC_13_13_0 (
            .in0(N__33336),
            .in1(N__56832),
            .in2(_gnd_net_),
            .in3(N__46882),
            .lcout(),
            .ltout(n26_adj_1506_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18221_4_lut_LC_13_13_1.C_ON=1'b0;
    defparam i18221_4_lut_LC_13_13_1.SEQ_MODE=4'b0000;
    defparam i18221_4_lut_LC_13_13_1.LUT_INIT=16'b0111010000110000;
    LogicCell40 i18221_4_lut_LC_13_13_1 (
            .in0(N__56833),
            .in1(N__57482),
            .in2(N__33325),
            .in3(N__33322),
            .lcout(),
            .ltout(n20816_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_2__bdd_4_lut_19561_LC_13_13_2.C_ON=1'b0;
    defparam comm_cmd_2__bdd_4_lut_19561_LC_13_13_2.SEQ_MODE=4'b0000;
    defparam comm_cmd_2__bdd_4_lut_19561_LC_13_13_2.LUT_INIT=16'b1110010010101010;
    LogicCell40 comm_cmd_2__bdd_4_lut_19561_LC_13_13_2 (
            .in0(N__47788),
            .in1(N__33238),
            .in2(N__33304),
            .in3(N__56289),
            .lcout(),
            .ltout(n22087_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22087_bdd_4_lut_LC_13_13_3.C_ON=1'b0;
    defparam n22087_bdd_4_lut_LC_13_13_3.SEQ_MODE=4'b0000;
    defparam n22087_bdd_4_lut_LC_13_13_3.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22087_bdd_4_lut_LC_13_13_3 (
            .in0(N__56290),
            .in1(N__33301),
            .in2(N__33286),
            .in3(N__33244),
            .lcout(),
            .ltout(n22090_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i2_LC_13_13_4.C_ON=1'b0;
    defparam comm_buf_1__i2_LC_13_13_4.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i2_LC_13_13_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 comm_buf_1__i2_LC_13_13_4 (
            .in0(_gnd_net_),
            .in1(N__35452),
            .in2(N__33283),
            .in3(N__53908),
            .lcout(comm_buf_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55118),
            .ce(N__38544),
            .sr(N__36807));
    defparam i18251_3_lut_LC_13_13_6.C_ON=1'b0;
    defparam i18251_3_lut_LC_13_13_6.SEQ_MODE=4'b0000;
    defparam i18251_3_lut_LC_13_13_6.LUT_INIT=16'b1100110010101010;
    LogicCell40 i18251_3_lut_LC_13_13_6 (
            .in0(N__33280),
            .in1(N__33271),
            .in2(_gnd_net_),
            .in3(N__57481),
            .lcout(n20846),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18220_3_lut_LC_13_13_7.C_ON=1'b0;
    defparam i18220_3_lut_LC_13_13_7.SEQ_MODE=4'b0000;
    defparam i18220_3_lut_LC_13_13_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 i18220_3_lut_LC_13_13_7 (
            .in0(N__57480),
            .in1(N__41596),
            .in2(_gnd_net_),
            .in3(N__36304),
            .lcout(n20815),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19477_LC_13_14_0.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19477_LC_13_14_0.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19477_LC_13_14_0.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_19477_LC_13_14_0 (
            .in0(N__33232),
            .in1(N__57532),
            .in2(N__33217),
            .in3(N__47782),
            .lcout(),
            .ltout(n22081_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22081_bdd_4_lut_LC_13_14_1.C_ON=1'b0;
    defparam n22081_bdd_4_lut_LC_13_14_1.SEQ_MODE=4'b0000;
    defparam n22081_bdd_4_lut_LC_13_14_1.LUT_INIT=16'b1110010111100000;
    LogicCell40 n22081_bdd_4_lut_LC_13_14_1 (
            .in0(N__47783),
            .in1(N__33469),
            .in2(N__33442),
            .in3(N__36124),
            .lcout(n22084),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_4_i26_3_lut_LC_13_14_2.C_ON=1'b0;
    defparam mux_129_Mux_4_i26_3_lut_LC_13_14_2.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_4_i26_3_lut_LC_13_14_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_129_Mux_4_i26_3_lut_LC_13_14_2 (
            .in0(N__33438),
            .in1(N__56840),
            .in2(_gnd_net_),
            .in3(N__46813),
            .lcout(),
            .ltout(n26_adj_1484_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19531_LC_13_14_3.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19531_LC_13_14_3.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19531_LC_13_14_3.LUT_INIT=16'b1101110110100000;
    LogicCell40 comm_cmd_1__bdd_4_lut_19531_LC_13_14_3 (
            .in0(N__47784),
            .in1(N__33421),
            .in2(N__33409),
            .in3(N__57483),
            .lcout(),
            .ltout(n22159_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22159_bdd_4_lut_LC_13_14_4.C_ON=1'b0;
    defparam n22159_bdd_4_lut_LC_13_14_4.SEQ_MODE=4'b0000;
    defparam n22159_bdd_4_lut_LC_13_14_4.LUT_INIT=16'b1111001011000010;
    LogicCell40 n22159_bdd_4_lut_LC_13_14_4 (
            .in0(N__36949),
            .in1(N__47785),
            .in2(N__33406),
            .in3(N__38395),
            .lcout(),
            .ltout(n22162_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1541671_i1_3_lut_LC_13_14_5.C_ON=1'b0;
    defparam i1541671_i1_3_lut_LC_13_14_5.SEQ_MODE=4'b0000;
    defparam i1541671_i1_3_lut_LC_13_14_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 i1541671_i1_3_lut_LC_13_14_5 (
            .in0(_gnd_net_),
            .in1(N__33403),
            .in2(N__33397),
            .in3(N__56287),
            .lcout(),
            .ltout(n30_adj_1493_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i4_LC_13_14_6.C_ON=1'b0;
    defparam comm_buf_1__i4_LC_13_14_6.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i4_LC_13_14_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 comm_buf_1__i4_LC_13_14_6 (
            .in0(_gnd_net_),
            .in1(N__35661),
            .in2(N__33394),
            .in3(N__54000),
            .lcout(comm_buf_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55127),
            .ce(N__38550),
            .sr(N__36790));
    defparam mux_129_Mux_3_i26_3_lut_LC_13_15_0.C_ON=1'b0;
    defparam mux_129_Mux_3_i26_3_lut_LC_13_15_0.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_3_i26_3_lut_LC_13_15_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_129_Mux_3_i26_3_lut_LC_13_15_0 (
            .in0(N__56841),
            .in1(N__33391),
            .in2(_gnd_net_),
            .in3(N__46851),
            .lcout(),
            .ltout(n26_adj_1502_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_LC_13_15_1.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_LC_13_15_1.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_LC_13_15_1.LUT_INIT=16'b1011101111000000;
    LogicCell40 comm_cmd_1__bdd_4_lut_LC_13_15_1 (
            .in0(N__33376),
            .in1(N__47780),
            .in2(N__33361),
            .in3(N__57550),
            .lcout(),
            .ltout(n22195_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22195_bdd_4_lut_LC_13_15_2.C_ON=1'b0;
    defparam n22195_bdd_4_lut_LC_13_15_2.SEQ_MODE=4'b0000;
    defparam n22195_bdd_4_lut_LC_13_15_2.LUT_INIT=16'b1110010111100000;
    LogicCell40 n22195_bdd_4_lut_LC_13_15_2 (
            .in0(N__47781),
            .in1(N__38833),
            .in2(N__33358),
            .in3(N__33355),
            .lcout(),
            .ltout(n22198_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1540465_i1_3_lut_LC_13_15_3.C_ON=1'b0;
    defparam i1540465_i1_3_lut_LC_13_15_3.SEQ_MODE=4'b0000;
    defparam i1540465_i1_3_lut_LC_13_15_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 i1540465_i1_3_lut_LC_13_15_3 (
            .in0(_gnd_net_),
            .in1(N__33502),
            .in2(N__33589),
            .in3(N__56288),
            .lcout(),
            .ltout(n30_adj_1503_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i3_LC_13_15_4.C_ON=1'b0;
    defparam comm_buf_1__i3_LC_13_15_4.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i3_LC_13_15_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 comm_buf_1__i3_LC_13_15_4 (
            .in0(_gnd_net_),
            .in1(N__35569),
            .in2(N__33586),
            .in3(N__53909),
            .lcout(comm_buf_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55139),
            .ce(N__38545),
            .sr(N__36796));
    defparam comm_cmd_1__bdd_4_lut_19403_LC_13_15_5.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19403_LC_13_15_5.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19403_LC_13_15_5.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_1__bdd_4_lut_19403_LC_13_15_5 (
            .in0(N__33583),
            .in1(N__47778),
            .in2(N__33571),
            .in3(N__57549),
            .lcout(),
            .ltout(n22009_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22009_bdd_4_lut_LC_13_15_6.C_ON=1'b0;
    defparam n22009_bdd_4_lut_LC_13_15_6.SEQ_MODE=4'b0000;
    defparam n22009_bdd_4_lut_LC_13_15_6.LUT_INIT=16'b1110010111100000;
    LogicCell40 n22009_bdd_4_lut_LC_13_15_6 (
            .in0(N__47779),
            .in1(N__33541),
            .in2(N__33514),
            .in3(N__33511),
            .lcout(n22012),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipcnt_i0_i0_LC_13_16_0.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i0_LC_13_16_0.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i0_LC_13_16_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i0_LC_13_16_0 (
            .in0(_gnd_net_),
            .in1(N__46956),
            .in2(N__33496),
            .in3(_gnd_net_),
            .lcout(acadc_skipcnt_0),
            .ltout(),
            .carryin(bfn_13_16_0_),
            .carryout(n19311),
            .clk(INVacadc_skipcnt_i0_i0C_net),
            .ce(N__33936),
            .sr(N__33481));
    defparam add_73_2_THRU_CRY_0_LC_13_16_1.C_ON=1'b1;
    defparam add_73_2_THRU_CRY_0_LC_13_16_1.SEQ_MODE=4'b0000;
    defparam add_73_2_THRU_CRY_0_LC_13_16_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_73_2_THRU_CRY_0_LC_13_16_1 (
            .in0(_gnd_net_),
            .in1(N__52799),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n19311),
            .carryout(n19311_THRU_CRY_0_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_73_2_THRU_CRY_1_LC_13_16_2.C_ON=1'b1;
    defparam add_73_2_THRU_CRY_1_LC_13_16_2.SEQ_MODE=4'b0000;
    defparam add_73_2_THRU_CRY_1_LC_13_16_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_73_2_THRU_CRY_1_LC_13_16_2 (
            .in0(_gnd_net_),
            .in1(N__52803),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n19311_THRU_CRY_0_THRU_CO),
            .carryout(n19311_THRU_CRY_1_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_73_2_THRU_CRY_2_LC_13_16_3.C_ON=1'b1;
    defparam add_73_2_THRU_CRY_2_LC_13_16_3.SEQ_MODE=4'b0000;
    defparam add_73_2_THRU_CRY_2_LC_13_16_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_73_2_THRU_CRY_2_LC_13_16_3 (
            .in0(_gnd_net_),
            .in1(N__52800),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n19311_THRU_CRY_1_THRU_CO),
            .carryout(n19311_THRU_CRY_2_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_73_2_THRU_CRY_3_LC_13_16_4.C_ON=1'b1;
    defparam add_73_2_THRU_CRY_3_LC_13_16_4.SEQ_MODE=4'b0000;
    defparam add_73_2_THRU_CRY_3_LC_13_16_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_73_2_THRU_CRY_3_LC_13_16_4 (
            .in0(_gnd_net_),
            .in1(N__52804),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n19311_THRU_CRY_2_THRU_CO),
            .carryout(n19311_THRU_CRY_3_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_73_2_THRU_CRY_4_LC_13_16_5.C_ON=1'b1;
    defparam add_73_2_THRU_CRY_4_LC_13_16_5.SEQ_MODE=4'b0000;
    defparam add_73_2_THRU_CRY_4_LC_13_16_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_73_2_THRU_CRY_4_LC_13_16_5 (
            .in0(_gnd_net_),
            .in1(N__52801),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n19311_THRU_CRY_3_THRU_CO),
            .carryout(n19311_THRU_CRY_4_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_73_2_THRU_CRY_5_LC_13_16_6.C_ON=1'b1;
    defparam add_73_2_THRU_CRY_5_LC_13_16_6.SEQ_MODE=4'b0000;
    defparam add_73_2_THRU_CRY_5_LC_13_16_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_73_2_THRU_CRY_5_LC_13_16_6 (
            .in0(_gnd_net_),
            .in1(N__52805),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n19311_THRU_CRY_4_THRU_CO),
            .carryout(n19311_THRU_CRY_5_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_73_2_THRU_CRY_6_LC_13_16_7.C_ON=1'b1;
    defparam add_73_2_THRU_CRY_6_LC_13_16_7.SEQ_MODE=4'b0000;
    defparam add_73_2_THRU_CRY_6_LC_13_16_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_73_2_THRU_CRY_6_LC_13_16_7 (
            .in0(_gnd_net_),
            .in1(N__52802),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n19311_THRU_CRY_5_THRU_CO),
            .carryout(n19311_THRU_CRY_6_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipcnt_i0_i1_LC_13_17_0.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i1_LC_13_17_0.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i1_LC_13_17_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i1_LC_13_17_0 (
            .in0(_gnd_net_),
            .in1(N__33675),
            .in2(_gnd_net_),
            .in3(N__33661),
            .lcout(acadc_skipcnt_1),
            .ltout(),
            .carryin(bfn_13_17_0_),
            .carryout(n19312),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__33923),
            .sr(N__33894));
    defparam acadc_skipcnt_i0_i2_LC_13_17_1.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i2_LC_13_17_1.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i2_LC_13_17_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i2_LC_13_17_1 (
            .in0(_gnd_net_),
            .in1(N__36333),
            .in2(_gnd_net_),
            .in3(N__33658),
            .lcout(acadc_skipcnt_2),
            .ltout(),
            .carryin(n19312),
            .carryout(n19313),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__33923),
            .sr(N__33894));
    defparam acadc_skipcnt_i0_i3_LC_13_17_2.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i3_LC_13_17_2.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i3_LC_13_17_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i3_LC_13_17_2 (
            .in0(_gnd_net_),
            .in1(N__33654),
            .in2(_gnd_net_),
            .in3(N__33637),
            .lcout(acadc_skipcnt_3),
            .ltout(),
            .carryin(n19313),
            .carryout(n19314),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__33923),
            .sr(N__33894));
    defparam acadc_skipcnt_i0_i4_LC_13_17_3.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i4_LC_13_17_3.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i4_LC_13_17_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i4_LC_13_17_3 (
            .in0(_gnd_net_),
            .in1(N__33630),
            .in2(_gnd_net_),
            .in3(N__33613),
            .lcout(acadc_skipcnt_4),
            .ltout(),
            .carryin(n19314),
            .carryout(n19315),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__33923),
            .sr(N__33894));
    defparam acadc_skipcnt_i0_i5_LC_13_17_4.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i5_LC_13_17_4.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i5_LC_13_17_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i5_LC_13_17_4 (
            .in0(_gnd_net_),
            .in1(N__33606),
            .in2(_gnd_net_),
            .in3(N__33592),
            .lcout(acadc_skipcnt_5),
            .ltout(),
            .carryin(n19315),
            .carryout(n19316),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__33923),
            .sr(N__33894));
    defparam acadc_skipcnt_i0_i6_LC_13_17_5.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i6_LC_13_17_5.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i6_LC_13_17_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i6_LC_13_17_5 (
            .in0(_gnd_net_),
            .in1(N__33753),
            .in2(_gnd_net_),
            .in3(N__33739),
            .lcout(acadc_skipcnt_6),
            .ltout(),
            .carryin(n19316),
            .carryout(n19317),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__33923),
            .sr(N__33894));
    defparam acadc_skipcnt_i0_i7_LC_13_17_6.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i7_LC_13_17_6.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i7_LC_13_17_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i7_LC_13_17_6 (
            .in0(_gnd_net_),
            .in1(N__36318),
            .in2(_gnd_net_),
            .in3(N__33736),
            .lcout(acadc_skipcnt_7),
            .ltout(),
            .carryin(n19317),
            .carryout(n19318),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__33923),
            .sr(N__33894));
    defparam acadc_skipcnt_i0_i8_LC_13_17_7.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i8_LC_13_17_7.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i8_LC_13_17_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i8_LC_13_17_7 (
            .in0(_gnd_net_),
            .in1(N__33729),
            .in2(_gnd_net_),
            .in3(N__33715),
            .lcout(acadc_skipcnt_8),
            .ltout(),
            .carryin(n19318),
            .carryout(n19319),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__33923),
            .sr(N__33894));
    defparam acadc_skipcnt_i0_i9_LC_13_18_0.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i9_LC_13_18_0.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i9_LC_13_18_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i9_LC_13_18_0 (
            .in0(_gnd_net_),
            .in1(N__36627),
            .in2(_gnd_net_),
            .in3(N__33712),
            .lcout(acadc_skipcnt_9),
            .ltout(),
            .carryin(bfn_13_18_0_),
            .carryout(n19320),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__33937),
            .sr(N__33898));
    defparam acadc_skipcnt_i0_i10_LC_13_18_1.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i10_LC_13_18_1.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i10_LC_13_18_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i10_LC_13_18_1 (
            .in0(_gnd_net_),
            .in1(N__38790),
            .in2(_gnd_net_),
            .in3(N__33709),
            .lcout(acadc_skipcnt_10),
            .ltout(),
            .carryin(n19320),
            .carryout(n19321),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__33937),
            .sr(N__33898));
    defparam acadc_skipcnt_i0_i11_LC_13_18_2.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i11_LC_13_18_2.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i11_LC_13_18_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i11_LC_13_18_2 (
            .in0(_gnd_net_),
            .in1(N__36411),
            .in2(_gnd_net_),
            .in3(N__33706),
            .lcout(acadc_skipcnt_11),
            .ltout(),
            .carryin(n19321),
            .carryout(n19322),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__33937),
            .sr(N__33898));
    defparam acadc_skipcnt_i0_i12_LC_13_18_3.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i12_LC_13_18_3.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i12_LC_13_18_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i12_LC_13_18_3 (
            .in0(_gnd_net_),
            .in1(N__38808),
            .in2(_gnd_net_),
            .in3(N__33703),
            .lcout(acadc_skipcnt_12),
            .ltout(),
            .carryin(n19322),
            .carryout(n19323),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__33937),
            .sr(N__33898));
    defparam acadc_skipcnt_i0_i13_LC_13_18_4.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i13_LC_13_18_4.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i13_LC_13_18_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i13_LC_13_18_4 (
            .in0(_gnd_net_),
            .in1(N__33696),
            .in2(_gnd_net_),
            .in3(N__33682),
            .lcout(acadc_skipcnt_13),
            .ltout(),
            .carryin(n19323),
            .carryout(n19324),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__33937),
            .sr(N__33898));
    defparam acadc_skipcnt_i0_i14_LC_13_18_5.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i14_LC_13_18_5.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i14_LC_13_18_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i14_LC_13_18_5 (
            .in0(_gnd_net_),
            .in1(N__36426),
            .in2(_gnd_net_),
            .in3(N__33679),
            .lcout(acadc_skipcnt_14),
            .ltout(),
            .carryin(n19324),
            .carryout(n19325),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__33937),
            .sr(N__33898));
    defparam acadc_skipcnt_i0_i15_LC_13_18_6.C_ON=1'b0;
    defparam acadc_skipcnt_i0_i15_LC_13_18_6.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i15_LC_13_18_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i15_LC_13_18_6 (
            .in0(_gnd_net_),
            .in1(N__36612),
            .in2(_gnd_net_),
            .in3(N__33940),
            .lcout(acadc_skipcnt_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__33937),
            .sr(N__33898));
    defparam \SIG_DDS.tmp_buf_i12_LC_13_19_1 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i12_LC_13_19_1 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i12_LC_13_19_1 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \SIG_DDS.tmp_buf_i12_LC_13_19_1  (
            .in0(N__55878),
            .in1(N__55660),
            .in2(N__33877),
            .in3(N__33868),
            .lcout(\SIG_DDS.tmp_buf_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55196),
            .ce(N__40315),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i2_LC_13_19_3 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i2_LC_13_19_3 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i2_LC_13_19_3 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \SIG_DDS.tmp_buf_i2_LC_13_19_3  (
            .in0(N__55879),
            .in1(N__55661),
            .in2(N__33829),
            .in3(N__42754),
            .lcout(\SIG_DDS.tmp_buf_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55196),
            .ce(N__40315),
            .sr(_gnd_net_));
    defparam \comm_spi.data_rx_i0_12197_12198_reset_LC_14_3_0 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i0_12197_12198_reset_LC_14_3_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i0_12197_12198_reset_LC_14_3_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.data_rx_i0_12197_12198_reset_LC_14_3_0  (
            .in0(N__37425),
            .in1(N__34996),
            .in2(_gnd_net_),
            .in3(N__33819),
            .lcout(\comm_spi.n14600 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52441),
            .ce(),
            .sr(N__33796));
    defparam \ADC_VDC.genclk.i18725_4_lut_LC_14_4_0 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i18725_4_lut_LC_14_4_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i18725_4_lut_LC_14_4_0 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \ADC_VDC.genclk.i18725_4_lut_LC_14_4_0  (
            .in0(N__37017),
            .in1(N__37110),
            .in2(N__37063),
            .in3(N__37125),
            .lcout(),
            .ltout(\ADC_VDC.genclk.n21172_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i18906_4_lut_LC_14_4_1 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i18906_4_lut_LC_14_4_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i18906_4_lut_LC_14_4_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i18906_4_lut_LC_14_4_1  (
            .in0(N__33769),
            .in1(N__33760),
            .in2(N__33784),
            .in3(N__35002),
            .lcout(\ADC_VDC.genclk.n21166 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i12_4_lut_adj_27_LC_14_4_2 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i12_4_lut_adj_27_LC_14_4_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i12_4_lut_adj_27_LC_14_4_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i12_4_lut_adj_27_LC_14_4_2  (
            .in0(N__37170),
            .in1(N__37251),
            .in2(N__37498),
            .in3(N__37218),
            .lcout(\ADC_VDC.genclk.n28_adj_1400 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i10_4_lut_adj_28_LC_14_4_3 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i10_4_lut_adj_28_LC_14_4_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i10_4_lut_adj_28_LC_14_4_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i10_4_lut_adj_28_LC_14_4_3  (
            .in0(N__37077),
            .in1(N__37185),
            .in2(N__37039),
            .in3(N__37269),
            .lcout(\ADC_VDC.genclk.n26_adj_1401 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i11_4_lut_adj_29_LC_14_4_4 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i11_4_lut_adj_29_LC_14_4_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i11_4_lut_adj_29_LC_14_4_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i11_4_lut_adj_29_LC_14_4_4  (
            .in0(N__37203),
            .in1(N__37092),
            .in2(N__37288),
            .in3(N__37236),
            .lcout(\ADC_VDC.genclk.n27_adj_1402 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.imosi_44_12183_12184_reset_LC_14_5_0 .C_ON=1'b0;
    defparam \comm_spi.imosi_44_12183_12184_reset_LC_14_5_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.imosi_44_12183_12184_reset_LC_14_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \comm_spi.imosi_44_12183_12184_reset_LC_14_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37342),
            .lcout(\comm_spi.n14586 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55074),
            .ce(),
            .sr(N__37300));
    defparam \ADC_VDC.genclk.div_state_i1_LC_14_6_1 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.div_state_i1_LC_14_6_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.div_state_i1_LC_14_6_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ADC_VDC.genclk.div_state_i1_LC_14_6_1  (
            .in0(_gnd_net_),
            .in1(N__34974),
            .in2(_gnd_net_),
            .in3(N__34918),
            .lcout(\ADC_VDC.genclk.div_state_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVADC_VDC.genclk.div_state_i1C_net ),
            .ce(N__34885),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_2_lut_LC_14_6_4 .C_ON=1'b0;
    defparam \ADC_VDC.i1_2_lut_LC_14_6_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_2_lut_LC_14_6_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \ADC_VDC.i1_2_lut_LC_14_6_4  (
            .in0(N__34872),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34747),
            .lcout(\ADC_VDC.n62 ),
            .ltout(\ADC_VDC.n62_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i16006_4_lut_LC_14_6_5 .C_ON=1'b0;
    defparam \ADC_VDC.i16006_4_lut_LC_14_6_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i16006_4_lut_LC_14_6_5 .LUT_INIT=16'b1001100010111010;
    LogicCell40 \ADC_VDC.i16006_4_lut_LC_14_6_5  (
            .in0(N__34566),
            .in1(N__34375),
            .in2(N__34162),
            .in3(N__34155),
            .lcout(\ADC_VDC.n11736 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_137_Mux_7_i2_3_lut_LC_14_7_0.C_ON=1'b0;
    defparam mux_137_Mux_7_i2_3_lut_LC_14_7_0.SEQ_MODE=4'b0000;
    defparam mux_137_Mux_7_i2_3_lut_LC_14_7_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_137_Mux_7_i2_3_lut_LC_14_7_0 (
            .in0(N__34003),
            .in1(N__35230),
            .in2(_gnd_net_),
            .in3(N__51622),
            .lcout(),
            .ltout(n2_adj_1559_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i7_LC_14_7_1.C_ON=1'b0;
    defparam comm_tx_buf_i7_LC_14_7_1.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i7_LC_14_7_1.LUT_INIT=16'b1111101001000100;
    LogicCell40 comm_tx_buf_i7_LC_14_7_1 (
            .in0(N__50101),
            .in1(N__33988),
            .in2(N__33979),
            .in3(N__35044),
            .lcout(comm_tx_buf_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55077),
            .ce(N__47124),
            .sr(N__47056));
    defparam mux_137_Mux_7_i4_3_lut_LC_14_7_2.C_ON=1'b0;
    defparam mux_137_Mux_7_i4_3_lut_LC_14_7_2.SEQ_MODE=4'b0000;
    defparam mux_137_Mux_7_i4_3_lut_LC_14_7_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_137_Mux_7_i4_3_lut_LC_14_7_2 (
            .in0(N__35110),
            .in1(N__33976),
            .in2(_gnd_net_),
            .in3(N__51620),
            .lcout(n4_adj_1560),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19043_2_lut_LC_14_7_3.C_ON=1'b0;
    defparam i19043_2_lut_LC_14_7_3.SEQ_MODE=4'b0000;
    defparam i19043_2_lut_LC_14_7_3.LUT_INIT=16'b0101010100000000;
    LogicCell40 i19043_2_lut_LC_14_7_3 (
            .in0(N__51621),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33964),
            .lcout(),
            .ltout(n21276_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_1__bdd_4_lut_LC_14_7_4.C_ON=1'b0;
    defparam comm_index_1__bdd_4_lut_LC_14_7_4.SEQ_MODE=4'b0000;
    defparam comm_index_1__bdd_4_lut_LC_14_7_4.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_index_1__bdd_4_lut_LC_14_7_4 (
            .in0(N__35053),
            .in1(N__49529),
            .in2(N__35047),
            .in3(N__50100),
            .lcout(n22105),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i19164_4_lut_3_lut_LC_14_7_6 .C_ON=1'b0;
    defparam \comm_spi.i19164_4_lut_3_lut_LC_14_7_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19164_4_lut_3_lut_LC_14_7_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \comm_spi.i19164_4_lut_3_lut_LC_14_7_6  (
            .in0(N__44271),
            .in1(N__37391),
            .in2(_gnd_net_),
            .in3(N__55409),
            .lcout(\comm_spi.n14588 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_100_2_lut_LC_14_7_7 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_100_2_lut_LC_14_7_7 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_100_2_lut_LC_14_7_7 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \comm_spi.RESET_I_0_100_2_lut_LC_14_7_7  (
            .in0(N__55408),
            .in1(_gnd_net_),
            .in2(N__37396),
            .in3(_gnd_net_),
            .lcout(\comm_spi.data_tx_7__N_766 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_0__bdd_4_lut_19379_LC_14_8_0.C_ON=1'b0;
    defparam comm_index_0__bdd_4_lut_19379_LC_14_8_0.SEQ_MODE=4'b0000;
    defparam comm_index_0__bdd_4_lut_19379_LC_14_8_0.LUT_INIT=16'b1110101001001010;
    LogicCell40 comm_index_0__bdd_4_lut_19379_LC_14_8_0 (
            .in0(N__51638),
            .in1(N__35173),
            .in2(N__49543),
            .in3(N__35038),
            .lcout(),
            .ltout(n21985_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n21985_bdd_4_lut_LC_14_8_1.C_ON=1'b0;
    defparam n21985_bdd_4_lut_LC_14_8_1.SEQ_MODE=4'b0000;
    defparam n21985_bdd_4_lut_LC_14_8_1.LUT_INIT=16'b1111010010100100;
    LogicCell40 n21985_bdd_4_lut_LC_14_8_1 (
            .in0(N__49536),
            .in1(N__38712),
            .in2(N__35026),
            .in3(N__42815),
            .lcout(),
            .ltout(n21988_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i2_LC_14_8_2.C_ON=1'b0;
    defparam comm_tx_buf_i2_LC_14_8_2.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i2_LC_14_8_2.LUT_INIT=16'b1111101001010000;
    LogicCell40 comm_tx_buf_i2_LC_14_8_2 (
            .in0(N__50077),
            .in1(_gnd_net_),
            .in2(N__35023),
            .in3(N__35059),
            .lcout(comm_tx_buf_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55085),
            .ce(N__47136),
            .sr(N__47057));
    defparam i14920_3_lut_LC_14_8_3.C_ON=1'b0;
    defparam i14920_3_lut_LC_14_8_3.SEQ_MODE=4'b0000;
    defparam i14920_3_lut_LC_14_8_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 i14920_3_lut_LC_14_8_3 (
            .in0(N__35131),
            .in1(N__41354),
            .in2(_gnd_net_),
            .in3(N__50075),
            .lcout(),
            .ltout(n17304_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18311_4_lut_LC_14_8_4.C_ON=1'b0;
    defparam i18311_4_lut_LC_14_8_4.SEQ_MODE=4'b0000;
    defparam i18311_4_lut_LC_14_8_4.LUT_INIT=16'b0100010011110000;
    LogicCell40 i18311_4_lut_LC_14_8_4 (
            .in0(N__50076),
            .in1(N__35020),
            .in2(N__35008),
            .in3(N__49537),
            .lcout(),
            .ltout(n20906_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i0_LC_14_8_5.C_ON=1'b0;
    defparam comm_tx_buf_i0_LC_14_8_5.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i0_LC_14_8_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 comm_tx_buf_i0_LC_14_8_5 (
            .in0(_gnd_net_),
            .in1(N__38113),
            .in2(N__35005),
            .in3(N__51641),
            .lcout(comm_tx_buf_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55085),
            .ce(N__47136),
            .sr(N__47057));
    defparam mux_137_Mux_2_i4_3_lut_LC_14_8_6.C_ON=1'b0;
    defparam mux_137_Mux_2_i4_3_lut_LC_14_8_6.SEQ_MODE=4'b0000;
    defparam mux_137_Mux_2_i4_3_lut_LC_14_8_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_137_Mux_2_i4_3_lut_LC_14_8_6 (
            .in0(N__51639),
            .in1(N__35356),
            .in2(_gnd_net_),
            .in3(N__35098),
            .lcout(),
            .ltout(n4_adj_1568_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18191_4_lut_LC_14_8_7.C_ON=1'b0;
    defparam i18191_4_lut_LC_14_8_7.SEQ_MODE=4'b0000;
    defparam i18191_4_lut_LC_14_8_7.LUT_INIT=16'b0101000011011000;
    LogicCell40 i18191_4_lut_LC_14_8_7 (
            .in0(N__49535),
            .in1(N__35086),
            .in2(N__35062),
            .in3(N__51640),
            .lcout(n20786),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_rx_i7_LC_14_9_0 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i7_LC_14_9_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i7_LC_14_9_0 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \comm_spi.data_rx_i7_LC_14_9_0  (
            .in0(N__46376),
            .in1(N__35757),
            .in2(_gnd_net_),
            .in3(N__46332),
            .lcout(comm_rx_buf_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52443),
            .ce(),
            .sr(N__55431));
    defparam \comm_spi.data_rx_i6_LC_14_9_1 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i6_LC_14_9_1 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i6_LC_14_9_1 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \comm_spi.data_rx_i6_LC_14_9_1  (
            .in0(N__46331),
            .in1(N__37953),
            .in2(_gnd_net_),
            .in3(N__46375),
            .lcout(comm_rx_buf_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52443),
            .ce(),
            .sr(N__55431));
    defparam \comm_spi.data_rx_i5_LC_14_9_2 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i5_LC_14_9_2 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i5_LC_14_9_2 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \comm_spi.data_rx_i5_LC_14_9_2  (
            .in0(N__46374),
            .in1(N__35617),
            .in2(_gnd_net_),
            .in3(N__46330),
            .lcout(comm_rx_buf_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52443),
            .ce(),
            .sr(N__55431));
    defparam \comm_spi.data_rx_i4_LC_14_9_3 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i4_LC_14_9_3 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i4_LC_14_9_3 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \comm_spi.data_rx_i4_LC_14_9_3  (
            .in0(N__46329),
            .in1(N__35509),
            .in2(_gnd_net_),
            .in3(N__46373),
            .lcout(comm_rx_buf_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52443),
            .ce(),
            .sr(N__55431));
    defparam \comm_spi.data_rx_i3_LC_14_9_4 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i3_LC_14_9_4 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i3_LC_14_9_4 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \comm_spi.data_rx_i3_LC_14_9_4  (
            .in0(N__46372),
            .in1(N__35401),
            .in2(_gnd_net_),
            .in3(N__46328),
            .lcout(comm_rx_buf_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52443),
            .ce(),
            .sr(N__55431));
    defparam \comm_spi.data_rx_i2_LC_14_9_5 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i2_LC_14_9_5 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i2_LC_14_9_5 .LUT_INIT=16'b1100110010001000;
    LogicCell40 \comm_spi.data_rx_i2_LC_14_9_5  (
            .in0(N__46327),
            .in1(N__35933),
            .in2(_gnd_net_),
            .in3(N__46371),
            .lcout(comm_rx_buf_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52443),
            .ce(),
            .sr(N__55431));
    defparam \comm_spi.data_rx_i1_LC_14_9_6 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i1_LC_14_9_6 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i1_LC_14_9_6 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \comm_spi.data_rx_i1_LC_14_9_6  (
            .in0(N__46370),
            .in1(N__46326),
            .in2(_gnd_net_),
            .in3(N__36241),
            .lcout(comm_rx_buf_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52443),
            .ce(),
            .sr(N__55431));
    defparam comm_buf_2__i0_LC_14_10_0.C_ON=1'b0;
    defparam comm_buf_2__i0_LC_14_10_0.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i0_LC_14_10_0.LUT_INIT=16'b1110111000100010;
    LogicCell40 comm_buf_2__i0_LC_14_10_0 (
            .in0(N__35239),
            .in1(N__53938),
            .in2(_gnd_net_),
            .in3(N__36233),
            .lcout(comm_buf_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55099),
            .ce(N__37921),
            .sr(N__38350));
    defparam comm_buf_2__i7_LC_14_10_1.C_ON=1'b0;
    defparam comm_buf_2__i7_LC_14_10_1.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i7_LC_14_10_1.LUT_INIT=16'b1111010110100000;
    LogicCell40 comm_buf_2__i7_LC_14_10_1 (
            .in0(N__53937),
            .in1(_gnd_net_),
            .in2(N__36858),
            .in3(N__47428),
            .lcout(comm_buf_2_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55099),
            .ce(N__37921),
            .sr(N__38350));
    defparam comm_buf_2__i6_LC_14_10_2.C_ON=1'b0;
    defparam comm_buf_2__i6_LC_14_10_2.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i6_LC_14_10_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_2__i6_LC_14_10_2 (
            .in0(N__35758),
            .in1(N__35221),
            .in2(_gnd_net_),
            .in3(N__53941),
            .lcout(comm_buf_2_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55099),
            .ce(N__37921),
            .sr(N__38350));
    defparam comm_buf_2__i4_LC_14_10_3.C_ON=1'b0;
    defparam comm_buf_2__i4_LC_14_10_3.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i4_LC_14_10_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_2__i4_LC_14_10_3 (
            .in0(N__53936),
            .in1(N__35618),
            .in2(_gnd_net_),
            .in3(N__56053),
            .lcout(comm_buf_2_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55099),
            .ce(N__37921),
            .sr(N__38350));
    defparam comm_buf_2__i3_LC_14_10_4.C_ON=1'b0;
    defparam comm_buf_2__i3_LC_14_10_4.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i3_LC_14_10_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_2__i3_LC_14_10_4 (
            .in0(N__35510),
            .in1(N__35203),
            .in2(_gnd_net_),
            .in3(N__53940),
            .lcout(comm_buf_2_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55099),
            .ce(N__37921),
            .sr(N__38350));
    defparam comm_buf_2__i2_LC_14_10_5.C_ON=1'b0;
    defparam comm_buf_2__i2_LC_14_10_5.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i2_LC_14_10_5.LUT_INIT=16'b1111010110100000;
    LogicCell40 comm_buf_2__i2_LC_14_10_5 (
            .in0(N__53935),
            .in1(_gnd_net_),
            .in2(N__35420),
            .in3(N__35185),
            .lcout(comm_buf_2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55099),
            .ce(N__37921),
            .sr(N__38350));
    defparam comm_buf_2__i1_LC_14_10_6.C_ON=1'b0;
    defparam comm_buf_2__i1_LC_14_10_6.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i1_LC_14_10_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_2__i1_LC_14_10_6 (
            .in0(N__35934),
            .in1(N__35164),
            .in2(_gnd_net_),
            .in3(N__53939),
            .lcout(comm_buf_2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55099),
            .ce(N__37921),
            .sr(N__38350));
    defparam comm_buf_5__i0_LC_14_11_0.C_ON=1'b0;
    defparam comm_buf_5__i0_LC_14_11_0.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i0_LC_14_11_0.LUT_INIT=16'b1110111000100010;
    LogicCell40 comm_buf_5__i0_LC_14_11_0 (
            .in0(N__35143),
            .in1(N__53946),
            .in2(_gnd_net_),
            .in3(N__36237),
            .lcout(comm_buf_5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55108),
            .ce(N__38104),
            .sr(N__38092));
    defparam comm_buf_5__i7_LC_14_11_1.C_ON=1'b0;
    defparam comm_buf_5__i7_LC_14_11_1.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i7_LC_14_11_1.LUT_INIT=16'b1111010110100000;
    LogicCell40 comm_buf_5__i7_LC_14_11_1 (
            .in0(N__53945),
            .in1(_gnd_net_),
            .in2(N__36880),
            .in3(N__35119),
            .lcout(comm_buf_5_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55108),
            .ce(N__38104),
            .sr(N__38092));
    defparam comm_buf_5__i6_LC_14_11_2.C_ON=1'b0;
    defparam comm_buf_5__i6_LC_14_11_2.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i6_LC_14_11_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_5__i6_LC_14_11_2 (
            .in0(N__35779),
            .in1(N__35716),
            .in2(_gnd_net_),
            .in3(N__53949),
            .lcout(comm_buf_5_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55108),
            .ce(N__38104),
            .sr(N__38092));
    defparam comm_buf_5__i5_LC_14_11_3.C_ON=1'b0;
    defparam comm_buf_5__i5_LC_14_11_3.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i5_LC_14_11_3.LUT_INIT=16'b1111010110100000;
    LogicCell40 comm_buf_5__i5_LC_14_11_3 (
            .in0(N__53944),
            .in1(_gnd_net_),
            .in2(N__37994),
            .in3(N__35689),
            .lcout(comm_buf_5_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55108),
            .ce(N__38104),
            .sr(N__38092));
    defparam comm_buf_5__i4_LC_14_11_4.C_ON=1'b0;
    defparam comm_buf_5__i4_LC_14_11_4.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i4_LC_14_11_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_5__i4_LC_14_11_4 (
            .in0(N__35636),
            .in1(N__35584),
            .in2(_gnd_net_),
            .in3(N__53948),
            .lcout(comm_buf_5_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55108),
            .ce(N__38104),
            .sr(N__38092));
    defparam comm_buf_5__i3_LC_14_11_5.C_ON=1'b0;
    defparam comm_buf_5__i3_LC_14_11_5.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i3_LC_14_11_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_5__i3_LC_14_11_5 (
            .in0(N__53943),
            .in1(N__35530),
            .in2(_gnd_net_),
            .in3(N__35482),
            .lcout(comm_buf_5_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55108),
            .ce(N__38104),
            .sr(N__38092));
    defparam comm_buf_5__i2_LC_14_11_6.C_ON=1'b0;
    defparam comm_buf_5__i2_LC_14_11_6.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i2_LC_14_11_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_5__i2_LC_14_11_6 (
            .in0(N__35421),
            .in1(N__35368),
            .in2(_gnd_net_),
            .in3(N__53947),
            .lcout(comm_buf_5_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55108),
            .ce(N__38104),
            .sr(N__38092));
    defparam comm_buf_5__i1_LC_14_11_7.C_ON=1'b0;
    defparam comm_buf_5__i1_LC_14_11_7.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i1_LC_14_11_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_5__i1_LC_14_11_7 (
            .in0(N__53942),
            .in1(N__35951),
            .in2(_gnd_net_),
            .in3(N__35347),
            .lcout(comm_buf_5_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55108),
            .ce(N__38104),
            .sr(N__38092));
    defparam i18242_3_lut_LC_14_12_0.C_ON=1'b0;
    defparam i18242_3_lut_LC_14_12_0.SEQ_MODE=4'b0000;
    defparam i18242_3_lut_LC_14_12_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 i18242_3_lut_LC_14_12_0 (
            .in0(N__57552),
            .in1(N__35335),
            .in2(_gnd_net_),
            .in3(N__35245),
            .lcout(n20837),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_1_i19_3_lut_LC_14_12_1.C_ON=1'b0;
    defparam mux_129_Mux_1_i19_3_lut_LC_14_12_1.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_1_i19_3_lut_LC_14_12_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_129_Mux_1_i19_3_lut_LC_14_12_1 (
            .in0(N__56950),
            .in1(N__35308),
            .in2(_gnd_net_),
            .in3(N__35283),
            .lcout(n19_adj_1508),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_2__bdd_4_lut_19457_LC_14_12_2.C_ON=1'b0;
    defparam comm_cmd_2__bdd_4_lut_19457_LC_14_12_2.SEQ_MODE=4'b0000;
    defparam comm_cmd_2__bdd_4_lut_19457_LC_14_12_2.LUT_INIT=16'b1110101001100010;
    LogicCell40 comm_cmd_2__bdd_4_lut_19457_LC_14_12_2 (
            .in0(N__47847),
            .in1(N__56264),
            .in2(N__36079),
            .in3(N__36001),
            .lcout(),
            .ltout(n22069_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22069_bdd_4_lut_LC_14_12_3.C_ON=1'b0;
    defparam n22069_bdd_4_lut_LC_14_12_3.SEQ_MODE=4'b0000;
    defparam n22069_bdd_4_lut_LC_14_12_3.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22069_bdd_4_lut_LC_14_12_3 (
            .in0(N__56265),
            .in1(N__36067),
            .in2(N__36049),
            .in3(N__36046),
            .lcout(n22072),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_1_i26_3_lut_LC_14_12_4.C_ON=1'b0;
    defparam mux_129_Mux_1_i26_3_lut_LC_14_12_4.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_1_i26_3_lut_LC_14_12_4.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_129_Mux_1_i26_3_lut_LC_14_12_4 (
            .in0(N__36040),
            .in1(N__56949),
            .in2(_gnd_net_),
            .in3(N__46908),
            .lcout(),
            .ltout(n26_adj_1509_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18230_4_lut_LC_14_12_5.C_ON=1'b0;
    defparam i18230_4_lut_LC_14_12_5.SEQ_MODE=4'b0000;
    defparam i18230_4_lut_LC_14_12_5.LUT_INIT=16'b0111010000110000;
    LogicCell40 i18230_4_lut_LC_14_12_5 (
            .in0(N__56951),
            .in1(N__57551),
            .in2(N__36025),
            .in3(N__36022),
            .lcout(n20825),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i1_LC_14_12_6.C_ON=1'b0;
    defparam comm_buf_1__i1_LC_14_12_6.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i1_LC_14_12_6.LUT_INIT=16'b1011101110001000;
    LogicCell40 comm_buf_1__i1_LC_14_12_6 (
            .in0(N__35971),
            .in1(N__54031),
            .in2(_gnd_net_),
            .in3(N__35905),
            .lcout(comm_buf_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55119),
            .ce(N__38523),
            .sr(N__36780));
    defparam mux_129_Mux_0_i26_3_lut_LC_14_13_1.C_ON=1'b0;
    defparam mux_129_Mux_0_i26_3_lut_LC_14_13_1.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_0_i26_3_lut_LC_14_13_1.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_129_Mux_0_i26_3_lut_LC_14_13_1 (
            .in0(N__35899),
            .in1(N__56831),
            .in2(_gnd_net_),
            .in3(N__46935),
            .lcout(),
            .ltout(n26_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19452_LC_14_13_2.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19452_LC_14_13_2.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19452_LC_14_13_2.LUT_INIT=16'b1011100011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_19452_LC_14_13_2 (
            .in0(N__35881),
            .in1(N__57479),
            .in2(N__35863),
            .in3(N__47726),
            .lcout(),
            .ltout(n22021_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22021_bdd_4_lut_LC_14_13_3.C_ON=1'b0;
    defparam n22021_bdd_4_lut_LC_14_13_3.SEQ_MODE=4'b0000;
    defparam n22021_bdd_4_lut_LC_14_13_3.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22021_bdd_4_lut_LC_14_13_3 (
            .in0(N__47727),
            .in1(N__35860),
            .in2(N__35833),
            .in3(N__41752),
            .lcout(n22024),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1541068_i1_3_lut_LC_14_13_5.C_ON=1'b0;
    defparam i1541068_i1_3_lut_LC_14_13_5.SEQ_MODE=4'b0000;
    defparam i1541068_i1_3_lut_LC_14_13_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 i1541068_i1_3_lut_LC_14_13_5 (
            .in0(N__35830),
            .in1(N__35824),
            .in2(_gnd_net_),
            .in3(N__56269),
            .lcout(),
            .ltout(n30_adj_1478_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i0_LC_14_13_6.C_ON=1'b0;
    defparam comm_buf_1__i0_LC_14_13_6.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i0_LC_14_13_6.LUT_INIT=16'b1111110000110000;
    LogicCell40 comm_buf_1__i0_LC_14_13_6 (
            .in0(_gnd_net_),
            .in1(N__54032),
            .in2(N__36262),
            .in3(N__36253),
            .lcout(comm_buf_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55128),
            .ce(N__38533),
            .sr(N__36795));
    defparam \ADC_VAC.ADC_DATA_i5_LC_14_14_0 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i5_LC_14_14_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i5_LC_14_14_0 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC.ADC_DATA_i5_LC_14_14_0  (
            .in0(N__48526),
            .in1(N__48350),
            .in2(N__38304),
            .in3(N__36165),
            .lcout(buf_adcdata_vac_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55140),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i13_LC_14_14_1 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i13_LC_14_14_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i13_LC_14_14_1 .LUT_INIT=16'b1011100000110000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i13_LC_14_14_1  (
            .in0(N__48349),
            .in1(N__37884),
            .in2(N__36166),
            .in3(N__47967),
            .lcout(cmd_rdadctmp_13_adj_1430),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55140),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i14_LC_14_14_2 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i14_LC_14_14_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i14_LC_14_14_2 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i14_LC_14_14_2  (
            .in0(N__37885),
            .in1(N__36164),
            .in2(N__38759),
            .in3(N__48351),
            .lcout(cmd_rdadctmp_14_adj_1429),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55140),
            .ce(),
            .sr(_gnd_net_));
    defparam i12345_2_lut_LC_14_14_3.C_ON=1'b0;
    defparam i12345_2_lut_LC_14_14_3.SEQ_MODE=4'b0000;
    defparam i12345_2_lut_LC_14_14_3.LUT_INIT=16'b1100110000000000;
    LogicCell40 i12345_2_lut_LC_14_14_3 (
            .in0(_gnd_net_),
            .in1(N__54600),
            .in2(_gnd_net_),
            .in3(N__38497),
            .lcout(n14742),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i6_LC_14_14_4.C_ON=1'b0;
    defparam buf_dds1_i6_LC_14_14_4.SEQ_MODE=4'b1000;
    defparam buf_dds1_i6_LC_14_14_4.LUT_INIT=16'b1110001000000000;
    LogicCell40 buf_dds1_i6_LC_14_14_4 (
            .in0(N__36108),
            .in1(N__45876),
            .in2(N__51430),
            .in3(N__45987),
            .lcout(buf_dds1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55140),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_4_i16_3_lut_LC_14_14_5.C_ON=1'b0;
    defparam mux_129_Mux_4_i16_3_lut_LC_14_14_5.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_4_i16_3_lut_LC_14_14_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_129_Mux_4_i16_3_lut_LC_14_14_5 (
            .in0(N__36151),
            .in1(N__42711),
            .in2(_gnd_net_),
            .in3(N__56983),
            .lcout(n16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_6_i16_3_lut_LC_14_14_6.C_ON=1'b0;
    defparam mux_129_Mux_6_i16_3_lut_LC_14_14_6.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_6_i16_3_lut_LC_14_14_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_129_Mux_6_i16_3_lut_LC_14_14_6 (
            .in0(N__56984),
            .in1(N__36104),
            .in2(_gnd_net_),
            .in3(N__42654),
            .lcout(n16_adj_1488),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18229_3_lut_LC_14_14_7.C_ON=1'b0;
    defparam i18229_3_lut_LC_14_14_7.SEQ_MODE=4'b0000;
    defparam i18229_3_lut_LC_14_14_7.LUT_INIT=16'b1110111001000100;
    LogicCell40 i18229_3_lut_LC_14_14_7 (
            .in0(N__57525),
            .in1(N__36564),
            .in2(_gnd_net_),
            .in3(N__38374),
            .lcout(n20824),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_354_Mux_2_i15_4_lut_LC_14_15_0.C_ON=1'b0;
    defparam comm_state_3__I_0_354_Mux_2_i15_4_lut_LC_14_15_0.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_354_Mux_2_i15_4_lut_LC_14_15_0.LUT_INIT=16'b0011101100001000;
    LogicCell40 comm_state_3__I_0_354_Mux_2_i15_4_lut_LC_14_15_0 (
            .in0(N__36636),
            .in1(N__54670),
            .in2(N__51984),
            .in3(N__41841),
            .lcout(data_index_9_N_212_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7_4_lut_LC_14_15_1.C_ON=1'b0;
    defparam i7_4_lut_LC_14_15_1.SEQ_MODE=4'b0000;
    defparam i7_4_lut_LC_14_15_1.LUT_INIT=16'b0111110110111110;
    LogicCell40 i7_4_lut_LC_14_15_1 (
            .in0(N__36430),
            .in1(N__36412),
            .in2(N__45477),
            .in3(N__36653),
            .lcout(n23_adj_1586),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6412_3_lut_LC_14_15_2.C_ON=1'b0;
    defparam i6412_3_lut_LC_14_15_2.SEQ_MODE=4'b0000;
    defparam i6412_3_lut_LC_14_15_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 i6412_3_lut_LC_14_15_2 (
            .in0(N__41827),
            .in1(N__36378),
            .in2(_gnd_net_),
            .in3(N__43273),
            .lcout(n8_adj_1543),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i2_LC_14_15_3.C_ON=1'b0;
    defparam acadc_skipCount_i2_LC_14_15_3.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i2_LC_14_15_3.LUT_INIT=16'b0111001101000000;
    LogicCell40 acadc_skipCount_i2_LC_14_15_3 (
            .in0(N__51893),
            .in1(N__39313),
            .in2(N__42808),
            .in3(N__36302),
            .lcout(acadc_skipCount_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55153),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i2_LC_14_15_4.C_ON=1'b0;
    defparam data_index_i2_LC_14_15_4.SEQ_MODE=4'b1000;
    defparam data_index_i2_LC_14_15_4.LUT_INIT=16'b0011101100001000;
    LogicCell40 data_index_i2_LC_14_15_4 (
            .in0(N__36637),
            .in1(N__54671),
            .in2(N__51985),
            .in3(N__41842),
            .lcout(data_index_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55153),
            .ce(),
            .sr(_gnd_net_));
    defparam i6_4_lut_LC_14_15_5.C_ON=1'b0;
    defparam i6_4_lut_LC_14_15_5.SEQ_MODE=4'b0000;
    defparam i6_4_lut_LC_14_15_5.LUT_INIT=16'b0111101111011110;
    LogicCell40 i6_4_lut_LC_14_15_5 (
            .in0(N__36334),
            .in1(N__36319),
            .in2(N__36303),
            .in3(N__36977),
            .lcout(),
            .ltout(n22_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i14_4_lut_LC_14_15_6.C_ON=1'b0;
    defparam i14_4_lut_LC_14_15_6.SEQ_MODE=4'b0000;
    defparam i14_4_lut_LC_14_15_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i14_4_lut_LC_14_15_6 (
            .in0(N__36280),
            .in1(N__38776),
            .in2(N__36274),
            .in3(N__36574),
            .lcout(n30_adj_1571),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i7_LC_14_15_7.C_ON=1'b0;
    defparam acadc_skipCount_i7_LC_14_15_7.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i7_LC_14_15_7.LUT_INIT=16'b0111001101000000;
    LogicCell40 acadc_skipCount_i7_LC_14_15_7 (
            .in0(N__51894),
            .in1(N__39314),
            .in2(N__42619),
            .in3(N__36978),
            .lcout(acadc_skipCount_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55153),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i4_LC_14_16_0.C_ON=1'b0;
    defparam buf_control_i4_LC_14_16_0.SEQ_MODE=4'b1000;
    defparam buf_control_i4_LC_14_16_0.LUT_INIT=16'b1110111000100010;
    LogicCell40 buf_control_i4_LC_14_16_0 (
            .in0(N__44744),
            .in1(N__43847),
            .in2(_gnd_net_),
            .in3(N__42135),
            .lcout(VDC_RNG0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55168),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i15_LC_14_16_1.C_ON=1'b0;
    defparam acadc_skipCount_i15_LC_14_16_1.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i15_LC_14_16_1.LUT_INIT=16'b1011101110001000;
    LogicCell40 acadc_skipCount_i15_LC_14_16_1 (
            .in0(N__45766),
            .in1(N__39273),
            .in2(_gnd_net_),
            .in3(N__36588),
            .lcout(acadc_skipCount_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55168),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_7_i26_3_lut_LC_14_16_2.C_ON=1'b0;
    defparam mux_129_Mux_7_i26_3_lut_LC_14_16_2.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_7_i26_3_lut_LC_14_16_2.LUT_INIT=16'b1100110010101010;
    LogicCell40 mux_129_Mux_7_i26_3_lut_LC_14_16_2 (
            .in0(N__47376),
            .in1(N__36682),
            .in2(_gnd_net_),
            .in3(N__56954),
            .lcout(n26_adj_1623),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i14_LC_14_16_3.C_ON=1'b0;
    defparam acadc_skipCount_i14_LC_14_16_3.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i14_LC_14_16_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 acadc_skipCount_i14_LC_14_16_3 (
            .in0(N__41528),
            .in1(N__39272),
            .in2(_gnd_net_),
            .in3(N__36657),
            .lcout(acadc_skipCount_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55168),
            .ce(),
            .sr(_gnd_net_));
    defparam i6422_3_lut_LC_14_16_4.C_ON=1'b0;
    defparam i6422_3_lut_LC_14_16_4.SEQ_MODE=4'b0000;
    defparam i6422_3_lut_LC_14_16_4.LUT_INIT=16'b1100110010101010;
    LogicCell40 i6422_3_lut_LC_14_16_4 (
            .in0(N__42788),
            .in1(N__41861),
            .in2(_gnd_net_),
            .in3(N__43277),
            .lcout(n8_adj_1545),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i6_LC_14_16_5.C_ON=1'b0;
    defparam buf_control_i6_LC_14_16_5.SEQ_MODE=4'b1000;
    defparam buf_control_i6_LC_14_16_5.LUT_INIT=16'b1111000010101010;
    LogicCell40 buf_control_i6_LC_14_16_5 (
            .in0(N__55949),
            .in1(_gnd_net_),
            .in2(N__41535),
            .in3(N__43848),
            .lcout(buf_control_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55168),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_4_lut_adj_175_LC_14_16_6.C_ON=1'b0;
    defparam i1_2_lut_4_lut_adj_175_LC_14_16_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_4_lut_adj_175_LC_14_16_6.LUT_INIT=16'b1111111111111011;
    LogicCell40 i1_2_lut_4_lut_adj_175_LC_14_16_6 (
            .in0(N__57493),
            .in1(N__56955),
            .in2(N__45382),
            .in3(N__47836),
            .lcout(n20626),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i8_4_lut_LC_14_16_7.C_ON=1'b0;
    defparam i8_4_lut_LC_14_16_7.SEQ_MODE=4'b0000;
    defparam i8_4_lut_LC_14_16_7.LUT_INIT=16'b0111101111011110;
    LogicCell40 i8_4_lut_LC_14_16_7 (
            .in0(N__36628),
            .in1(N__36613),
            .in2(N__36921),
            .in3(N__36587),
            .lcout(n24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i1_LC_14_17_0.C_ON=1'b0;
    defparam acadc_skipCount_i1_LC_14_17_0.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i1_LC_14_17_0.LUT_INIT=16'b0011000010111000;
    LogicCell40 acadc_skipCount_i1_LC_14_17_0 (
            .in0(N__43374),
            .in1(N__39285),
            .in2(N__36568),
            .in3(N__52087),
            .lcout(acadc_skipCount_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55183),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_301_LC_14_17_1.C_ON=1'b0;
    defparam i1_4_lut_adj_301_LC_14_17_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_301_LC_14_17_1.LUT_INIT=16'b1100000011000100;
    LogicCell40 i1_4_lut_adj_301_LC_14_17_1 (
            .in0(N__36538),
            .in1(N__54675),
            .in2(N__52159),
            .in3(N__41626),
            .lcout(n12391),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19350_LC_14_17_2.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19350_LC_14_17_2.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19350_LC_14_17_2.LUT_INIT=16'b1110011010100010;
    LogicCell40 comm_cmd_1__bdd_4_lut_19350_LC_14_17_2 (
            .in0(N__57539),
            .in1(N__47844),
            .in2(N__37003),
            .in3(N__36991),
            .lcout(),
            .ltout(n21949_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n21949_bdd_4_lut_LC_14_17_3.C_ON=1'b0;
    defparam n21949_bdd_4_lut_LC_14_17_3.SEQ_MODE=4'b0000;
    defparam n21949_bdd_4_lut_LC_14_17_3.LUT_INIT=16'b1110010111100000;
    LogicCell40 n21949_bdd_4_lut_LC_14_17_3 (
            .in0(N__47845),
            .in1(N__41569),
            .in2(N__36985),
            .in3(N__36982),
            .lcout(),
            .ltout(n21952_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1535641_i1_3_lut_LC_14_17_4.C_ON=1'b0;
    defparam i1535641_i1_3_lut_LC_14_17_4.SEQ_MODE=4'b0000;
    defparam i1535641_i1_3_lut_LC_14_17_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 i1535641_i1_3_lut_LC_14_17_4 (
            .in0(_gnd_net_),
            .in1(N__36964),
            .in2(N__36952),
            .in3(N__56317),
            .lcout(n30_adj_1624),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i4_LC_14_17_5.C_ON=1'b0;
    defparam acadc_skipCount_i4_LC_14_17_5.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i4_LC_14_17_5.LUT_INIT=16'b0101110100001000;
    LogicCell40 acadc_skipCount_i4_LC_14_17_5 (
            .in0(N__39286),
            .in1(N__46647),
            .in2(N__52160),
            .in3(N__36947),
            .lcout(acadc_skipCount_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55183),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i9_LC_14_17_7.C_ON=1'b0;
    defparam acadc_skipCount_i9_LC_14_17_7.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i9_LC_14_17_7.LUT_INIT=16'b0101110100001000;
    LogicCell40 acadc_skipCount_i9_LC_14_17_7 (
            .in0(N__39287),
            .in1(N__44127),
            .in2(N__52161),
            .in3(N__36920),
            .lcout(acadc_skipCount_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55183),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i7_LC_14_18_0.C_ON=1'b0;
    defparam comm_buf_1__i7_LC_14_18_0.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i7_LC_14_18_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 comm_buf_1__i7_LC_14_18_0 (
            .in0(N__36894),
            .in1(N__54090),
            .in2(_gnd_net_),
            .in3(N__36814),
            .lcout(comm_buf_1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55197),
            .ce(N__38540),
            .sr(N__36803));
    defparam \SIG_DDS.i19068_4_lut_LC_14_19_3 .C_ON=1'b0;
    defparam \SIG_DDS.i19068_4_lut_LC_14_19_3 .SEQ_MODE=4'b0000;
    defparam \SIG_DDS.i19068_4_lut_LC_14_19_3 .LUT_INIT=16'b1010101000100110;
    LogicCell40 \SIG_DDS.i19068_4_lut_LC_14_19_3  (
            .in0(N__55866),
            .in1(N__55737),
            .in2(N__53025),
            .in3(N__55628),
            .lcout(\SIG_DDS.n12700 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i3_LC_14_19_4 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i3_LC_14_19_4 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i3_LC_14_19_4 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \SIG_DDS.tmp_buf_i3_LC_14_19_4  (
            .in0(N__55629),
            .in1(N__55867),
            .in2(N__36724),
            .in3(N__36697),
            .lcout(\SIG_DDS.tmp_buf_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55210),
            .ce(N__40314),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i4_LC_14_19_5 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i4_LC_14_19_5 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i4_LC_14_19_5 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \SIG_DDS.tmp_buf_i4_LC_14_19_5  (
            .in0(N__55868),
            .in1(N__55630),
            .in2(N__36691),
            .in3(N__42712),
            .lcout(\SIG_DDS.tmp_buf_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55210),
            .ce(N__40314),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i5_LC_14_19_6 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i5_LC_14_19_6 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i5_LC_14_19_6 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \SIG_DDS.tmp_buf_i5_LC_14_19_6  (
            .in0(N__55631),
            .in1(N__55869),
            .in2(N__37156),
            .in3(N__43065),
            .lcout(\SIG_DDS.tmp_buf_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55210),
            .ce(N__40314),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i6_LC_14_19_7 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i6_LC_14_19_7 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i6_LC_14_19_7 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \SIG_DDS.tmp_buf_i6_LC_14_19_7  (
            .in0(N__55870),
            .in1(N__55632),
            .in2(N__37147),
            .in3(N__42658),
            .lcout(\SIG_DDS.tmp_buf_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55210),
            .ce(N__40314),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.t0on_i0_LC_15_3_0 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i0_LC_15_3_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i0_LC_15_3_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i0_LC_15_3_0  (
            .in0(_gnd_net_),
            .in1(N__37126),
            .in2(_gnd_net_),
            .in3(N__37114),
            .lcout(\ADC_VDC.genclk.t0on_0 ),
            .ltout(),
            .carryin(bfn_15_3_0_),
            .carryout(\ADC_VDC.genclk.n19425 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__37483),
            .sr(N__37452));
    defparam \ADC_VDC.genclk.t0on_i1_LC_15_3_1 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i1_LC_15_3_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i1_LC_15_3_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i1_LC_15_3_1  (
            .in0(_gnd_net_),
            .in1(N__37111),
            .in2(N__52828),
            .in3(N__37099),
            .lcout(\ADC_VDC.genclk.t0on_1 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19425 ),
            .carryout(\ADC_VDC.genclk.n19426 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__37483),
            .sr(N__37452));
    defparam \ADC_VDC.genclk.t0on_i2_LC_15_3_2 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i2_LC_15_3_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i2_LC_15_3_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i2_LC_15_3_2  (
            .in0(_gnd_net_),
            .in1(N__52776),
            .in2(N__37096),
            .in3(N__37081),
            .lcout(\ADC_VDC.genclk.t0on_2 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19426 ),
            .carryout(\ADC_VDC.genclk.n19427 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__37483),
            .sr(N__37452));
    defparam \ADC_VDC.genclk.t0on_i3_LC_15_3_3 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i3_LC_15_3_3 .SEQ_MODE=4'b1001;
    defparam \ADC_VDC.genclk.t0on_i3_LC_15_3_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i3_LC_15_3_3  (
            .in0(_gnd_net_),
            .in1(N__37078),
            .in2(N__52829),
            .in3(N__37066),
            .lcout(\ADC_VDC.genclk.t0on_3 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19427 ),
            .carryout(\ADC_VDC.genclk.n19428 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__37483),
            .sr(N__37452));
    defparam \ADC_VDC.genclk.t0on_i4_LC_15_3_4 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i4_LC_15_3_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i4_LC_15_3_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i4_LC_15_3_4  (
            .in0(_gnd_net_),
            .in1(N__52780),
            .in2(N__37062),
            .in3(N__37042),
            .lcout(\ADC_VDC.genclk.t0on_4 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19428 ),
            .carryout(\ADC_VDC.genclk.n19429 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__37483),
            .sr(N__37452));
    defparam \ADC_VDC.genclk.t0on_i5_LC_15_3_5 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i5_LC_15_3_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i5_LC_15_3_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i5_LC_15_3_5  (
            .in0(_gnd_net_),
            .in1(N__37038),
            .in2(N__52830),
            .in3(N__37024),
            .lcout(\ADC_VDC.genclk.t0on_5 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19429 ),
            .carryout(\ADC_VDC.genclk.n19430 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__37483),
            .sr(N__37452));
    defparam \ADC_VDC.genclk.t0on_i6_LC_15_3_6 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i6_LC_15_3_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i6_LC_15_3_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i6_LC_15_3_6  (
            .in0(_gnd_net_),
            .in1(N__52784),
            .in2(N__37021),
            .in3(N__37006),
            .lcout(\ADC_VDC.genclk.t0on_6 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19430 ),
            .carryout(\ADC_VDC.genclk.n19431 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__37483),
            .sr(N__37452));
    defparam \ADC_VDC.genclk.t0on_i7_LC_15_3_7 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i7_LC_15_3_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i7_LC_15_3_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i7_LC_15_3_7  (
            .in0(_gnd_net_),
            .in1(N__37287),
            .in2(N__52831),
            .in3(N__37273),
            .lcout(\ADC_VDC.genclk.t0on_7 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19431 ),
            .carryout(\ADC_VDC.genclk.n19432 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__37483),
            .sr(N__37452));
    defparam \ADC_VDC.genclk.t0on_i8_LC_15_4_0 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i8_LC_15_4_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i8_LC_15_4_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i8_LC_15_4_0  (
            .in0(_gnd_net_),
            .in1(N__37270),
            .in2(N__52794),
            .in3(N__37258),
            .lcout(\ADC_VDC.genclk.t0on_8 ),
            .ltout(),
            .carryin(bfn_15_4_0_),
            .carryout(\ADC_VDC.genclk.n19433 ),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__37482),
            .sr(N__37456));
    defparam \ADC_VDC.genclk.t0on_i9_LC_15_4_1 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i9_LC_15_4_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i9_LC_15_4_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i9_LC_15_4_1  (
            .in0(_gnd_net_),
            .in1(N__52719),
            .in2(N__37255),
            .in3(N__37240),
            .lcout(\ADC_VDC.genclk.t0on_9 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19433 ),
            .carryout(\ADC_VDC.genclk.n19434 ),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__37482),
            .sr(N__37456));
    defparam \ADC_VDC.genclk.t0on_i10_LC_15_4_2 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i10_LC_15_4_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i10_LC_15_4_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i10_LC_15_4_2  (
            .in0(_gnd_net_),
            .in1(N__37237),
            .in2(N__52791),
            .in3(N__37225),
            .lcout(\ADC_VDC.genclk.t0on_10 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19434 ),
            .carryout(\ADC_VDC.genclk.n19435 ),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__37482),
            .sr(N__37456));
    defparam \ADC_VDC.genclk.t0on_i11_LC_15_4_3 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i11_LC_15_4_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i11_LC_15_4_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i11_LC_15_4_3  (
            .in0(_gnd_net_),
            .in1(N__52707),
            .in2(N__37222),
            .in3(N__37207),
            .lcout(\ADC_VDC.genclk.t0on_11 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19435 ),
            .carryout(\ADC_VDC.genclk.n19436 ),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__37482),
            .sr(N__37456));
    defparam \ADC_VDC.genclk.t0on_i12_LC_15_4_4 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i12_LC_15_4_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i12_LC_15_4_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i12_LC_15_4_4  (
            .in0(_gnd_net_),
            .in1(N__37204),
            .in2(N__52792),
            .in3(N__37192),
            .lcout(\ADC_VDC.genclk.t0on_12 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19436 ),
            .carryout(\ADC_VDC.genclk.n19437 ),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__37482),
            .sr(N__37456));
    defparam \ADC_VDC.genclk.t0on_i13_LC_15_4_5 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i13_LC_15_4_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i13_LC_15_4_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i13_LC_15_4_5  (
            .in0(_gnd_net_),
            .in1(N__52711),
            .in2(N__37189),
            .in3(N__37174),
            .lcout(\ADC_VDC.genclk.t0on_13 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19437 ),
            .carryout(\ADC_VDC.genclk.n19438 ),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__37482),
            .sr(N__37456));
    defparam \ADC_VDC.genclk.t0on_i14_LC_15_4_6 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i14_LC_15_4_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i14_LC_15_4_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i14_LC_15_4_6  (
            .in0(_gnd_net_),
            .in1(N__37171),
            .in2(N__52793),
            .in3(N__37159),
            .lcout(\ADC_VDC.genclk.t0on_14 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19438 ),
            .carryout(\ADC_VDC.genclk.n19439 ),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__37482),
            .sr(N__37456));
    defparam \ADC_VDC.genclk.t0on_i15_LC_15_4_7 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.t0on_i15_LC_15_4_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i15_LC_15_4_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ADC_VDC.genclk.t0on_i15_LC_15_4_7  (
            .in0(N__37497),
            .in1(N__52715),
            .in2(_gnd_net_),
            .in3(N__37501),
            .lcout(\ADC_VDC.genclk.t0on_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__37482),
            .sr(N__37456));
    defparam \comm_spi.imosi_44_12183_12184_set_LC_15_5_0 .C_ON=1'b0;
    defparam \comm_spi.imosi_44_12183_12184_set_LC_15_5_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.imosi_44_12183_12184_set_LC_15_5_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \comm_spi.imosi_44_12183_12184_set_LC_15_5_0  (
            .in0(N__37355),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\comm_spi.n14585 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55075),
            .ce(),
            .sr(N__37363));
    defparam \comm_spi.MISO_48_12187_12188_set_LC_15_6_0 .C_ON=1'b0;
    defparam \comm_spi.MISO_48_12187_12188_set_LC_15_6_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.MISO_48_12187_12188_set_LC_15_6_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \comm_spi.MISO_48_12187_12188_set_LC_15_6_0  (
            .in0(N__44323),
            .in1(N__44310),
            .in2(_gnd_net_),
            .in3(N__44270),
            .lcout(\comm_spi.n14589 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.MISO_48_12187_12188_setC_net ),
            .ce(),
            .sr(N__40256));
    defparam \comm_spi.RESET_I_0_105_2_lut_LC_15_6_1 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_105_2_lut_LC_15_6_1 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_105_2_lut_LC_15_6_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \comm_spi.RESET_I_0_105_2_lut_LC_15_6_1  (
            .in0(N__55424),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37376),
            .lcout(\comm_spi.data_tx_7__N_781 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_92_2_lut_LC_15_6_2 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_92_2_lut_LC_15_6_2 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_92_2_lut_LC_15_6_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \comm_spi.RESET_I_0_92_2_lut_LC_15_6_2  (
            .in0(_gnd_net_),
            .in1(N__37395),
            .in2(_gnd_net_),
            .in3(N__55421),
            .lcout(\comm_spi.data_tx_7__N_758 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_97_2_lut_LC_15_6_3 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_97_2_lut_LC_15_6_3 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_97_2_lut_LC_15_6_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \comm_spi.RESET_I_0_97_2_lut_LC_15_6_3  (
            .in0(N__55426),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37377),
            .lcout(\comm_spi.data_tx_7__N_763 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i19179_4_lut_3_lut_LC_15_6_4 .C_ON=1'b0;
    defparam \comm_spi.i19179_4_lut_3_lut_LC_15_6_4 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19179_4_lut_3_lut_LC_15_6_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.i19179_4_lut_3_lut_LC_15_6_4  (
            .in0(N__37378),
            .in1(N__37718),
            .in2(_gnd_net_),
            .in3(N__55427),
            .lcout(\comm_spi.n22644 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_88_2_lut_LC_15_6_5 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_88_2_lut_LC_15_6_5 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_88_2_lut_LC_15_6_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \comm_spi.RESET_I_0_88_2_lut_LC_15_6_5  (
            .in0(N__55423),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37356),
            .lcout(\comm_spi.imosi_N_744 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_89_2_lut_LC_15_6_6 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_89_2_lut_LC_15_6_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_89_2_lut_LC_15_6_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \comm_spi.RESET_I_0_89_2_lut_LC_15_6_6  (
            .in0(N__37357),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55422),
            .lcout(\comm_spi.imosi_N_745 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_95_2_lut_LC_15_6_7 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_95_2_lut_LC_15_6_7 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_95_2_lut_LC_15_6_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \comm_spi.RESET_I_0_95_2_lut_LC_15_6_7  (
            .in0(N__55425),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53164),
            .lcout(\comm_spi.data_tx_7__N_761 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i3_12209_12210_reset_LC_15_7_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i3_12209_12210_reset_LC_15_7_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i3_12209_12210_reset_LC_15_7_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i3_12209_12210_reset_LC_15_7_0  (
            .in0(N__37719),
            .in1(N__37662),
            .in2(_gnd_net_),
            .in3(N__37689),
            .lcout(\comm_spi.n14612 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52407),
            .ce(),
            .sr(N__37702));
    defparam \comm_spi.data_tx_i2_12205_12206_reset_LC_15_8_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i2_12205_12206_reset_LC_15_8_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i2_12205_12206_reset_LC_15_8_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i2_12205_12206_reset_LC_15_8_0  (
            .in0(N__50220),
            .in1(N__52468),
            .in2(_gnd_net_),
            .in3(N__52518),
            .lcout(\comm_spi.n14608 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52424),
            .ce(),
            .sr(N__37678));
    defparam \comm_spi.data_tx_i2_12205_12206_set_LC_15_9_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i2_12205_12206_set_LC_15_9_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i2_12205_12206_set_LC_15_9_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i2_12205_12206_set_LC_15_9_0  (
            .in0(N__50221),
            .in1(N__52461),
            .in2(_gnd_net_),
            .in3(N__52522),
            .lcout(\comm_spi.n14607 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52442),
            .ce(),
            .sr(N__37645));
    defparam \comm_spi.i19184_4_lut_3_lut_LC_15_9_1 .C_ON=1'b0;
    defparam \comm_spi.i19184_4_lut_3_lut_LC_15_9_1 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19184_4_lut_3_lut_LC_15_9_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.i19184_4_lut_3_lut_LC_15_9_1  (
            .in0(N__55429),
            .in1(N__37633),
            .in2(_gnd_net_),
            .in3(N__46191),
            .lcout(\comm_spi.n22641 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i19189_4_lut_3_lut_LC_15_9_2 .C_ON=1'b0;
    defparam \comm_spi.i19189_4_lut_3_lut_LC_15_9_2 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19189_4_lut_3_lut_LC_15_9_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \comm_spi.i19189_4_lut_3_lut_LC_15_9_2  (
            .in0(N__46257),
            .in1(N__53160),
            .in2(_gnd_net_),
            .in3(N__55430),
            .lcout(\comm_spi.n22638 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15011_2_lut_LC_15_9_4.C_ON=1'b0;
    defparam i15011_2_lut_LC_15_9_4.SEQ_MODE=4'b0000;
    defparam i15011_2_lut_LC_15_9_4.LUT_INIT=16'b1010000010100000;
    LogicCell40 i15011_2_lut_LC_15_9_4 (
            .in0(N__41169),
            .in1(_gnd_net_),
            .in2(N__41197),
            .in3(_gnd_net_),
            .lcout(n17393),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18832_2_lut_LC_15_9_5.C_ON=1'b0;
    defparam i18832_2_lut_LC_15_9_5.SEQ_MODE=4'b0000;
    defparam i18832_2_lut_LC_15_9_5.LUT_INIT=16'b0011001100000000;
    LogicCell40 i18832_2_lut_LC_15_9_5 (
            .in0(_gnd_net_),
            .in1(N__37606),
            .in2(_gnd_net_),
            .in3(N__38897),
            .lcout(n21067),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_4_lut_adj_229_LC_15_10_0.C_ON=1'b0;
    defparam i1_3_lut_4_lut_adj_229_LC_15_10_0.SEQ_MODE=4'b0000;
    defparam i1_3_lut_4_lut_adj_229_LC_15_10_0.LUT_INIT=16'b1101111111011101;
    LogicCell40 i1_3_lut_4_lut_adj_229_LC_15_10_0 (
            .in0(N__51239),
            .in1(N__54486),
            .in2(N__54001),
            .in3(N__37516),
            .lcout(),
            .ltout(n11839_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_152_LC_15_10_1.C_ON=1'b0;
    defparam i1_4_lut_adj_152_LC_15_10_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_152_LC_15_10_1.LUT_INIT=16'b1100000010000000;
    LogicCell40 i1_4_lut_adj_152_LC_15_10_1 (
            .in0(N__46500),
            .in1(N__49216),
            .in2(N__37909),
            .in3(N__37905),
            .lcout(n11846),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_284_LC_15_10_2.C_ON=1'b0;
    defparam i1_4_lut_adj_284_LC_15_10_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_284_LC_15_10_2.LUT_INIT=16'b1111000001000000;
    LogicCell40 i1_4_lut_adj_284_LC_15_10_2 (
            .in0(N__51240),
            .in1(N__37906),
            .in2(N__49235),
            .in3(N__54487),
            .lcout(n14722),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6817_2_lut_LC_15_10_3.C_ON=1'b0;
    defparam i6817_2_lut_LC_15_10_3.SEQ_MODE=4'b0000;
    defparam i6817_2_lut_LC_15_10_3.LUT_INIT=16'b0101010100000000;
    LogicCell40 i6817_2_lut_LC_15_10_3 (
            .in0(N__53838),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53487),
            .lcout(n9222),
            .ltout(n9222_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_303_LC_15_10_4.C_ON=1'b0;
    defparam i1_4_lut_adj_303_LC_15_10_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_303_LC_15_10_4.LUT_INIT=16'b1010100010001000;
    LogicCell40 i1_4_lut_adj_303_LC_15_10_4 (
            .in0(N__49215),
            .in1(N__54485),
            .in2(N__37894),
            .in3(N__51238),
            .lcout(n12322),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i41_4_lut_LC_15_10_5.C_ON=1'b0;
    defparam i41_4_lut_LC_15_10_5.SEQ_MODE=4'b0000;
    defparam i41_4_lut_LC_15_10_5.LUT_INIT=16'b0100000000101100;
    LogicCell40 i41_4_lut_LC_15_10_5 (
            .in0(N__56945),
            .in1(N__47851),
            .in2(N__57447),
            .in3(N__56270),
            .lcout(),
            .ltout(n24_adj_1579_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18910_2_lut_LC_15_10_6.C_ON=1'b0;
    defparam i18910_2_lut_LC_15_10_6.SEQ_MODE=4'b0000;
    defparam i18910_2_lut_LC_15_10_6.LUT_INIT=16'b1111000000000000;
    LogicCell40 i18910_2_lut_LC_15_10_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__37891),
            .in3(N__44401),
            .lcout(),
            .ltout(n21079_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i42_4_lut_LC_15_10_7.C_ON=1'b0;
    defparam i42_4_lut_LC_15_10_7.SEQ_MODE=4'b0000;
    defparam i42_4_lut_LC_15_10_7.LUT_INIT=16'b0111001001010000;
    LogicCell40 i42_4_lut_LC_15_10_7 (
            .in0(N__53839),
            .in1(N__50078),
            .in2(N__37888),
            .in3(N__46581),
            .lcout(n16_adj_1570),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15209_2_lut_3_lut_LC_15_11_0.C_ON=1'b0;
    defparam i15209_2_lut_3_lut_LC_15_11_0.SEQ_MODE=4'b0000;
    defparam i15209_2_lut_3_lut_LC_15_11_0.LUT_INIT=16'b0000000001000100;
    LogicCell40 i15209_2_lut_3_lut_LC_15_11_0 (
            .in0(N__53874),
            .in1(N__43347),
            .in2(_gnd_net_),
            .in3(N__51207),
            .lcout(n14_adj_1529),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i15_LC_15_11_1 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i15_LC_15_11_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i15_LC_15_11_1 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i15_LC_15_11_1  (
            .in0(N__45179),
            .in1(N__37871),
            .in2(N__48358),
            .in3(N__38767),
            .lcout(cmd_rdadctmp_15_adj_1428),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55120),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_291_LC_15_11_2.C_ON=1'b0;
    defparam i1_4_lut_adj_291_LC_15_11_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_291_LC_15_11_2.LUT_INIT=16'b1000110010001000;
    LogicCell40 i1_4_lut_adj_291_LC_15_11_2 (
            .in0(N__49910),
            .in1(N__49860),
            .in2(N__53521),
            .in3(N__38131),
            .lcout(n12080),
            .ltout(n12080_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12352_2_lut_LC_15_11_3.C_ON=1'b0;
    defparam i12352_2_lut_LC_15_11_3.SEQ_MODE=4'b0000;
    defparam i12352_2_lut_LC_15_11_3.LUT_INIT=16'b1111000000000000;
    LogicCell40 i12352_2_lut_LC_15_11_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38125),
            .in3(N__54488),
            .lcout(n14749),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22129_bdd_4_lut_LC_15_11_4.C_ON=1'b0;
    defparam n22129_bdd_4_lut_LC_15_11_4.SEQ_MODE=4'b0000;
    defparam n22129_bdd_4_lut_LC_15_11_4.LUT_INIT=16'b1110111001010000;
    LogicCell40 n22129_bdd_4_lut_LC_15_11_4 (
            .in0(N__49523),
            .in1(N__38122),
            .in2(N__43525),
            .in3(N__38047),
            .lcout(n22132),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_299_LC_15_11_5.C_ON=1'b0;
    defparam i1_3_lut_adj_299_LC_15_11_5.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_299_LC_15_11_5.LUT_INIT=16'b1010101010001000;
    LogicCell40 i1_3_lut_adj_299_LC_15_11_5 (
            .in0(N__49859),
            .in1(N__49909),
            .in2(_gnd_net_),
            .in3(N__51454),
            .lcout(n12206),
            .ltout(n12206_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12373_2_lut_LC_15_11_6.C_ON=1'b0;
    defparam i12373_2_lut_LC_15_11_6.SEQ_MODE=4'b0000;
    defparam i12373_2_lut_LC_15_11_6.LUT_INIT=16'b1010000010100000;
    LogicCell40 i12373_2_lut_LC_15_11_6 (
            .in0(N__54489),
            .in1(_gnd_net_),
            .in2(N__38095),
            .in3(_gnd_net_),
            .lcout(n14770),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_2__bdd_4_lut_LC_15_11_7.C_ON=1'b0;
    defparam comm_index_2__bdd_4_lut_LC_15_11_7.SEQ_MODE=4'b0000;
    defparam comm_index_2__bdd_4_lut_LC_15_11_7.LUT_INIT=16'b1101100010101010;
    LogicCell40 comm_index_2__bdd_4_lut_LC_15_11_7 (
            .in0(N__50087),
            .in1(N__38083),
            .in2(N__38056),
            .in3(N__49522),
            .lcout(n22129),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_5_i22_3_lut_LC_15_12_0.C_ON=1'b0;
    defparam mux_130_Mux_5_i22_3_lut_LC_15_12_0.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_5_i22_3_lut_LC_15_12_0.LUT_INIT=16'b1100110010101010;
    LogicCell40 mux_130_Mux_5_i22_3_lut_LC_15_12_0 (
            .in0(N__49077),
            .in1(N__38275),
            .in2(_gnd_net_),
            .in3(N__47848),
            .lcout(),
            .ltout(n22_adj_1599_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_5_i30_3_lut_LC_15_12_1.C_ON=1'b0;
    defparam mux_130_Mux_5_i30_3_lut_LC_15_12_1.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_5_i30_3_lut_LC_15_12_1.LUT_INIT=16'b1010101011110000;
    LogicCell40 mux_130_Mux_5_i30_3_lut_LC_15_12_1 (
            .in0(N__38041),
            .in1(_gnd_net_),
            .in2(N__38029),
            .in3(N__56259),
            .lcout(),
            .ltout(n30_adj_1600_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_2__i5_LC_15_12_2.C_ON=1'b0;
    defparam comm_buf_2__i5_LC_15_12_2.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i5_LC_15_12_2.LUT_INIT=16'b1111110000110000;
    LogicCell40 comm_buf_2__i5_LC_15_12_2 (
            .in0(_gnd_net_),
            .in1(N__54033),
            .in2(N__38026),
            .in3(N__37981),
            .lcout(comm_buf_2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55129),
            .ce(N__37920),
            .sr(N__38346));
    defparam mux_130_Mux_5_i19_3_lut_LC_15_12_3.C_ON=1'b0;
    defparam mux_130_Mux_5_i19_3_lut_LC_15_12_3.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_5_i19_3_lut_LC_15_12_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_130_Mux_5_i19_3_lut_LC_15_12_3 (
            .in0(N__56953),
            .in1(N__38329),
            .in2(_gnd_net_),
            .in3(N__38303),
            .lcout(n19_adj_1598),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_2__bdd_4_lut_19491_LC_15_12_4.C_ON=1'b0;
    defparam comm_index_2__bdd_4_lut_19491_LC_15_12_4.SEQ_MODE=4'b0000;
    defparam comm_index_2__bdd_4_lut_19491_LC_15_12_4.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_index_2__bdd_4_lut_19491_LC_15_12_4 (
            .in0(N__38269),
            .in1(N__50088),
            .in2(N__38263),
            .in3(N__49524),
            .lcout(),
            .ltout(n22123_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22123_bdd_4_lut_LC_15_12_5.C_ON=1'b0;
    defparam n22123_bdd_4_lut_LC_15_12_5.SEQ_MODE=4'b0000;
    defparam n22123_bdd_4_lut_LC_15_12_5.LUT_INIT=16'b1110010111100000;
    LogicCell40 n22123_bdd_4_lut_LC_15_12_5 (
            .in0(N__49525),
            .in1(N__38242),
            .in2(N__38224),
            .in3(N__44871),
            .lcout(n22126),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_283_LC_15_12_6.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_283_LC_15_12_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_283_LC_15_12_6.LUT_INIT=16'b1011101111111111;
    LogicCell40 i1_2_lut_3_lut_adj_283_LC_15_12_6 (
            .in0(N__38209),
            .in1(N__56952),
            .in2(_gnd_net_),
            .in3(N__56260),
            .lcout(n11324),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_272_LC_15_12_7.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_272_LC_15_12_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_272_LC_15_12_7.LUT_INIT=16'b1111111110111011;
    LogicCell40 i1_2_lut_3_lut_adj_272_LC_15_12_7 (
            .in0(N__53499),
            .in1(N__56258),
            .in2(_gnd_net_),
            .in3(N__38208),
            .lcout(n20613),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i2_LC_15_13_0.C_ON=1'b0;
    defparam buf_control_i2_LC_15_13_0.SEQ_MODE=4'b1000;
    defparam buf_control_i2_LC_15_13_0.LUT_INIT=16'b0101110100001000;
    LogicCell40 buf_control_i2_LC_15_13_0 (
            .in0(N__43864),
            .in1(N__38719),
            .in2(N__52147),
            .in3(N__38162),
            .lcout(SELIRNG0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55141),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i5_LC_15_13_1.C_ON=1'b0;
    defparam req_data_cnt_i5_LC_15_13_1.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i5_LC_15_13_1.LUT_INIT=16'b1011101110001000;
    LogicCell40 req_data_cnt_i5_LC_15_13_1 (
            .in0(N__50136),
            .in1(N__42005),
            .in2(_gnd_net_),
            .in3(N__38417),
            .lcout(req_data_cnt_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55141),
            .ce(),
            .sr(_gnd_net_));
    defparam i15204_2_lut_3_lut_LC_15_13_2.C_ON=1'b0;
    defparam i15204_2_lut_3_lut_LC_15_13_2.SEQ_MODE=4'b0000;
    defparam i15204_2_lut_3_lut_LC_15_13_2.LUT_INIT=16'b0001000100000000;
    LogicCell40 i15204_2_lut_3_lut_LC_15_13_2 (
            .in0(N__54027),
            .in1(N__51282),
            .in2(_gnd_net_),
            .in3(N__44108),
            .lcout(n14_adj_1552),
            .ltout(n14_adj_1552_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i9_LC_15_13_3.C_ON=1'b0;
    defparam req_data_cnt_i9_LC_15_13_3.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i9_LC_15_13_3.LUT_INIT=16'b1111001111000000;
    LogicCell40 req_data_cnt_i9_LC_15_13_3 (
            .in0(_gnd_net_),
            .in1(N__42006),
            .in2(N__38134),
            .in3(N__41646),
            .lcout(req_data_cnt_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55141),
            .ce(),
            .sr(_gnd_net_));
    defparam i15202_2_lut_3_lut_LC_15_13_4.C_ON=1'b0;
    defparam i15202_2_lut_3_lut_LC_15_13_4.SEQ_MODE=4'b0000;
    defparam i15202_2_lut_3_lut_LC_15_13_4.LUT_INIT=16'b0000000000100010;
    LogicCell40 i15202_2_lut_3_lut_LC_15_13_4 (
            .in0(N__43796),
            .in1(N__51283),
            .in2(_gnd_net_),
            .in3(N__53957),
            .lcout(n14_adj_1550),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15_4_lut_adj_315_LC_15_13_5.C_ON=1'b0;
    defparam i15_4_lut_adj_315_LC_15_13_5.SEQ_MODE=4'b0000;
    defparam i15_4_lut_adj_315_LC_15_13_5.LUT_INIT=16'b1100111101000111;
    LogicCell40 i15_4_lut_adj_315_LC_15_13_5 (
            .in0(N__43299),
            .in1(N__54668),
            .in2(N__42353),
            .in3(N__52065),
            .lcout(n12254),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i15_LC_15_13_6.C_ON=1'b0;
    defparam req_data_cnt_i15_LC_15_13_6.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i15_LC_15_13_6.LUT_INIT=16'b1111010110100000;
    LogicCell40 req_data_cnt_i15_LC_15_13_6 (
            .in0(N__42004),
            .in1(_gnd_net_),
            .in2(N__45768),
            .in3(N__41684),
            .lcout(req_data_cnt_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55141),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_290_LC_15_13_7.C_ON=1'b0;
    defparam i1_4_lut_adj_290_LC_15_13_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_290_LC_15_13_7.LUT_INIT=16'b1000101010001000;
    LogicCell40 i1_4_lut_adj_290_LC_15_13_7 (
            .in0(N__49858),
            .in1(N__49908),
            .in2(N__53532),
            .in3(N__40813),
            .lcout(n12007),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i4_LC_15_14_0.C_ON=1'b0;
    defparam req_data_cnt_i4_LC_15_14_0.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i4_LC_15_14_0.LUT_INIT=16'b1111110000001100;
    LogicCell40 req_data_cnt_i4_LC_15_14_0 (
            .in0(_gnd_net_),
            .in1(N__38390),
            .in2(N__42025),
            .in3(N__38469),
            .lcout(req_data_cnt_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55154),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i1_LC_15_14_1.C_ON=1'b0;
    defparam req_data_cnt_i1_LC_15_14_1.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i1_LC_15_14_1.LUT_INIT=16'b1011101110001000;
    LogicCell40 req_data_cnt_i1_LC_15_14_1 (
            .in0(N__38442),
            .in1(N__42019),
            .in2(_gnd_net_),
            .in3(N__38373),
            .lcout(req_data_cnt_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55154),
            .ce(),
            .sr(_gnd_net_));
    defparam i4_4_lut_LC_15_14_2.C_ON=1'b0;
    defparam i4_4_lut_LC_15_14_2.SEQ_MODE=4'b0000;
    defparam i4_4_lut_LC_15_14_2.LUT_INIT=16'b0111110110111110;
    LogicCell40 i4_4_lut_LC_15_14_2 (
            .in0(N__46852),
            .in1(N__46782),
            .in2(N__38418),
            .in3(N__38825),
            .lcout(n20_adj_1496),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_adj_69_LC_15_14_3.C_ON=1'b0;
    defparam i2_4_lut_adj_69_LC_15_14_3.SEQ_MODE=4'b0000;
    defparam i2_4_lut_adj_69_LC_15_14_3.LUT_INIT=16'b0111101111011110;
    LogicCell40 i2_4_lut_adj_69_LC_15_14_3 (
            .in0(N__46812),
            .in1(N__46912),
            .in2(N__38394),
            .in3(N__38372),
            .lcout(),
            .ltout(n18_adj_1553_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i13_4_lut_LC_15_14_4.C_ON=1'b0;
    defparam i13_4_lut_LC_15_14_4.SEQ_MODE=4'b0000;
    defparam i13_4_lut_LC_15_14_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i13_4_lut_LC_15_14_4 (
            .in0(N__38359),
            .in1(N__41875),
            .in2(N__38353),
            .in3(N__41698),
            .lcout(),
            .ltout(n29_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_80_LC_15_14_5.C_ON=1'b0;
    defparam i1_3_lut_adj_80_LC_15_14_5.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_80_LC_15_14_5.LUT_INIT=16'b1100110011001111;
    LogicCell40 i1_3_lut_adj_80_LC_15_14_5 (
            .in0(_gnd_net_),
            .in1(N__38937),
            .in2(N__38902),
            .in3(N__42151),
            .lcout(n16_adj_1609),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i3_LC_15_14_6.C_ON=1'b0;
    defparam req_data_cnt_i3_LC_15_14_6.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i3_LC_15_14_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 req_data_cnt_i3_LC_15_14_6 (
            .in0(N__42020),
            .in1(N__38865),
            .in2(_gnd_net_),
            .in3(N__38826),
            .lcout(req_data_cnt_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55154),
            .ce(),
            .sr(_gnd_net_));
    defparam i5_4_lut_LC_15_15_0.C_ON=1'b0;
    defparam i5_4_lut_LC_15_15_0.SEQ_MODE=4'b0000;
    defparam i5_4_lut_LC_15_15_0.LUT_INIT=16'b0111110110111110;
    LogicCell40 i5_4_lut_LC_15_15_0 (
            .in0(N__38812),
            .in1(N__38794),
            .in2(N__38613),
            .in3(N__44717),
            .lcout(n21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_6__I_0_363_i9_2_lut_3_lut_LC_15_15_1.C_ON=1'b0;
    defparam comm_cmd_6__I_0_363_i9_2_lut_3_lut_LC_15_15_1.SEQ_MODE=4'b0000;
    defparam comm_cmd_6__I_0_363_i9_2_lut_3_lut_LC_15_15_1.LUT_INIT=16'b1111111111101110;
    LogicCell40 comm_cmd_6__I_0_363_i9_2_lut_3_lut_LC_15_15_1 (
            .in0(N__57548),
            .in1(N__56966),
            .in2(_gnd_net_),
            .in3(N__47843),
            .lcout(),
            .ltout(n9_adj_1408_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_271_LC_15_15_2.C_ON=1'b0;
    defparam i1_4_lut_adj_271_LC_15_15_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_271_LC_15_15_2.LUT_INIT=16'b1100110100000000;
    LogicCell40 i1_4_lut_adj_271_LC_15_15_2 (
            .in0(N__41622),
            .in1(N__51914),
            .in2(N__38770),
            .in3(N__54625),
            .lcout(n11901),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i12_LC_15_15_3.C_ON=1'b0;
    defparam acadc_skipCount_i12_LC_15_15_3.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i12_LC_15_15_3.LUT_INIT=16'b1100110010101010;
    LogicCell40 acadc_skipCount_i12_LC_15_15_3 (
            .in0(N__44718),
            .in1(N__42139),
            .in2(_gnd_net_),
            .in3(N__39315),
            .lcout(acadc_skipCount_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55169),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i6_LC_15_15_4 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i6_LC_15_15_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i6_LC_15_15_4 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i6_LC_15_15_4  (
            .in0(N__48314),
            .in1(N__48504),
            .in2(N__38763),
            .in3(N__40853),
            .lcout(buf_adcdata_vac_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55169),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i10_LC_15_15_5.C_ON=1'b0;
    defparam acadc_skipCount_i10_LC_15_15_5.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i10_LC_15_15_5.LUT_INIT=16'b0011000010101010;
    LogicCell40 acadc_skipCount_i10_LC_15_15_5 (
            .in0(N__38612),
            .in1(N__51978),
            .in2(N__38734),
            .in3(N__39316),
            .lcout(acadc_skipCount_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55169),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i12_LC_15_15_6.C_ON=1'b0;
    defparam req_data_cnt_i12_LC_15_15_6.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i12_LC_15_15_6.LUT_INIT=16'b1111010110100000;
    LogicCell40 req_data_cnt_i12_LC_15_15_6 (
            .in0(N__42024),
            .in1(_gnd_net_),
            .in2(N__42145),
            .in3(N__56397),
            .lcout(req_data_cnt_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55169),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i11_LC_15_15_7.C_ON=1'b0;
    defparam acadc_skipCount_i11_LC_15_15_7.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i11_LC_15_15_7.LUT_INIT=16'b0111001101000000;
    LogicCell40 acadc_skipCount_i11_LC_15_15_7 (
            .in0(N__51915),
            .in1(N__39317),
            .in2(N__43816),
            .in3(N__45470),
            .lcout(acadc_skipCount_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55169),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_276_LC_15_16_0.C_ON=1'b0;
    defparam i1_4_lut_adj_276_LC_15_16_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_276_LC_15_16_0.LUT_INIT=16'b1010000010100010;
    LogicCell40 i1_4_lut_adj_276_LC_15_16_0 (
            .in0(N__54624),
            .in1(N__45561),
            .in2(N__52062),
            .in3(N__45380),
            .lcout(n12367),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i4_LC_15_16_1.C_ON=1'b0;
    defparam data_index_i4_LC_15_16_1.SEQ_MODE=4'b1000;
    defparam data_index_i4_LC_15_16_1.LUT_INIT=16'b0101110100001000;
    LogicCell40 data_index_i4_LC_15_16_1 (
            .in0(N__54709),
            .in1(N__39043),
            .in2(N__52061),
            .in3(N__42490),
            .lcout(data_index_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55184),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_4_lut_adj_84_LC_15_16_2.C_ON=1'b0;
    defparam i3_4_lut_adj_84_LC_15_16_2.SEQ_MODE=4'b0000;
    defparam i3_4_lut_adj_84_LC_15_16_2.LUT_INIT=16'b1111111111111011;
    LogicCell40 i3_4_lut_adj_84_LC_15_16_2 (
            .in0(N__53522),
            .in1(N__47835),
            .in2(N__39183),
            .in3(N__57395),
            .lcout(n8780),
            .ltout(n8780_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i14930_3_lut_LC_15_16_3.C_ON=1'b0;
    defparam i14930_3_lut_LC_15_16_3.SEQ_MODE=4'b0000;
    defparam i14930_3_lut_LC_15_16_3.LUT_INIT=16'b1111110000001100;
    LogicCell40 i14930_3_lut_LC_15_16_3 (
            .in0(_gnd_net_),
            .in1(N__41347),
            .in2(N__39160),
            .in3(N__42840),
            .lcout(n17314),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12226_2_lut_LC_15_16_4.C_ON=1'b0;
    defparam i12226_2_lut_LC_15_16_4.SEQ_MODE=4'b0000;
    defparam i12226_2_lut_LC_15_16_4.LUT_INIT=16'b0101010100000000;
    LogicCell40 i12226_2_lut_LC_15_16_4 (
            .in0(N__39150),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48631),
            .lcout(n14632),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i7_LC_15_16_5.C_ON=1'b0;
    defparam buf_dds0_i7_LC_15_16_5.SEQ_MODE=4'b1000;
    defparam buf_dds0_i7_LC_15_16_5.LUT_INIT=16'b0101000011001100;
    LogicCell40 buf_dds0_i7_LC_15_16_5 (
            .in0(N__51951),
            .in1(N__39057),
            .in2(N__42615),
            .in3(N__45693),
            .lcout(buf_dds0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55184),
            .ce(),
            .sr(_gnd_net_));
    defparam i6402_3_lut_LC_15_16_6.C_ON=1'b0;
    defparam i6402_3_lut_LC_15_16_6.SEQ_MODE=4'b0000;
    defparam i6402_3_lut_LC_15_16_6.LUT_INIT=16'b1100110010101010;
    LogicCell40 i6402_3_lut_LC_15_16_6 (
            .in0(N__46654),
            .in1(N__42508),
            .in2(_gnd_net_),
            .in3(N__43284),
            .lcout(n8_adj_1541),
            .ltout(n8_adj_1541_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_354_Mux_4_i15_4_lut_LC_15_16_7.C_ON=1'b0;
    defparam comm_state_3__I_0_354_Mux_4_i15_4_lut_LC_15_16_7.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_354_Mux_4_i15_4_lut_LC_15_16_7.LUT_INIT=16'b0111001101000000;
    LogicCell40 comm_state_3__I_0_354_Mux_4_i15_4_lut_LC_15_16_7 (
            .in0(N__51950),
            .in1(N__54623),
            .in2(N__39037),
            .in3(N__42489),
            .lcout(data_index_9_N_212_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_count_i0_i0_LC_15_17_0.C_ON=1'b1;
    defparam data_count_i0_i0_LC_15_17_0.SEQ_MODE=4'b1000;
    defparam data_count_i0_i0_LC_15_17_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i0_LC_15_17_0 (
            .in0(_gnd_net_),
            .in1(N__46986),
            .in2(N__40097),
            .in3(_gnd_net_),
            .lcout(data_count_0),
            .ltout(),
            .carryin(bfn_15_17_0_),
            .carryout(n19287),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__48655),
            .sr(N__48586));
    defparam data_count_i0_i1_LC_15_17_1.C_ON=1'b1;
    defparam data_count_i0_i1_LC_15_17_1.SEQ_MODE=4'b1000;
    defparam data_count_i0_i1_LC_15_17_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i1_LC_15_17_1 (
            .in0(_gnd_net_),
            .in1(N__39986),
            .in2(_gnd_net_),
            .in3(N__39967),
            .lcout(data_count_1),
            .ltout(),
            .carryin(n19287),
            .carryout(n19288),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__48655),
            .sr(N__48586));
    defparam data_count_i0_i2_LC_15_17_2.C_ON=1'b1;
    defparam data_count_i0_i2_LC_15_17_2.SEQ_MODE=4'b1000;
    defparam data_count_i0_i2_LC_15_17_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i2_LC_15_17_2 (
            .in0(_gnd_net_),
            .in1(N__39881),
            .in2(_gnd_net_),
            .in3(N__39859),
            .lcout(data_count_2),
            .ltout(),
            .carryin(n19288),
            .carryout(n19289),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__48655),
            .sr(N__48586));
    defparam data_count_i0_i3_LC_15_17_3.C_ON=1'b1;
    defparam data_count_i0_i3_LC_15_17_3.SEQ_MODE=4'b1000;
    defparam data_count_i0_i3_LC_15_17_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i3_LC_15_17_3 (
            .in0(_gnd_net_),
            .in1(N__39779),
            .in2(_gnd_net_),
            .in3(N__39757),
            .lcout(data_count_3),
            .ltout(),
            .carryin(n19289),
            .carryout(n19290),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__48655),
            .sr(N__48586));
    defparam data_count_i0_i4_LC_15_17_4.C_ON=1'b1;
    defparam data_count_i0_i4_LC_15_17_4.SEQ_MODE=4'b1000;
    defparam data_count_i0_i4_LC_15_17_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i4_LC_15_17_4 (
            .in0(_gnd_net_),
            .in1(N__39671),
            .in2(_gnd_net_),
            .in3(N__39649),
            .lcout(data_count_4),
            .ltout(),
            .carryin(n19290),
            .carryout(n19291),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__48655),
            .sr(N__48586));
    defparam data_count_i0_i5_LC_15_17_5.C_ON=1'b1;
    defparam data_count_i0_i5_LC_15_17_5.SEQ_MODE=4'b1000;
    defparam data_count_i0_i5_LC_15_17_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i5_LC_15_17_5 (
            .in0(_gnd_net_),
            .in1(N__39563),
            .in2(_gnd_net_),
            .in3(N__39541),
            .lcout(data_count_5),
            .ltout(),
            .carryin(n19291),
            .carryout(n19292),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__48655),
            .sr(N__48586));
    defparam data_count_i0_i6_LC_15_17_6.C_ON=1'b1;
    defparam data_count_i0_i6_LC_15_17_6.SEQ_MODE=4'b1000;
    defparam data_count_i0_i6_LC_15_17_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i6_LC_15_17_6 (
            .in0(_gnd_net_),
            .in1(N__39458),
            .in2(_gnd_net_),
            .in3(N__39436),
            .lcout(data_count_6),
            .ltout(),
            .carryin(n19292),
            .carryout(n19293),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__48655),
            .sr(N__48586));
    defparam data_count_i0_i7_LC_15_17_7.C_ON=1'b1;
    defparam data_count_i0_i7_LC_15_17_7.SEQ_MODE=4'b1000;
    defparam data_count_i0_i7_LC_15_17_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i7_LC_15_17_7 (
            .in0(_gnd_net_),
            .in1(N__39356),
            .in2(_gnd_net_),
            .in3(N__39334),
            .lcout(data_count_7),
            .ltout(),
            .carryin(n19293),
            .carryout(n19294),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__48655),
            .sr(N__48586));
    defparam data_count_i0_i8_LC_15_18_0.C_ON=1'b1;
    defparam data_count_i0_i8_LC_15_18_0.SEQ_MODE=4'b1000;
    defparam data_count_i0_i8_LC_15_18_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i8_LC_15_18_0 (
            .in0(_gnd_net_),
            .in1(N__40523),
            .in2(_gnd_net_),
            .in3(N__40501),
            .lcout(data_count_8),
            .ltout(),
            .carryin(bfn_15_18_0_),
            .carryout(n19295),
            .clk(INVdata_count_i0_i8C_net),
            .ce(N__48663),
            .sr(N__48596));
    defparam data_count_i0_i9_LC_15_18_1.C_ON=1'b0;
    defparam data_count_i0_i9_LC_15_18_1.SEQ_MODE=4'b1000;
    defparam data_count_i0_i9_LC_15_18_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i9_LC_15_18_1 (
            .in0(_gnd_net_),
            .in1(N__40412),
            .in2(_gnd_net_),
            .in3(N__40498),
            .lcout(data_count_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVdata_count_i0_i8C_net),
            .ce(N__48663),
            .sr(N__48596));
    defparam \SIG_DDS.tmp_buf_i15_LC_15_19_1 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i15_LC_15_19_1 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i15_LC_15_19_1 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \SIG_DDS.tmp_buf_i15_LC_15_19_1  (
            .in0(N__55872),
            .in1(N__55634),
            .in2(N__40390),
            .in3(N__45591),
            .lcout(tmp_buf_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55221),
            .ce(N__40316),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i0_LC_15_19_7 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i0_LC_15_19_7 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i0_LC_15_19_7 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \SIG_DDS.tmp_buf_i0_LC_15_19_7  (
            .in0(N__55871),
            .in1(N__55633),
            .in2(N__42916),
            .in3(N__40375),
            .lcout(\SIG_DDS.tmp_buf_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55221),
            .ce(N__40316),
            .sr(_gnd_net_));
    defparam \comm_spi.i19199_4_lut_3_lut_LC_16_3_4 .C_ON=1'b0;
    defparam \comm_spi.i19199_4_lut_3_lut_LC_16_3_4 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19199_4_lut_3_lut_LC_16_3_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \comm_spi.i19199_4_lut_3_lut_LC_16_3_4  (
            .in0(N__40229),
            .in1(N__40288),
            .in2(_gnd_net_),
            .in3(N__55472),
            .lcout(\comm_spi.n22623 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i7_12190_12191_set_LC_16_4_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i7_12190_12191_set_LC_16_4_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i7_12190_12191_set_LC_16_4_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i7_12190_12191_set_LC_16_4_0  (
            .in0(N__40230),
            .in1(N__43546),
            .in2(_gnd_net_),
            .in3(N__43641),
            .lcout(\comm_spi.n14592 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52319),
            .ce(),
            .sr(N__40260));
    defparam \comm_spi.data_tx_i7_12190_12191_reset_LC_16_5_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i7_12190_12191_reset_LC_16_5_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i7_12190_12191_reset_LC_16_5_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \comm_spi.data_tx_i7_12190_12191_reset_LC_16_5_0  (
            .in0(N__43645),
            .in1(N__40234),
            .in2(_gnd_net_),
            .in3(N__43545),
            .lcout(\comm_spi.n14593 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52391),
            .ce(),
            .sr(N__44233));
    defparam \comm_spi.imiso_83_12193_12194_reset_LC_16_6_0 .C_ON=1'b0;
    defparam \comm_spi.imiso_83_12193_12194_reset_LC_16_6_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.imiso_83_12193_12194_reset_LC_16_6_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.imiso_83_12193_12194_reset_LC_16_6_0  (
            .in0(N__40209),
            .in1(N__40185),
            .in2(_gnd_net_),
            .in3(N__44283),
            .lcout(\comm_spi.n14596 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.imiso_83_12193_12194_resetC_net ),
            .ce(),
            .sr(N__44232));
    defparam clk_cnt_3761_3762__i2_LC_16_7_0.C_ON=1'b0;
    defparam clk_cnt_3761_3762__i2_LC_16_7_0.SEQ_MODE=4'b1000;
    defparam clk_cnt_3761_3762__i2_LC_16_7_0.LUT_INIT=16'b0101010110101010;
    LogicCell40 clk_cnt_3761_3762__i2_LC_16_7_0 (
            .in0(N__41165),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41189),
            .lcout(clk_cnt_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56024),
            .ce(),
            .sr(N__40723));
    defparam clk_cnt_3761_3762__i1_LC_16_7_1.C_ON=1'b0;
    defparam clk_cnt_3761_3762__i1_LC_16_7_1.SEQ_MODE=4'b1000;
    defparam clk_cnt_3761_3762__i1_LC_16_7_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 clk_cnt_3761_3762__i1_LC_16_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41164),
            .lcout(clk_cnt_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56024),
            .ce(),
            .sr(N__40723));
    defparam i1_4_lut_adj_162_LC_16_8_0.C_ON=1'b0;
    defparam i1_4_lut_adj_162_LC_16_8_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_162_LC_16_8_0.LUT_INIT=16'b1010000010100010;
    LogicCell40 i1_4_lut_adj_162_LC_16_8_0 (
            .in0(N__44418),
            .in1(N__57547),
            .in2(N__40711),
            .in3(N__47833),
            .lcout(comm_state_3_N_412_3),
            .ltout(comm_state_3_N_412_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18743_2_lut_LC_16_8_1.C_ON=1'b0;
    defparam i18743_2_lut_LC_16_8_1.SEQ_MODE=4'b0000;
    defparam i18743_2_lut_LC_16_8_1.LUT_INIT=16'b0101000001010000;
    LogicCell40 i18743_2_lut_LC_16_8_1 (
            .in0(N__53491),
            .in1(_gnd_net_),
            .in2(N__40690),
            .in3(_gnd_net_),
            .lcout(n21162),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15273_2_lut_LC_16_8_2.C_ON=1'b0;
    defparam i15273_2_lut_LC_16_8_2.SEQ_MODE=4'b0000;
    defparam i15273_2_lut_LC_16_8_2.LUT_INIT=16'b1111111110101010;
    LogicCell40 i15273_2_lut_LC_16_8_2 (
            .in0(N__53686),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53489),
            .lcout(n17656),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18105_2_lut_LC_16_8_3.C_ON=1'b0;
    defparam i18105_2_lut_LC_16_8_3.SEQ_MODE=4'b0000;
    defparam i18105_2_lut_LC_16_8_3.LUT_INIT=16'b1000100010001000;
    LogicCell40 i18105_2_lut_LC_16_8_3 (
            .in0(N__53490),
            .in1(N__53685),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(n20700_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_273_LC_16_8_4.C_ON=1'b0;
    defparam i1_4_lut_adj_273_LC_16_8_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_273_LC_16_8_4.LUT_INIT=16'b1010101000000010;
    LogicCell40 i1_4_lut_adj_273_LC_16_8_4 (
            .in0(N__49210),
            .in1(N__51197),
            .in2(N__40687),
            .in3(N__54367),
            .lcout(n11411),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam flagcntwd_303_LC_16_8_5.C_ON=1'b0;
    defparam flagcntwd_303_LC_16_8_5.SEQ_MODE=4'b1000;
    defparam flagcntwd_303_LC_16_8_5.LUT_INIT=16'b1101110111011101;
    LogicCell40 flagcntwd_303_LC_16_8_5 (
            .in0(N__53492),
            .in1(N__53687),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(flagcntwd),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55100),
            .ce(N__40660),
            .sr(N__40648));
    defparam i1_2_lut_adj_249_LC_16_8_6.C_ON=1'b0;
    defparam i1_2_lut_adj_249_LC_16_8_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_249_LC_16_8_6.LUT_INIT=16'b1111111111001100;
    LogicCell40 i1_2_lut_adj_249_LC_16_8_6 (
            .in0(_gnd_net_),
            .in1(N__51196),
            .in2(_gnd_net_),
            .in3(N__53488),
            .lcout(n11333),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i11_4_lut_adj_223_LC_16_9_0.C_ON=1'b0;
    defparam i11_4_lut_adj_223_LC_16_9_0.SEQ_MODE=4'b0000;
    defparam i11_4_lut_adj_223_LC_16_9_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i11_4_lut_adj_223_LC_16_9_0 (
            .in0(N__44487),
            .in1(N__44631),
            .in2(N__44689),
            .in3(N__44539),
            .lcout(n27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15200_2_lut_3_lut_LC_16_9_1.C_ON=1'b0;
    defparam i15200_2_lut_3_lut_LC_16_9_1.SEQ_MODE=4'b0000;
    defparam i15200_2_lut_3_lut_LC_16_9_1.LUT_INIT=16'b0000000001000100;
    LogicCell40 i15200_2_lut_3_lut_LC_16_9_1 (
            .in0(N__53871),
            .in1(N__40784),
            .in2(_gnd_net_),
            .in3(N__51106),
            .lcout(n14_adj_1548),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15201_2_lut_3_lut_LC_16_9_2.C_ON=1'b0;
    defparam i15201_2_lut_3_lut_LC_16_9_2.SEQ_MODE=4'b0000;
    defparam i15201_2_lut_3_lut_LC_16_9_2.LUT_INIT=16'b0000000000100010;
    LogicCell40 i15201_2_lut_3_lut_LC_16_9_2 (
            .in0(N__46700),
            .in1(N__51074),
            .in2(_gnd_net_),
            .in3(N__53872),
            .lcout(n14_adj_1549),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9_4_lut_LC_16_9_3.C_ON=1'b0;
    defparam i9_4_lut_LC_16_9_3.SEQ_MODE=4'b0000;
    defparam i9_4_lut_LC_16_9_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i9_4_lut_LC_16_9_3 (
            .in0(N__44616),
            .in1(N__44454),
            .in2(N__44572),
            .in3(N__44506),
            .lcout(n25_adj_1616),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18268_3_lut_LC_16_9_4.C_ON=1'b0;
    defparam i18268_3_lut_LC_16_9_4.SEQ_MODE=4'b0000;
    defparam i18268_3_lut_LC_16_9_4.LUT_INIT=16'b1110111001010101;
    LogicCell40 i18268_3_lut_LC_16_9_4 (
            .in0(N__53494),
            .in1(N__49790),
            .in2(_gnd_net_),
            .in3(N__53873),
            .lcout(n20863),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_LC_16_9_5.C_ON=1'b0;
    defparam i2_2_lut_LC_16_9_5.SEQ_MODE=4'b0000;
    defparam i2_2_lut_LC_16_9_5.LUT_INIT=16'b1010101011111111;
    LogicCell40 i2_2_lut_LC_16_9_5 (
            .in0(N__49791),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53493),
            .lcout(n14514),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_73_LC_16_9_6.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_73_LC_16_9_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_73_LC_16_9_6.LUT_INIT=16'b1010101010001000;
    LogicCell40 i1_2_lut_3_lut_adj_73_LC_16_9_6 (
            .in0(N__49211),
            .in1(N__54372),
            .in2(_gnd_net_),
            .in3(N__51073),
            .lcout(n20556),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12_4_lut_adj_221_LC_16_9_7.C_ON=1'b0;
    defparam i12_4_lut_adj_221_LC_16_9_7.SEQ_MODE=4'b0000;
    defparam i12_4_lut_adj_221_LC_16_9_7.LUT_INIT=16'b1111111111111110;
    LogicCell40 i12_4_lut_adj_221_LC_16_9_7 (
            .in0(N__44586),
            .in1(N__44953),
            .in2(N__44671),
            .in3(N__44520),
            .lcout(n28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10_4_lut_adj_222_LC_16_10_0.C_ON=1'b0;
    defparam i10_4_lut_adj_222_LC_16_10_0.SEQ_MODE=4'b0000;
    defparam i10_4_lut_adj_222_LC_16_10_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i10_4_lut_adj_222_LC_16_10_0 (
            .in0(N__44553),
            .in1(N__44601),
            .in2(N__44650),
            .in3(N__44473),
            .lcout(),
            .ltout(n26_adj_1625_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15_4_lut_adj_227_LC_16_10_1.C_ON=1'b0;
    defparam i15_4_lut_adj_227_LC_16_10_1.SEQ_MODE=4'b0000;
    defparam i15_4_lut_adj_227_LC_16_10_1.LUT_INIT=16'b1111111111111110;
    LogicCell40 i15_4_lut_adj_227_LC_16_10_1 (
            .in0(N__40747),
            .in1(N__40741),
            .in2(N__40735),
            .in3(N__40732),
            .lcout(),
            .ltout(n19553_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7_4_lut_adj_228_LC_16_10_2.C_ON=1'b0;
    defparam i7_4_lut_adj_228_LC_16_10_2.SEQ_MODE=4'b0000;
    defparam i7_4_lut_adj_228_LC_16_10_2.LUT_INIT=16'b0000100000000000;
    LogicCell40 i7_4_lut_adj_228_LC_16_10_2 (
            .in0(N__44931),
            .in1(N__53038),
            .in2(N__40726),
            .in3(N__41203),
            .lcout(n14700),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12387_3_lut_LC_16_10_3.C_ON=1'b0;
    defparam i12387_3_lut_LC_16_10_3.SEQ_MODE=4'b0000;
    defparam i12387_3_lut_LC_16_10_3.LUT_INIT=16'b1000100010101010;
    LogicCell40 i12387_3_lut_LC_16_10_3 (
            .in0(N__47081),
            .in1(N__54537),
            .in2(_gnd_net_),
            .in3(N__49302),
            .lcout(n14784),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_6_i22_3_lut_LC_16_10_4.C_ON=1'b0;
    defparam mux_130_Mux_6_i22_3_lut_LC_16_10_4.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_6_i22_3_lut_LC_16_10_4.LUT_INIT=16'b1100110010101010;
    LogicCell40 mux_130_Mux_6_i22_3_lut_LC_16_10_4 (
            .in0(N__48564),
            .in1(N__40831),
            .in2(_gnd_net_),
            .in3(N__47832),
            .lcout(n22_adj_1594),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_adj_225_LC_16_10_7.C_ON=1'b0;
    defparam i2_2_lut_adj_225_LC_16_10_7.SEQ_MODE=4'b0000;
    defparam i2_2_lut_adj_225_LC_16_10_7.LUT_INIT=16'b1010101000000000;
    LogicCell40 i2_2_lut_adj_225_LC_16_10_7 (
            .in0(N__44703),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44967),
            .lcout(n10_adj_1582),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_RTD_287_LC_16_11_0.C_ON=1'b0;
    defparam clk_RTD_287_LC_16_11_0.SEQ_MODE=4'b1000;
    defparam clk_RTD_287_LC_16_11_0.LUT_INIT=16'b0110011010101010;
    LogicCell40 clk_RTD_287_LC_16_11_0 (
            .in0(N__40961),
            .in1(N__41196),
            .in2(_gnd_net_),
            .in3(N__41170),
            .lcout(clk_RTD),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56026),
            .ce(),
            .sr(_gnd_net_));
    defparam SecClk_292_LC_16_11_1.C_ON=1'b0;
    defparam SecClk_292_LC_16_11_1.SEQ_MODE=4'b1000;
    defparam SecClk_292_LC_16_11_1.LUT_INIT=16'b0011001111001100;
    LogicCell40 SecClk_292_LC_16_11_1 (
            .in0(_gnd_net_),
            .in1(N__40906),
            .in2(_gnd_net_),
            .in3(N__44902),
            .lcout(TEST_LED),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56026),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_6_i19_3_lut_LC_16_11_2.C_ON=1'b0;
    defparam mux_130_Mux_6_i19_3_lut_LC_16_11_2.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_6_i19_3_lut_LC_16_11_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_130_Mux_6_i19_3_lut_LC_16_11_2 (
            .in0(N__40888),
            .in1(N__40860),
            .in2(_gnd_net_),
            .in3(N__56939),
            .lcout(n19_adj_1593),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i45_4_lut_LC_16_11_3.C_ON=1'b0;
    defparam i45_4_lut_LC_16_11_3.SEQ_MODE=4'b0000;
    defparam i45_4_lut_LC_16_11_3.LUT_INIT=16'b1110110000100000;
    LogicCell40 i45_4_lut_LC_16_11_3 (
            .in0(N__44411),
            .in1(N__53837),
            .in2(N__40825),
            .in3(N__46996),
            .lcout(n20_adj_1607),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_3_lut_LC_16_11_5.C_ON=1'b0;
    defparam i2_2_lut_3_lut_LC_16_11_5.SEQ_MODE=4'b0000;
    defparam i2_2_lut_3_lut_LC_16_11_5.LUT_INIT=16'b1011101111111111;
    LogicCell40 i2_2_lut_3_lut_LC_16_11_5 (
            .in0(N__56940),
            .in1(N__57543),
            .in2(_gnd_net_),
            .in3(N__47754),
            .lcout(n10553),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_137_Mux_4_i4_3_lut_LC_16_11_6.C_ON=1'b0;
    defparam mux_137_Mux_4_i4_3_lut_LC_16_11_6.SEQ_MODE=4'b0000;
    defparam mux_137_Mux_4_i4_3_lut_LC_16_11_6.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_137_Mux_4_i4_3_lut_LC_16_11_6 (
            .in0(N__40804),
            .in1(N__51579),
            .in2(_gnd_net_),
            .in3(N__40795),
            .lcout(n4_adj_1566),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18184_3_lut_LC_16_11_7.C_ON=1'b0;
    defparam i18184_3_lut_LC_16_11_7.SEQ_MODE=4'b0000;
    defparam i18184_3_lut_LC_16_11_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 i18184_3_lut_LC_16_11_7 (
            .in0(N__56938),
            .in1(N__41469),
            .in2(_gnd_net_),
            .in3(N__47343),
            .lcout(n20779),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_57_LC_16_12_0.C_ON=1'b0;
    defparam i1_4_lut_adj_57_LC_16_12_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_57_LC_16_12_0.LUT_INIT=16'b1100000011010000;
    LogicCell40 i1_4_lut_adj_57_LC_16_12_0 (
            .in0(N__45562),
            .in1(N__52063),
            .in2(N__54669),
            .in3(N__41615),
            .lcout(n12415),
            .ltout(n12415_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i6_LC_16_12_1.C_ON=1'b0;
    defparam req_data_cnt_i6_LC_16_12_1.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i6_LC_16_12_1.LUT_INIT=16'b1010111110100000;
    LogicCell40 req_data_cnt_i6_LC_16_12_1 (
            .in0(N__51376),
            .in1(_gnd_net_),
            .in2(N__41440),
            .in3(N__41718),
            .lcout(req_data_cnt_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55142),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i5_LC_16_12_2.C_ON=1'b0;
    defparam buf_cfgRTD_i5_LC_16_12_2.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i5_LC_16_12_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 buf_cfgRTD_i5_LC_16_12_2 (
            .in0(N__45292),
            .in1(N__44800),
            .in2(_gnd_net_),
            .in3(N__41386),
            .lcout(buf_cfgRTD_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55142),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i13_LC_16_12_3.C_ON=1'b0;
    defparam req_data_cnt_i13_LC_16_12_3.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i13_LC_16_12_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 req_data_cnt_i13_LC_16_12_3 (
            .in0(N__44799),
            .in1(N__41987),
            .in2(_gnd_net_),
            .in3(N__45087),
            .lcout(req_data_cnt_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55142),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i0_LC_16_12_4.C_ON=1'b0;
    defparam req_data_cnt_i0_LC_16_12_4.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i0_LC_16_12_4.LUT_INIT=16'b0111010100100000;
    LogicCell40 req_data_cnt_i0_LC_16_12_4 (
            .in0(N__41990),
            .in1(N__52064),
            .in2(N__41363),
            .in3(N__41744),
            .lcout(req_data_cnt_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55142),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i2_LC_16_12_5.C_ON=1'b0;
    defparam req_data_cnt_i2_LC_16_12_5.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i2_LC_16_12_5.LUT_INIT=16'b1011101110001000;
    LogicCell40 req_data_cnt_i2_LC_16_12_5 (
            .in0(N__41284),
            .in1(N__41988),
            .in2(_gnd_net_),
            .in3(N__41591),
            .lcout(req_data_cnt_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55142),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i7_LC_16_12_6.C_ON=1'b0;
    defparam req_data_cnt_i7_LC_16_12_6.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i7_LC_16_12_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 req_data_cnt_i7_LC_16_12_6 (
            .in0(N__41989),
            .in1(N__41263),
            .in2(_gnd_net_),
            .in3(N__41565),
            .lcout(req_data_cnt_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55142),
            .ce(),
            .sr(_gnd_net_));
    defparam i1536244_i1_3_lut_LC_16_12_7.C_ON=1'b0;
    defparam i1536244_i1_3_lut_LC_16_12_7.SEQ_MODE=4'b0000;
    defparam i1536244_i1_3_lut_LC_16_12_7.LUT_INIT=16'b1010101011001100;
    LogicCell40 i1536244_i1_3_lut_LC_16_12_7 (
            .in0(N__45028),
            .in1(N__41242),
            .in2(_gnd_net_),
            .in3(N__56315),
            .lcout(n30_adj_1520),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i11_LC_16_13_1.C_ON=1'b0;
    defparam req_data_cnt_i11_LC_16_13_1.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i11_LC_16_13_1.LUT_INIT=16'b0101110100001000;
    LogicCell40 req_data_cnt_i11_LC_16_13_1 (
            .in0(N__41992),
            .in1(N__43802),
            .in2(N__52158),
            .in3(N__45255),
            .lcout(req_data_cnt_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55155),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i8_LC_16_13_2.C_ON=1'b0;
    defparam req_data_cnt_i8_LC_16_13_2.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i8_LC_16_13_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 req_data_cnt_i8_LC_16_13_2 (
            .in0(N__41782),
            .in1(N__41991),
            .in2(_gnd_net_),
            .in3(N__41895),
            .lcout(req_data_cnt_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55155),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_74_LC_16_13_3.C_ON=1'b0;
    defparam i1_4_lut_adj_74_LC_16_13_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_74_LC_16_13_3.LUT_INIT=16'b0111101111011110;
    LogicCell40 i1_4_lut_adj_74_LC_16_13_3 (
            .in0(N__46936),
            .in1(N__47412),
            .in2(N__41751),
            .in3(N__41714),
            .lcout(n17_adj_1554),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i8_4_lut_adj_55_LC_16_13_4.C_ON=1'b0;
    defparam i8_4_lut_adj_55_LC_16_13_4.SEQ_MODE=4'b0000;
    defparam i8_4_lut_adj_55_LC_16_13_4.LUT_INIT=16'b0111101111011110;
    LogicCell40 i8_4_lut_adj_55_LC_16_13_4 (
            .in0(N__48682),
            .in1(N__47307),
            .in2(N__41691),
            .in3(N__41642),
            .lcout(n24_adj_1530),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_4_lut_LC_16_13_5.C_ON=1'b0;
    defparam i1_2_lut_4_lut_LC_16_13_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_4_lut_LC_16_13_5.LUT_INIT=16'b1111111110111111;
    LogicCell40 i1_2_lut_4_lut_LC_16_13_5 (
            .in0(N__56803),
            .in1(N__47790),
            .in2(N__57533),
            .in3(N__41614),
            .lcout(n10540),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6_4_lut_adj_56_LC_16_13_6.C_ON=1'b0;
    defparam i6_4_lut_adj_56_LC_16_13_6.SEQ_MODE=4'b0000;
    defparam i6_4_lut_adj_56_LC_16_13_6.LUT_INIT=16'b0111101111011110;
    LogicCell40 i6_4_lut_adj_56_LC_16_13_6 (
            .in0(N__46881),
            .in1(N__47377),
            .in2(N__41592),
            .in3(N__41561),
            .lcout(n22_adj_1492),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_adj_313_LC_16_14_0.C_ON=1'b0;
    defparam i2_3_lut_adj_313_LC_16_14_0.SEQ_MODE=4'b0000;
    defparam i2_3_lut_adj_313_LC_16_14_0.LUT_INIT=16'b1111111110111011;
    LogicCell40 i2_3_lut_adj_313_LC_16_14_0 (
            .in0(N__51659),
            .in1(N__51200),
            .in2(_gnd_net_),
            .in3(N__53956),
            .lcout(n10579),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i14_LC_16_14_1.C_ON=1'b0;
    defparam req_data_cnt_i14_LC_16_14_1.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i14_LC_16_14_1.LUT_INIT=16'b1011101110001000;
    LogicCell40 req_data_cnt_i14_LC_16_14_1 (
            .in0(N__41506),
            .in1(N__42008),
            .in2(_gnd_net_),
            .in3(N__45231),
            .lcout(req_data_cnt_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55170),
            .ce(),
            .sr(_gnd_net_));
    defparam i5_4_lut_adj_59_LC_16_14_2.C_ON=1'b0;
    defparam i5_4_lut_adj_59_LC_16_14_2.SEQ_MODE=4'b0000;
    defparam i5_4_lut_adj_59_LC_16_14_2.LUT_INIT=16'b0111110110111110;
    LogicCell40 i5_4_lut_adj_59_LC_16_14_2 (
            .in0(N__47221),
            .in1(N__41912),
            .in2(N__47278),
            .in3(N__56387),
            .lcout(),
            .ltout(n21_adj_1494_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i14_4_lut_adj_79_LC_16_14_3.C_ON=1'b0;
    defparam i14_4_lut_adj_79_LC_16_14_3.SEQ_MODE=4'b0000;
    defparam i14_4_lut_adj_79_LC_16_14_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i14_4_lut_adj_79_LC_16_14_3 (
            .in0(N__42169),
            .in1(N__45211),
            .in2(N__42160),
            .in3(N__42157),
            .lcout(n30_adj_1597),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i4_LC_16_14_4.C_ON=1'b0;
    defparam buf_cfgRTD_i4_LC_16_14_4.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i4_LC_16_14_4.LUT_INIT=16'b1011101110001000;
    LogicCell40 buf_cfgRTD_i4_LC_16_14_4 (
            .in0(N__42119),
            .in1(N__45279),
            .in2(_gnd_net_),
            .in3(N__42044),
            .lcout(buf_cfgRTD_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55170),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i10_LC_16_14_5.C_ON=1'b0;
    defparam req_data_cnt_i10_LC_16_14_5.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i10_LC_16_14_5.LUT_INIT=16'b1110111000100010;
    LogicCell40 req_data_cnt_i10_LC_16_14_5 (
            .in0(N__41913),
            .in1(N__42007),
            .in2(_gnd_net_),
            .in3(N__41950),
            .lcout(req_data_cnt_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55170),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_4_lut_LC_16_14_6.C_ON=1'b0;
    defparam i3_4_lut_LC_16_14_6.SEQ_MODE=4'b0000;
    defparam i3_4_lut_LC_16_14_6.LUT_INIT=16'b0111101111011110;
    LogicCell40 i3_4_lut_LC_16_14_6 (
            .in0(N__47200),
            .in1(N__47344),
            .in2(N__45091),
            .in3(N__41891),
            .lcout(n19_adj_1499),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_125_2_lut_LC_16_15_0.C_ON=1'b1;
    defparam add_125_2_lut_LC_16_15_0.SEQ_MODE=4'b0000;
    defparam add_125_2_lut_LC_16_15_0.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_125_2_lut_LC_16_15_0 (
            .in0(N__42841),
            .in1(N__42839),
            .in2(N__42339),
            .in3(N__41869),
            .lcout(n7_adj_1515),
            .ltout(),
            .carryin(bfn_16_15_0_),
            .carryout(n19326),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_125_3_lut_LC_16_15_1.C_ON=1'b1;
    defparam add_125_3_lut_LC_16_15_1.SEQ_MODE=4'b0000;
    defparam add_125_3_lut_LC_16_15_1.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_125_3_lut_LC_16_15_1 (
            .in0(N__43321),
            .in1(N__43320),
            .in2(N__42343),
            .in3(N__41866),
            .lcout(n7_adj_1546),
            .ltout(),
            .carryin(n19326),
            .carryout(n19327),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_125_4_lut_LC_16_15_2.C_ON=1'b1;
    defparam add_125_4_lut_LC_16_15_2.SEQ_MODE=4'b0000;
    defparam add_125_4_lut_LC_16_15_2.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_125_4_lut_LC_16_15_2 (
            .in0(N__41863),
            .in1(N__41862),
            .in2(N__42340),
            .in3(N__41830),
            .lcout(n7_adj_1544),
            .ltout(),
            .carryin(n19327),
            .carryout(n19328),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_125_5_lut_LC_16_15_3.C_ON=1'b1;
    defparam add_125_5_lut_LC_16_15_3.SEQ_MODE=4'b0000;
    defparam add_125_5_lut_LC_16_15_3.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_125_5_lut_LC_16_15_3 (
            .in0(N__41826),
            .in1(N__41825),
            .in2(N__42344),
            .in3(N__41785),
            .lcout(n7_adj_1542),
            .ltout(),
            .carryin(n19328),
            .carryout(n19329),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_125_6_lut_LC_16_15_4.C_ON=1'b1;
    defparam add_125_6_lut_LC_16_15_4.SEQ_MODE=4'b0000;
    defparam add_125_6_lut_LC_16_15_4.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_125_6_lut_LC_16_15_4 (
            .in0(N__42507),
            .in1(N__42506),
            .in2(N__42341),
            .in3(N__42481),
            .lcout(n7_adj_1540),
            .ltout(),
            .carryin(n19329),
            .carryout(n19330),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_125_7_lut_LC_16_15_5.C_ON=1'b1;
    defparam add_125_7_lut_LC_16_15_5.SEQ_MODE=4'b0000;
    defparam add_125_7_lut_LC_16_15_5.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_125_7_lut_LC_16_15_5 (
            .in0(N__46038),
            .in1(N__46037),
            .in2(N__42345),
            .in3(N__42478),
            .lcout(n17336),
            .ltout(),
            .carryin(n19330),
            .carryout(n19331),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_125_8_lut_LC_16_15_6.C_ON=1'b1;
    defparam add_125_8_lut_LC_16_15_6.SEQ_MODE=4'b0000;
    defparam add_125_8_lut_LC_16_15_6.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_125_8_lut_LC_16_15_6 (
            .in0(N__42679),
            .in1(N__42678),
            .in2(N__42342),
            .in3(N__42475),
            .lcout(n7_adj_1537),
            .ltout(),
            .carryin(n19331),
            .carryout(n19332),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_125_9_lut_LC_16_15_7.C_ON=1'b1;
    defparam add_125_9_lut_LC_16_15_7.SEQ_MODE=4'b0000;
    defparam add_125_9_lut_LC_16_15_7.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_125_9_lut_LC_16_15_7 (
            .in0(N__42472),
            .in1(N__42471),
            .in2(N__42346),
            .in3(N__42412),
            .lcout(n7_adj_1535),
            .ltout(),
            .carryin(n19332),
            .carryout(n19333),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_125_10_lut_LC_16_16_0.C_ON=1'b1;
    defparam add_125_10_lut_LC_16_16_0.SEQ_MODE=4'b0000;
    defparam add_125_10_lut_LC_16_16_0.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_125_10_lut_LC_16_16_0 (
            .in0(N__42409),
            .in1(N__42408),
            .in2(N__42358),
            .in3(N__42361),
            .lcout(n7_adj_1533),
            .ltout(),
            .carryin(bfn_16_16_0_),
            .carryout(n19334),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_125_11_lut_LC_16_16_1.C_ON=1'b0;
    defparam add_125_11_lut_LC_16_16_1.SEQ_MODE=4'b0000;
    defparam add_125_11_lut_LC_16_16_1.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_125_11_lut_LC_16_16_1 (
            .in0(N__42725),
            .in1(N__42726),
            .in2(N__42357),
            .in3(N__42268),
            .lcout(n7_adj_1531),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i9_LC_16_16_2.C_ON=1'b0;
    defparam data_index_i9_LC_16_16_2.SEQ_MODE=4'b1000;
    defparam data_index_i9_LC_16_16_2.LUT_INIT=16'b0101110100001000;
    LogicCell40 data_index_i9_LC_16_16_2 (
            .in0(N__54635),
            .in1(N__43038),
            .in2(N__52033),
            .in3(N__43023),
            .lcout(data_index_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55199),
            .ce(),
            .sr(_gnd_net_));
    defparam i14955_3_lut_LC_16_16_3.C_ON=1'b0;
    defparam i14955_3_lut_LC_16_16_3.SEQ_MODE=4'b0000;
    defparam i14955_3_lut_LC_16_16_3.LUT_INIT=16'b1100110010101010;
    LogicCell40 i14955_3_lut_LC_16_16_3 (
            .in0(N__50183),
            .in1(N__46042),
            .in2(_gnd_net_),
            .in3(N__43275),
            .lcout(n17338),
            .ltout(n17338_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i14957_4_lut_LC_16_16_4.C_ON=1'b0;
    defparam i14957_4_lut_LC_16_16_4.SEQ_MODE=4'b0000;
    defparam i14957_4_lut_LC_16_16_4.LUT_INIT=16'b0111001101000000;
    LogicCell40 i14957_4_lut_LC_16_16_4 (
            .in0(N__51920),
            .in1(N__54610),
            .in2(N__42265),
            .in3(N__46053),
            .lcout(data_index_9_N_212_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i0_LC_16_16_5.C_ON=1'b0;
    defparam data_index_i0_LC_16_16_5.SEQ_MODE=4'b1000;
    defparam data_index_i0_LC_16_16_5.LUT_INIT=16'b0100111001000100;
    LogicCell40 data_index_i0_LC_16_16_5 (
            .in0(N__54611),
            .in1(N__42873),
            .in2(N__52077),
            .in3(N__42855),
            .lcout(data_index_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55199),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i2_LC_16_16_6.C_ON=1'b0;
    defparam buf_dds0_i2_LC_16_16_6.SEQ_MODE=4'b1000;
    defparam buf_dds0_i2_LC_16_16_6.LUT_INIT=16'b0111010100100000;
    LogicCell40 buf_dds0_i2_LC_16_16_6 (
            .in0(N__45697),
            .in1(N__51979),
            .in2(N__42822),
            .in3(N__42746),
            .lcout(buf_dds0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55199),
            .ce(),
            .sr(_gnd_net_));
    defparam i6352_3_lut_LC_16_16_7.C_ON=1'b0;
    defparam i6352_3_lut_LC_16_16_7.SEQ_MODE=4'b0000;
    defparam i6352_3_lut_LC_16_16_7.LUT_INIT=16'b1100110010101010;
    LogicCell40 i6352_3_lut_LC_16_16_7 (
            .in0(N__44107),
            .in1(N__42727),
            .in2(_gnd_net_),
            .in3(N__43274),
            .lcout(n8_adj_1532),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i4_LC_16_17_0.C_ON=1'b0;
    defparam buf_dds0_i4_LC_16_17_0.SEQ_MODE=4'b1000;
    defparam buf_dds0_i4_LC_16_17_0.LUT_INIT=16'b0101000011001100;
    LogicCell40 buf_dds0_i4_LC_16_17_0 (
            .in0(N__51975),
            .in1(N__42701),
            .in2(N__46665),
            .in3(N__45675),
            .lcout(buf_dds0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55212),
            .ce(),
            .sr(_gnd_net_));
    defparam i6382_3_lut_LC_16_17_1.C_ON=1'b0;
    defparam i6382_3_lut_LC_16_17_1.SEQ_MODE=4'b0000;
    defparam i6382_3_lut_LC_16_17_1.LUT_INIT=16'b1100110010101010;
    LogicCell40 i6382_3_lut_LC_16_17_1 (
            .in0(N__51431),
            .in1(N__42677),
            .in2(_gnd_net_),
            .in3(N__43276),
            .lcout(n8_adj_1538),
            .ltout(n8_adj_1538_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i6_LC_16_17_2.C_ON=1'b0;
    defparam data_index_i6_LC_16_17_2.SEQ_MODE=4'b1000;
    defparam data_index_i6_LC_16_17_2.LUT_INIT=16'b0111001101000000;
    LogicCell40 data_index_i6_LC_16_17_2 (
            .in0(N__51976),
            .in1(N__54705),
            .in2(N__42682),
            .in3(N__43981),
            .lcout(data_index_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55212),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i6_LC_16_17_3.C_ON=1'b0;
    defparam buf_dds0_i6_LC_16_17_3.SEQ_MODE=4'b1000;
    defparam buf_dds0_i6_LC_16_17_3.LUT_INIT=16'b0111010100100000;
    LogicCell40 buf_dds0_i6_LC_16_17_3 (
            .in0(N__45676),
            .in1(N__51977),
            .in2(N__51438),
            .in3(N__42644),
            .lcout(buf_dds0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55212),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i7_LC_16_17_4.C_ON=1'b0;
    defparam buf_dds1_i7_LC_16_17_4.SEQ_MODE=4'b1000;
    defparam buf_dds1_i7_LC_16_17_4.LUT_INIT=16'b1010000010001000;
    LogicCell40 buf_dds1_i7_LC_16_17_4 (
            .in0(N__45965),
            .in1(N__42530),
            .in2(N__42625),
            .in3(N__45829),
            .lcout(buf_dds1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55212),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i0_LC_16_17_6.C_ON=1'b0;
    defparam buf_control_i0_LC_16_17_6.SEQ_MODE=4'b1000;
    defparam buf_control_i0_LC_16_17_6.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_control_i0_LC_16_17_6 (
            .in0(N__51974),
            .in1(N__43865),
            .in2(N__43532),
            .in3(N__50285),
            .lcout(buf_control_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55212),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i1_LC_16_18_1.C_ON=1'b0;
    defparam data_index_i1_LC_16_18_1.SEQ_MODE=4'b1000;
    defparam data_index_i1_LC_16_18_1.LUT_INIT=16'b0101110100001000;
    LogicCell40 data_index_i1_LC_16_18_1 (
            .in0(N__54704),
            .in1(N__43228),
            .in2(N__52043),
            .in3(N__43219),
            .lcout(data_index_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55222),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i8_LC_16_18_3.C_ON=1'b0;
    defparam buf_dds0_i8_LC_16_18_3.SEQ_MODE=4'b1000;
    defparam buf_dds0_i8_LC_16_18_3.LUT_INIT=16'b0101110100001000;
    LogicCell40 buf_dds0_i8_LC_16_18_3 (
            .in0(N__45696),
            .in1(N__43524),
            .in2(N__52042),
            .in3(N__43409),
            .lcout(buf_dds0_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55222),
            .ce(),
            .sr(_gnd_net_));
    defparam i6432_3_lut_LC_16_18_4.C_ON=1'b0;
    defparam i6432_3_lut_LC_16_18_4.SEQ_MODE=4'b0000;
    defparam i6432_3_lut_LC_16_18_4.LUT_INIT=16'b1100110010101010;
    LogicCell40 i6432_3_lut_LC_16_18_4 (
            .in0(N__43375),
            .in1(N__43319),
            .in2(_gnd_net_),
            .in3(N__43291),
            .lcout(n8_adj_1547),
            .ltout(n8_adj_1547_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_354_Mux_1_i15_4_lut_LC_16_18_5.C_ON=1'b0;
    defparam comm_state_3__I_0_354_Mux_1_i15_4_lut_LC_16_18_5.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_354_Mux_1_i15_4_lut_LC_16_18_5.LUT_INIT=16'b0111001101000000;
    LogicCell40 comm_state_3__I_0_354_Mux_1_i15_4_lut_LC_16_18_5 (
            .in0(N__51929),
            .in1(N__54597),
            .in2(N__43222),
            .in3(N__43218),
            .lcout(data_index_9_N_212_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i11_LC_16_18_6.C_ON=1'b0;
    defparam buf_dds0_i11_LC_16_18_6.SEQ_MODE=4'b1000;
    defparam buf_dds0_i11_LC_16_18_6.LUT_INIT=16'b0011000010111000;
    LogicCell40 buf_dds0_i11_LC_16_18_6 (
            .in0(N__43821),
            .in1(N__45694),
            .in2(N__43097),
            .in3(N__51930),
            .lcout(buf_dds0_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55222),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i5_LC_16_18_7.C_ON=1'b0;
    defparam buf_dds0_i5_LC_16_18_7.SEQ_MODE=4'b1000;
    defparam buf_dds0_i5_LC_16_18_7.LUT_INIT=16'b0111010100100000;
    LogicCell40 buf_dds0_i5_LC_16_18_7 (
            .in0(N__45695),
            .in1(N__51983),
            .in2(N__50190),
            .in3(N__43055),
            .lcout(buf_dds0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55222),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_354_Mux_9_i15_4_lut_LC_16_19_0.C_ON=1'b0;
    defparam comm_state_3__I_0_354_Mux_9_i15_4_lut_LC_16_19_0.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_354_Mux_9_i15_4_lut_LC_16_19_0.LUT_INIT=16'b0101110100001000;
    LogicCell40 comm_state_3__I_0_354_Mux_9_i15_4_lut_LC_16_19_0 (
            .in0(N__54703),
            .in1(N__43039),
            .in2(N__52124),
            .in3(N__43024),
            .lcout(data_index_9_N_212_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.MOSI_31_LC_16_19_2 .C_ON=1'b0;
    defparam \SIG_DDS.MOSI_31_LC_16_19_2 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.MOSI_31_LC_16_19_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \SIG_DDS.MOSI_31_LC_16_19_2  (
            .in0(N__42915),
            .in1(N__42885),
            .in2(_gnd_net_),
            .in3(N__55566),
            .lcout(DDS_MOSI),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55231),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i1_LC_16_19_3.C_ON=1'b0;
    defparam buf_control_i1_LC_16_19_3.SEQ_MODE=4'b1000;
    defparam buf_control_i1_LC_16_19_3.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_control_i1_LC_16_19_3 (
            .in0(N__52059),
            .in1(N__43872),
            .in2(N__44147),
            .in3(N__44009),
            .lcout(DDS_RNG_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55231),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_354_Mux_6_i15_4_lut_LC_16_19_4.C_ON=1'b0;
    defparam comm_state_3__I_0_354_Mux_6_i15_4_lut_LC_16_19_4.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_354_Mux_6_i15_4_lut_LC_16_19_4.LUT_INIT=16'b0101110100001000;
    LogicCell40 comm_state_3__I_0_354_Mux_6_i15_4_lut_LC_16_19_4 (
            .in0(N__54702),
            .in1(N__43990),
            .in2(N__52123),
            .in3(N__43980),
            .lcout(data_index_9_N_212_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i3_LC_16_19_5.C_ON=1'b0;
    defparam buf_control_i3_LC_16_19_5.SEQ_MODE=4'b1000;
    defparam buf_control_i3_LC_16_19_5.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_control_i3_LC_16_19_5 (
            .in0(N__52060),
            .in1(N__43873),
            .in2(N__43822),
            .in3(N__45497),
            .lcout(SELIRNG1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55231),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.bit_cnt_i0_LC_16_19_7 .C_ON=1'b0;
    defparam \SIG_DDS.bit_cnt_i0_LC_16_19_7 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.bit_cnt_i0_LC_16_19_7 .LUT_INIT=16'b0000000001011010;
    LogicCell40 \SIG_DDS.bit_cnt_i0_LC_16_19_7  (
            .in0(N__55567),
            .in1(_gnd_net_),
            .in2(N__43673),
            .in3(N__43710),
            .lcout(bit_cnt_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55231),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i6_12221_12222_reset_LC_17_3_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i6_12221_12222_reset_LC_17_3_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i6_12221_12222_reset_LC_17_3_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i6_12221_12222_reset_LC_17_3_0  (
            .in0(N__43573),
            .in1(N__46246),
            .in2(_gnd_net_),
            .in3(N__46293),
            .lcout(\comm_spi.n14624 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52416),
            .ce(),
            .sr(N__43630));
    defparam \comm_spi.i19154_4_lut_3_lut_LC_17_4_3 .C_ON=1'b0;
    defparam \comm_spi.i19154_4_lut_3_lut_LC_17_4_3 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19154_4_lut_3_lut_LC_17_4_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.i19154_4_lut_3_lut_LC_17_4_3  (
            .in0(N__52960),
            .in1(N__43612),
            .in2(_gnd_net_),
            .in3(N__55428),
            .lcout(\comm_spi.n22626 ),
            .ltout(\comm_spi.n22626_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i12181_3_lut_LC_17_4_4 .C_ON=1'b0;
    defparam \comm_spi.i12181_3_lut_LC_17_4_4 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i12181_3_lut_LC_17_4_4 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \comm_spi.i12181_3_lut_LC_17_4_4  (
            .in0(_gnd_net_),
            .in1(N__52969),
            .in2(N__43606),
            .in3(N__48769),
            .lcout(\comm_spi.iclk ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i12189_3_lut_LC_17_4_6 .C_ON=1'b0;
    defparam \comm_spi.i12189_3_lut_LC_17_4_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i12189_3_lut_LC_17_4_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \comm_spi.i12189_3_lut_LC_17_4_6  (
            .in0(N__44287),
            .in1(N__44242),
            .in2(_gnd_net_),
            .in3(N__43603),
            .lcout(ICE_SPI_MISO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i6_12221_12222_set_LC_17_5_4 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i6_12221_12222_set_LC_17_5_4 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i6_12221_12222_set_LC_17_5_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i6_12221_12222_set_LC_17_5_4  (
            .in0(N__43569),
            .in1(N__46242),
            .in2(_gnd_net_),
            .in3(N__46294),
            .lcout(\comm_spi.n14623 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52379),
            .ce(),
            .sr(N__44341));
    defparam \comm_spi.MISO_48_12187_12188_reset_LC_17_6_0 .C_ON=1'b0;
    defparam \comm_spi.MISO_48_12187_12188_reset_LC_17_6_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.MISO_48_12187_12188_reset_LC_17_6_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \comm_spi.MISO_48_12187_12188_reset_LC_17_6_0  (
            .in0(N__44322),
            .in1(N__44311),
            .in2(_gnd_net_),
            .in3(N__44282),
            .lcout(\comm_spi.n14590 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.MISO_48_12187_12188_resetC_net ),
            .ce(),
            .sr(N__44231));
    defparam comm_state_i1_LC_17_7_0.C_ON=1'b0;
    defparam comm_state_i1_LC_17_7_0.SEQ_MODE=4'b1000;
    defparam comm_state_i1_LC_17_7_0.LUT_INIT=16'b0101110100001000;
    LogicCell40 comm_state_i1_LC_17_7_0 (
            .in0(N__54249),
            .in1(N__44428),
            .in2(N__52113),
            .in3(N__44179),
            .lcout(comm_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55101),
            .ce(N__44161),
            .sr(_gnd_net_));
    defparam comm_state_1__bdd_4_lut_LC_17_7_1.C_ON=1'b0;
    defparam comm_state_1__bdd_4_lut_LC_17_7_1.SEQ_MODE=4'b0000;
    defparam comm_state_1__bdd_4_lut_LC_17_7_1.LUT_INIT=16'b1110010010101010;
    LogicCell40 comm_state_1__bdd_4_lut_LC_17_7_1 (
            .in0(N__53681),
            .in1(N__44197),
            .in2(N__52232),
            .in3(N__51110),
            .lcout(),
            .ltout(n21913_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n21913_bdd_4_lut_LC_17_7_2.C_ON=1'b0;
    defparam n21913_bdd_4_lut_LC_17_7_2.SEQ_MODE=4'b0000;
    defparam n21913_bdd_4_lut_LC_17_7_2.LUT_INIT=16'b1111010010100100;
    LogicCell40 n21913_bdd_4_lut_LC_17_7_2 (
            .in0(N__51111),
            .in1(N__53498),
            .in2(N__44182),
            .in3(N__44170),
            .lcout(n21916),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i227_2_lut_LC_17_7_3.C_ON=1'b0;
    defparam i227_2_lut_LC_17_7_3.SEQ_MODE=4'b0000;
    defparam i227_2_lut_LC_17_7_3.LUT_INIT=16'b0000000011001100;
    LogicCell40 i227_2_lut_LC_17_7_3 (
            .in0(_gnd_net_),
            .in1(N__49800),
            .in2(_gnd_net_),
            .in3(N__49641),
            .lcout(n1252),
            .ltout(n1252_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_342_Mux_1_i2_3_lut_4_lut_LC_17_7_4.C_ON=1'b0;
    defparam comm_state_3__I_0_342_Mux_1_i2_3_lut_4_lut_LC_17_7_4.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_342_Mux_1_i2_3_lut_4_lut_LC_17_7_4.LUT_INIT=16'b0000110010101010;
    LogicCell40 comm_state_3__I_0_342_Mux_1_i2_3_lut_4_lut_LC_17_7_4 (
            .in0(N__49798),
            .in1(N__53680),
            .in2(N__44173),
            .in3(N__53495),
            .lcout(n2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19013_4_lut_LC_17_7_5.C_ON=1'b0;
    defparam i19013_4_lut_LC_17_7_5.SEQ_MODE=4'b0000;
    defparam i19013_4_lut_LC_17_7_5.LUT_INIT=16'b0100010101000000;
    LogicCell40 i19013_4_lut_LC_17_7_5 (
            .in0(N__53679),
            .in1(N__49113),
            .in2(N__51199),
            .in3(N__49799),
            .lcout(),
            .ltout(n21088_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19124_4_lut_LC_17_7_6.C_ON=1'b0;
    defparam i19124_4_lut_LC_17_7_6.SEQ_MODE=4'b0000;
    defparam i19124_4_lut_LC_17_7_6.LUT_INIT=16'b1100111111011101;
    LogicCell40 i19124_4_lut_LC_17_7_6 (
            .in0(N__46303),
            .in1(N__54245),
            .in2(N__44164),
            .in3(N__53496),
            .lcout(n14_adj_1497),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_342_Mux_1_i8_3_lut_4_lut_LC_17_7_7.C_ON=1'b0;
    defparam comm_state_3__I_0_342_Mux_1_i8_3_lut_4_lut_LC_17_7_7.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_342_Mux_1_i8_3_lut_4_lut_LC_17_7_7.LUT_INIT=16'b0001000110110001;
    LogicCell40 comm_state_3__I_0_342_Mux_1_i8_3_lut_4_lut_LC_17_7_7 (
            .in0(N__53497),
            .in1(N__44440),
            .in2(N__53830),
            .in3(N__44434),
            .lcout(n8_adj_1555),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i458_2_lut_LC_17_8_0.C_ON=1'b0;
    defparam i458_2_lut_LC_17_8_0.SEQ_MODE=4'b0000;
    defparam i458_2_lut_LC_17_8_0.LUT_INIT=16'b0101010100000000;
    LogicCell40 i458_2_lut_LC_17_8_0 (
            .in0(N__49755),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__49632),
            .lcout(n2342),
            .ltout(n2342_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i32_4_lut_LC_17_8_1.C_ON=1'b0;
    defparam i32_4_lut_LC_17_8_1.SEQ_MODE=4'b0000;
    defparam i32_4_lut_LC_17_8_1.LUT_INIT=16'b1110001011000000;
    LogicCell40 i32_4_lut_LC_17_8_1 (
            .in0(N__51198),
            .in1(N__53658),
            .in2(N__44422),
            .in3(N__44419),
            .lcout(),
            .ltout(n15_adj_1602_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_i2_LC_17_8_2.C_ON=1'b0;
    defparam comm_state_i2_LC_17_8_2.SEQ_MODE=4'b1000;
    defparam comm_state_i2_LC_17_8_2.LUT_INIT=16'b1000100011111000;
    LogicCell40 comm_state_i2_LC_17_8_2 (
            .in0(N__44371),
            .in1(N__44362),
            .in2(N__44374),
            .in3(N__53512),
            .lcout(comm_state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55109),
            .ce(N__49555),
            .sr(N__54609));
    defparam i1_2_lut_adj_277_LC_17_8_3.C_ON=1'b0;
    defparam i1_2_lut_adj_277_LC_17_8_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_277_LC_17_8_3.LUT_INIT=16'b0011001100000000;
    LogicCell40 i1_2_lut_adj_277_LC_17_8_3 (
            .in0(_gnd_net_),
            .in1(N__49751),
            .in2(_gnd_net_),
            .in3(N__51105),
            .lcout(n20571),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_4_lut_adj_254_LC_17_8_4.C_ON=1'b0;
    defparam i1_2_lut_4_lut_adj_254_LC_17_8_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_4_lut_adj_254_LC_17_8_4.LUT_INIT=16'b1111111101111101;
    LogicCell40 i1_2_lut_4_lut_adj_254_LC_17_8_4 (
            .in0(N__53656),
            .in1(N__49492),
            .in2(N__49348),
            .in3(N__49324),
            .lcout(n20641),
            .ltout(n20641_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i33_3_lut_LC_17_8_5.C_ON=1'b0;
    defparam i33_3_lut_LC_17_8_5.SEQ_MODE=4'b0000;
    defparam i33_3_lut_LC_17_8_5.LUT_INIT=16'b1110010011100100;
    LogicCell40 i33_3_lut_LC_17_8_5 (
            .in0(N__53511),
            .in1(N__53657),
            .in2(N__44365),
            .in3(_gnd_net_),
            .lcout(n12_adj_1603),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i22_4_lut_4_lut_LC_17_8_6.C_ON=1'b0;
    defparam i22_4_lut_4_lut_LC_17_8_6.SEQ_MODE=4'b0000;
    defparam i22_4_lut_4_lut_LC_17_8_6.LUT_INIT=16'b0100011001000100;
    LogicCell40 i22_4_lut_4_lut_LC_17_8_6 (
            .in0(N__53655),
            .in1(N__53510),
            .in2(N__49782),
            .in3(N__49633),
            .lcout(n7_adj_1588),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_312_LC_17_8_7.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_312_LC_17_8_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_312_LC_17_8_7.LUT_INIT=16'b1110111011111111;
    LogicCell40 i1_2_lut_3_lut_adj_312_LC_17_8_7 (
            .in0(N__54238),
            .in1(N__53654),
            .in2(_gnd_net_),
            .in3(N__51104),
            .lcout(n20650),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam secclk_cnt_3765_3766__i1_LC_17_9_0.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i1_LC_17_9_0.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i1_LC_17_9_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i1_LC_17_9_0 (
            .in0(_gnd_net_),
            .in1(N__44587),
            .in2(_gnd_net_),
            .in3(N__44575),
            .lcout(secclk_cnt_0),
            .ltout(),
            .carryin(bfn_17_9_0_),
            .carryout(n19447),
            .clk(N__56025),
            .ce(),
            .sr(N__44910));
    defparam secclk_cnt_3765_3766__i2_LC_17_9_1.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i2_LC_17_9_1.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i2_LC_17_9_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i2_LC_17_9_1 (
            .in0(_gnd_net_),
            .in1(N__44571),
            .in2(_gnd_net_),
            .in3(N__44557),
            .lcout(secclk_cnt_1),
            .ltout(),
            .carryin(n19447),
            .carryout(n19448),
            .clk(N__56025),
            .ce(),
            .sr(N__44910));
    defparam secclk_cnt_3765_3766__i3_LC_17_9_2.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i3_LC_17_9_2.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i3_LC_17_9_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i3_LC_17_9_2 (
            .in0(_gnd_net_),
            .in1(N__44554),
            .in2(_gnd_net_),
            .in3(N__44542),
            .lcout(secclk_cnt_2),
            .ltout(),
            .carryin(n19448),
            .carryout(n19449),
            .clk(N__56025),
            .ce(),
            .sr(N__44910));
    defparam secclk_cnt_3765_3766__i4_LC_17_9_3.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i4_LC_17_9_3.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i4_LC_17_9_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i4_LC_17_9_3 (
            .in0(_gnd_net_),
            .in1(N__44535),
            .in2(_gnd_net_),
            .in3(N__44524),
            .lcout(secclk_cnt_3),
            .ltout(),
            .carryin(n19449),
            .carryout(n19450),
            .clk(N__56025),
            .ce(),
            .sr(N__44910));
    defparam secclk_cnt_3765_3766__i5_LC_17_9_4.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i5_LC_17_9_4.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i5_LC_17_9_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i5_LC_17_9_4 (
            .in0(_gnd_net_),
            .in1(N__44521),
            .in2(_gnd_net_),
            .in3(N__44509),
            .lcout(secclk_cnt_4),
            .ltout(),
            .carryin(n19450),
            .carryout(n19451),
            .clk(N__56025),
            .ce(),
            .sr(N__44910));
    defparam secclk_cnt_3765_3766__i6_LC_17_9_5.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i6_LC_17_9_5.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i6_LC_17_9_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i6_LC_17_9_5 (
            .in0(_gnd_net_),
            .in1(N__44505),
            .in2(_gnd_net_),
            .in3(N__44491),
            .lcout(secclk_cnt_5),
            .ltout(),
            .carryin(n19451),
            .carryout(n19452),
            .clk(N__56025),
            .ce(),
            .sr(N__44910));
    defparam secclk_cnt_3765_3766__i7_LC_17_9_6.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i7_LC_17_9_6.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i7_LC_17_9_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i7_LC_17_9_6 (
            .in0(_gnd_net_),
            .in1(N__44488),
            .in2(_gnd_net_),
            .in3(N__44476),
            .lcout(secclk_cnt_6),
            .ltout(),
            .carryin(n19452),
            .carryout(n19453),
            .clk(N__56025),
            .ce(),
            .sr(N__44910));
    defparam secclk_cnt_3765_3766__i8_LC_17_9_7.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i8_LC_17_9_7.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i8_LC_17_9_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i8_LC_17_9_7 (
            .in0(_gnd_net_),
            .in1(N__44472),
            .in2(_gnd_net_),
            .in3(N__44458),
            .lcout(secclk_cnt_7),
            .ltout(),
            .carryin(n19453),
            .carryout(n19454),
            .clk(N__56025),
            .ce(),
            .sr(N__44910));
    defparam secclk_cnt_3765_3766__i9_LC_17_10_0.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i9_LC_17_10_0.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i9_LC_17_10_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i9_LC_17_10_0 (
            .in0(_gnd_net_),
            .in1(N__44455),
            .in2(_gnd_net_),
            .in3(N__44443),
            .lcout(secclk_cnt_8),
            .ltout(),
            .carryin(bfn_17_10_0_),
            .carryout(n19455),
            .clk(N__56027),
            .ce(),
            .sr(N__44906));
    defparam secclk_cnt_3765_3766__i10_LC_17_10_1.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i10_LC_17_10_1.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i10_LC_17_10_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i10_LC_17_10_1 (
            .in0(_gnd_net_),
            .in1(N__44704),
            .in2(_gnd_net_),
            .in3(N__44692),
            .lcout(secclk_cnt_9),
            .ltout(),
            .carryin(n19455),
            .carryout(n19456),
            .clk(N__56027),
            .ce(),
            .sr(N__44906));
    defparam secclk_cnt_3765_3766__i11_LC_17_10_2.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i11_LC_17_10_2.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i11_LC_17_10_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i11_LC_17_10_2 (
            .in0(_gnd_net_),
            .in1(N__44688),
            .in2(_gnd_net_),
            .in3(N__44674),
            .lcout(secclk_cnt_10),
            .ltout(),
            .carryin(n19456),
            .carryout(n19457),
            .clk(N__56027),
            .ce(),
            .sr(N__44906));
    defparam secclk_cnt_3765_3766__i12_LC_17_10_3.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i12_LC_17_10_3.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i12_LC_17_10_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i12_LC_17_10_3 (
            .in0(_gnd_net_),
            .in1(N__44670),
            .in2(_gnd_net_),
            .in3(N__44656),
            .lcout(secclk_cnt_11),
            .ltout(),
            .carryin(n19457),
            .carryout(n19458),
            .clk(N__56027),
            .ce(),
            .sr(N__44906));
    defparam secclk_cnt_3765_3766__i13_LC_17_10_4.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i13_LC_17_10_4.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i13_LC_17_10_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i13_LC_17_10_4 (
            .in0(_gnd_net_),
            .in1(N__53067),
            .in2(_gnd_net_),
            .in3(N__44653),
            .lcout(secclk_cnt_12),
            .ltout(),
            .carryin(n19458),
            .carryout(n19459),
            .clk(N__56027),
            .ce(),
            .sr(N__44906));
    defparam secclk_cnt_3765_3766__i14_LC_17_10_5.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i14_LC_17_10_5.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i14_LC_17_10_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i14_LC_17_10_5 (
            .in0(_gnd_net_),
            .in1(N__44649),
            .in2(_gnd_net_),
            .in3(N__44635),
            .lcout(secclk_cnt_13),
            .ltout(),
            .carryin(n19459),
            .carryout(n19460),
            .clk(N__56027),
            .ce(),
            .sr(N__44906));
    defparam secclk_cnt_3765_3766__i15_LC_17_10_6.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i15_LC_17_10_6.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i15_LC_17_10_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i15_LC_17_10_6 (
            .in0(_gnd_net_),
            .in1(N__44632),
            .in2(_gnd_net_),
            .in3(N__44620),
            .lcout(secclk_cnt_14),
            .ltout(),
            .carryin(n19460),
            .carryout(n19461),
            .clk(N__56027),
            .ce(),
            .sr(N__44906));
    defparam secclk_cnt_3765_3766__i16_LC_17_10_7.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i16_LC_17_10_7.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i16_LC_17_10_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i16_LC_17_10_7 (
            .in0(_gnd_net_),
            .in1(N__44617),
            .in2(_gnd_net_),
            .in3(N__44605),
            .lcout(secclk_cnt_15),
            .ltout(),
            .carryin(n19461),
            .carryout(n19462),
            .clk(N__56027),
            .ce(),
            .sr(N__44906));
    defparam secclk_cnt_3765_3766__i17_LC_17_11_0.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i17_LC_17_11_0.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i17_LC_17_11_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i17_LC_17_11_0 (
            .in0(_gnd_net_),
            .in1(N__44602),
            .in2(_gnd_net_),
            .in3(N__44590),
            .lcout(secclk_cnt_16),
            .ltout(),
            .carryin(bfn_17_11_0_),
            .carryout(n19463),
            .clk(N__56028),
            .ce(),
            .sr(N__44911));
    defparam secclk_cnt_3765_3766__i18_LC_17_11_1.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i18_LC_17_11_1.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i18_LC_17_11_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i18_LC_17_11_1 (
            .in0(_gnd_net_),
            .in1(N__44968),
            .in2(_gnd_net_),
            .in3(N__44956),
            .lcout(secclk_cnt_17),
            .ltout(),
            .carryin(n19463),
            .carryout(n19464),
            .clk(N__56028),
            .ce(),
            .sr(N__44911));
    defparam secclk_cnt_3765_3766__i19_LC_17_11_2.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i19_LC_17_11_2.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i19_LC_17_11_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i19_LC_17_11_2 (
            .in0(_gnd_net_),
            .in1(N__44952),
            .in2(_gnd_net_),
            .in3(N__44938),
            .lcout(secclk_cnt_18),
            .ltout(),
            .carryin(n19464),
            .carryout(n19465),
            .clk(N__56028),
            .ce(),
            .sr(N__44911));
    defparam secclk_cnt_3765_3766__i20_LC_17_11_3.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i20_LC_17_11_3.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i20_LC_17_11_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i20_LC_17_11_3 (
            .in0(_gnd_net_),
            .in1(N__53103),
            .in2(_gnd_net_),
            .in3(N__44935),
            .lcout(secclk_cnt_19),
            .ltout(),
            .carryin(n19465),
            .carryout(n19466),
            .clk(N__56028),
            .ce(),
            .sr(N__44911));
    defparam secclk_cnt_3765_3766__i21_LC_17_11_4.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i21_LC_17_11_4.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i21_LC_17_11_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i21_LC_17_11_4 (
            .in0(_gnd_net_),
            .in1(N__44932),
            .in2(_gnd_net_),
            .in3(N__44920),
            .lcout(secclk_cnt_20),
            .ltout(),
            .carryin(n19466),
            .carryout(n19467),
            .clk(N__56028),
            .ce(),
            .sr(N__44911));
    defparam secclk_cnt_3765_3766__i22_LC_17_11_5.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i22_LC_17_11_5.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i22_LC_17_11_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i22_LC_17_11_5 (
            .in0(_gnd_net_),
            .in1(N__53088),
            .in2(_gnd_net_),
            .in3(N__44917),
            .lcout(secclk_cnt_21),
            .ltout(),
            .carryin(n19467),
            .carryout(n19468),
            .clk(N__56028),
            .ce(),
            .sr(N__44911));
    defparam secclk_cnt_3765_3766__i23_LC_17_11_6.C_ON=1'b0;
    defparam secclk_cnt_3765_3766__i23_LC_17_11_6.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i23_LC_17_11_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i23_LC_17_11_6 (
            .in0(_gnd_net_),
            .in1(N__53052),
            .in2(_gnd_net_),
            .in3(N__44914),
            .lcout(secclk_cnt_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56028),
            .ce(),
            .sr(N__44911));
    defparam i1_2_lut_3_lut_adj_307_LC_17_12_0.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_307_LC_17_12_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_307_LC_17_12_0.LUT_INIT=16'b0000000000100010;
    LogicCell40 i1_2_lut_3_lut_adj_307_LC_17_12_0 (
            .in0(N__44872),
            .in1(N__51204),
            .in2(_gnd_net_),
            .in3(N__53828),
            .lcout(n14_adj_1556),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_4_i23_3_lut_LC_17_12_1.C_ON=1'b0;
    defparam mux_128_Mux_4_i23_3_lut_LC_17_12_1.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_4_i23_3_lut_LC_17_12_1.LUT_INIT=16'b1110111000100010;
    LogicCell40 mux_128_Mux_4_i23_3_lut_LC_17_12_1 (
            .in0(N__44754),
            .in1(N__56927),
            .in2(_gnd_net_),
            .in3(N__44725),
            .lcout(n23_adj_1517),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_4_i22_3_lut_LC_17_12_2.C_ON=1'b0;
    defparam mux_130_Mux_4_i22_3_lut_LC_17_12_2.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_4_i22_3_lut_LC_17_12_2.LUT_INIT=16'b1100110010101010;
    LogicCell40 mux_130_Mux_4_i22_3_lut_LC_17_12_2 (
            .in0(N__48828),
            .in1(N__51310),
            .in2(_gnd_net_),
            .in3(N__47825),
            .lcout(n22_adj_1606),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12250_3_lut_LC_17_12_3.C_ON=1'b0;
    defparam i12250_3_lut_LC_17_12_3.SEQ_MODE=4'b0000;
    defparam i12250_3_lut_LC_17_12_3.LUT_INIT=16'b1101110100000000;
    LogicCell40 i12250_3_lut_LC_17_12_3 (
            .in0(N__51205),
            .in1(N__54451),
            .in2(_gnd_net_),
            .in3(N__45431),
            .lcout(n14652),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18804_2_lut_LC_17_12_4.C_ON=1'b0;
    defparam i18804_2_lut_LC_17_12_4.SEQ_MODE=4'b0000;
    defparam i18804_2_lut_LC_17_12_4.LUT_INIT=16'b0101010100000000;
    LogicCell40 i18804_2_lut_LC_17_12_4 (
            .in0(N__56928),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45086),
            .lcout(n21022),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_317_LC_17_12_5.C_ON=1'b0;
    defparam i1_4_lut_adj_317_LC_17_12_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_317_LC_17_12_5.LUT_INIT=16'b0111101111011110;
    LogicCell40 i1_4_lut_adj_317_LC_17_12_5 (
            .in0(N__45039),
            .in1(N__51578),
            .in2(N__50094),
            .in3(N__45445),
            .lcout(n4_adj_1576),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_length_i2_LC_17_12_6.C_ON=1'b0;
    defparam comm_length_i2_LC_17_12_6.SEQ_MODE=4'b1000;
    defparam comm_length_i2_LC_17_12_6.LUT_INIT=16'b0101000011001100;
    LogicCell40 comm_length_i2_LC_17_12_6 (
            .in0(N__56929),
            .in1(N__45040),
            .in2(N__45058),
            .in3(N__45432),
            .lcout(comm_length_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55156),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19355_LC_17_13_0.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19355_LC_17_13_0.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19355_LC_17_13_0.LUT_INIT=16'b1101101010001010;
    LogicCell40 comm_cmd_1__bdd_4_lut_19355_LC_17_13_0 (
            .in0(N__57535),
            .in1(N__44998),
            .in2(N__47849),
            .in3(N__44974),
            .lcout(),
            .ltout(n21955_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n21955_bdd_4_lut_LC_17_13_1.C_ON=1'b0;
    defparam n21955_bdd_4_lut_LC_17_13_1.SEQ_MODE=4'b0000;
    defparam n21955_bdd_4_lut_LC_17_13_1.LUT_INIT=16'b1111001011000010;
    LogicCell40 n21955_bdd_4_lut_LC_17_13_1 (
            .in0(N__45451),
            .in1(N__47829),
            .in2(N__45031),
            .in3(N__45022),
            .lcout(n21958),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18787_2_lut_LC_17_13_2.C_ON=1'b0;
    defparam i18787_2_lut_LC_17_13_2.SEQ_MODE=4'b0000;
    defparam i18787_2_lut_LC_17_13_2.LUT_INIT=16'b0100010001000100;
    LogicCell40 i18787_2_lut_LC_17_13_2 (
            .in0(N__56932),
            .in1(N__45254),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(n21024),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19055_2_lut_LC_17_13_3.C_ON=1'b0;
    defparam i19055_2_lut_LC_17_13_3.SEQ_MODE=4'b0000;
    defparam i19055_2_lut_LC_17_13_3.LUT_INIT=16'b0000000011001100;
    LogicCell40 i19055_2_lut_LC_17_13_3 (
            .in0(_gnd_net_),
            .in1(N__45016),
            .in2(_gnd_net_),
            .in3(N__56931),
            .lcout(n20950),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_3_i26_3_lut_LC_17_13_4.C_ON=1'b0;
    defparam mux_128_Mux_3_i26_3_lut_LC_17_13_4.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_3_i26_3_lut_LC_17_13_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_128_Mux_3_i26_3_lut_LC_17_13_4 (
            .in0(N__56930),
            .in1(N__44992),
            .in2(_gnd_net_),
            .in3(N__47240),
            .lcout(n26_adj_1519),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_3_i23_3_lut_LC_17_13_5.C_ON=1'b0;
    defparam mux_128_Mux_3_i23_3_lut_LC_17_13_5.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_3_i23_3_lut_LC_17_13_5.LUT_INIT=16'b1110111000100010;
    LogicCell40 mux_128_Mux_3_i23_3_lut_LC_17_13_5 (
            .in0(N__45510),
            .in1(N__56933),
            .in2(_gnd_net_),
            .in3(N__45478),
            .lcout(n23_adj_1518),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_length_i0_LC_17_13_6.C_ON=1'b0;
    defparam comm_length_i0_LC_17_13_6.SEQ_MODE=4'b1000;
    defparam comm_length_i0_LC_17_13_6.LUT_INIT=16'b0001001110100110;
    LogicCell40 comm_length_i0_LC_17_13_6 (
            .in0(N__57536),
            .in1(N__56311),
            .in2(N__56977),
            .in3(N__47831),
            .lcout(comm_length_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55171),
            .ce(N__45439),
            .sr(N__45403));
    defparam comm_length_i1_LC_17_13_7.C_ON=1'b0;
    defparam comm_length_i1_LC_17_13_7.SEQ_MODE=4'b1000;
    defparam comm_length_i1_LC_17_13_7.LUT_INIT=16'b1011110011101111;
    LogicCell40 comm_length_i1_LC_17_13_7 (
            .in0(N__47830),
            .in1(N__56934),
            .in2(N__56341),
            .in3(N__57537),
            .lcout(comm_length_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55171),
            .ce(N__45439),
            .sr(N__45403));
    defparam \ADC_IAC.ADC_DATA_i7_LC_17_14_0 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i7_LC_17_14_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i7_LC_17_14_0 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_IAC.ADC_DATA_i7_LC_17_14_0  (
            .in0(N__49008),
            .in1(N__50962),
            .in2(N__47880),
            .in3(N__45155),
            .lcout(buf_adcdata_iac_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55185),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_280_LC_17_14_2.C_ON=1'b0;
    defparam i1_4_lut_adj_280_LC_17_14_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_280_LC_17_14_2.LUT_INIT=16'b1000100010001010;
    LogicCell40 i1_4_lut_adj_280_LC_17_14_2 (
            .in0(N__54441),
            .in1(N__51782),
            .in2(N__45394),
            .in3(N__45376),
            .lcout(n12381),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7_4_lut_adj_58_LC_17_14_3.C_ON=1'b0;
    defparam i7_4_lut_adj_58_LC_17_14_3.SEQ_MODE=4'b0000;
    defparam i7_4_lut_adj_58_LC_17_14_3.LUT_INIT=16'b0111110110111110;
    LogicCell40 i7_4_lut_adj_58_LC_17_14_3 (
            .in0(N__48699),
            .in1(N__47241),
            .in2(N__45256),
            .in3(N__45227),
            .lcout(n23_adj_1491),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i7_LC_17_14_4 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i7_LC_17_14_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i7_LC_17_14_4 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i7_LC_17_14_4  (
            .in0(N__48535),
            .in1(N__48347),
            .in2(N__45201),
            .in3(N__47928),
            .lcout(buf_adcdata_vac_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55185),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i15_LC_17_14_5 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i15_LC_17_14_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i15_LC_17_14_5 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i15_LC_17_14_5  (
            .in0(N__50961),
            .in1(N__48798),
            .in2(N__45159),
            .in3(N__50519),
            .lcout(cmd_rdadctmp_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55185),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i16_LC_17_14_6 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i16_LC_17_14_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i16_LC_17_14_6 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i16_LC_17_14_6  (
            .in0(N__50518),
            .in1(N__45113),
            .in2(N__45163),
            .in3(N__50963),
            .lcout(cmd_rdadctmp_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55185),
            .ce(),
            .sr(_gnd_net_));
    defparam i46_2_lut_LC_17_14_7.C_ON=1'b0;
    defparam i46_2_lut_LC_17_14_7.SEQ_MODE=4'b0000;
    defparam i46_2_lut_LC_17_14_7.LUT_INIT=16'b0011001111001100;
    LogicCell40 i46_2_lut_LC_17_14_7 (
            .in0(_gnd_net_),
            .in1(N__49767),
            .in2(_gnd_net_),
            .in3(N__53987),
            .lcout(n23_adj_1574),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i5_LC_17_15_0.C_ON=1'b0;
    defparam data_index_i5_LC_17_15_0.SEQ_MODE=4'b1000;
    defparam data_index_i5_LC_17_15_0.LUT_INIT=16'b0010111100100000;
    LogicCell40 data_index_i5_LC_17_15_0 (
            .in0(N__46060),
            .in1(N__51786),
            .in2(N__54599),
            .in3(N__46054),
            .lcout(data_index_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55200),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_LC_17_15_2.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_LC_17_15_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_LC_17_15_2.LUT_INIT=16'b0001000011111111;
    LogicCell40 i1_2_lut_3_lut_4_lut_LC_17_15_2 (
            .in0(N__51206),
            .in1(N__53829),
            .in2(N__54598),
            .in3(N__45810),
            .lcout(n16708),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15037_2_lut_LC_17_15_4.C_ON=1'b0;
    defparam i15037_2_lut_LC_17_15_4.SEQ_MODE=4'b0000;
    defparam i15037_2_lut_LC_17_15_4.LUT_INIT=16'b1010101011111111;
    LogicCell40 i15037_2_lut_LC_17_15_4 (
            .in0(N__53986),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53466),
            .lcout(n3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_4_lut_adj_243_LC_17_15_7.C_ON=1'b0;
    defparam i1_2_lut_4_lut_adj_243_LC_17_15_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_4_lut_adj_243_LC_17_15_7.LUT_INIT=16'b1110111111111111;
    LogicCell40 i1_2_lut_4_lut_adj_243_LC_17_15_7 (
            .in0(N__49801),
            .in1(N__54433),
            .in2(N__51259),
            .in3(N__49645),
            .lcout(n4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_251_LC_17_16_4.C_ON=1'b0;
    defparam i1_4_lut_adj_251_LC_17_16_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_251_LC_17_16_4.LUT_INIT=16'b1000101011001111;
    LogicCell40 i1_4_lut_adj_251_LC_17_16_4 (
            .in0(N__49240),
            .in1(N__54440),
            .in2(N__50980),
            .in3(N__45933),
            .lcout(n11805),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i15_LC_17_17_1.C_ON=1'b0;
    defparam buf_dds0_i15_LC_17_17_1.SEQ_MODE=4'b1000;
    defparam buf_dds0_i15_LC_17_17_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 buf_dds0_i15_LC_17_17_1 (
            .in0(N__45767),
            .in1(N__45581),
            .in2(_gnd_net_),
            .in3(N__45674),
            .lcout(buf_dds0_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55223),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_188_i9_2_lut_3_lut_LC_17_17_4.C_ON=1'b0;
    defparam equal_188_i9_2_lut_3_lut_LC_17_17_4.SEQ_MODE=4'b0000;
    defparam equal_188_i9_2_lut_3_lut_LC_17_17_4.LUT_INIT=16'b1111111111011101;
    LogicCell40 equal_188_i9_2_lut_3_lut_LC_17_17_4 (
            .in0(N__57534),
            .in1(N__56989),
            .in2(_gnd_net_),
            .in3(N__47850),
            .lcout(n9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.dds_state_i1_LC_17_18_0 .C_ON=1'b0;
    defparam \SIG_DDS.dds_state_i1_LC_17_18_0 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.dds_state_i1_LC_17_18_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \SIG_DDS.dds_state_i1_LC_17_18_0  (
            .in0(_gnd_net_),
            .in1(N__55862),
            .in2(_gnd_net_),
            .in3(N__55739),
            .lcout(dds_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55232),
            .ce(N__45534),
            .sr(N__55659));
    defparam \comm_spi.data_tx_i5_12217_12218_reset_LC_18_4_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i5_12217_12218_reset_LC_18_4_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i5_12217_12218_reset_LC_18_4_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i5_12217_12218_reset_LC_18_4_0  (
            .in0(N__46273),
            .in1(N__46231),
            .in2(_gnd_net_),
            .in3(N__46138),
            .lcout(\comm_spi.n14620 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52417),
            .ce(),
            .sr(N__46282));
    defparam \comm_spi.data_tx_i5_12217_12218_set_LC_18_5_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i5_12217_12218_set_LC_18_5_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i5_12217_12218_set_LC_18_5_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i5_12217_12218_set_LC_18_5_0  (
            .in0(N__46269),
            .in1(N__46227),
            .in2(_gnd_net_),
            .in3(N__46137),
            .lcout(\comm_spi.n14619 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52426),
            .ce(),
            .sr(N__48709));
    defparam \comm_spi.data_tx_i4_12213_12214_set_LC_18_6_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i4_12213_12214_set_LC_18_6_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i4_12213_12214_set_LC_18_6_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i4_12213_12214_set_LC_18_6_0  (
            .in0(N__46207),
            .in1(N__46180),
            .in2(_gnd_net_),
            .in3(N__46159),
            .lcout(\comm_spi.n14615 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52360),
            .ce(),
            .sr(N__46216));
    defparam \comm_spi.data_tx_i4_12213_12214_reset_LC_18_7_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i4_12213_12214_reset_LC_18_7_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i4_12213_12214_reset_LC_18_7_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i4_12213_12214_reset_LC_18_7_0  (
            .in0(N__46206),
            .in1(N__46179),
            .in2(_gnd_net_),
            .in3(N__46155),
            .lcout(\comm_spi.n14616 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52430),
            .ce(),
            .sr(N__53131));
    defparam comm_state_3__I_0_342_Mux_3_i7_4_lut_LC_18_8_0.C_ON=1'b0;
    defparam comm_state_3__I_0_342_Mux_3_i7_4_lut_LC_18_8_0.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_342_Mux_3_i7_4_lut_LC_18_8_0.LUT_INIT=16'b1110111011110000;
    LogicCell40 comm_state_3__I_0_342_Mux_3_i7_4_lut_LC_18_8_0 (
            .in0(N__46120),
            .in1(N__52233),
            .in2(N__46111),
            .in3(N__51062),
            .lcout(),
            .ltout(n17658_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_i3_LC_18_8_1.C_ON=1'b0;
    defparam comm_state_i3_LC_18_8_1.SEQ_MODE=4'b1000;
    defparam comm_state_i3_LC_18_8_1.LUT_INIT=16'b0100010000001111;
    LogicCell40 comm_state_i3_LC_18_8_1 (
            .in0(N__51919),
            .in1(N__46096),
            .in2(N__46087),
            .in3(N__54176),
            .lcout(comm_state_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55121),
            .ce(N__46453),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_260_LC_18_8_4.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_260_LC_18_8_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_260_LC_18_8_4.LUT_INIT=16'b1111111111011101;
    LogicCell40 i1_2_lut_3_lut_adj_260_LC_18_8_4 (
            .in0(N__54175),
            .in1(N__51061),
            .in2(_gnd_net_),
            .in3(N__53637),
            .lcout(n12220),
            .ltout(n12220_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_LC_18_8_5.C_ON=1'b0;
    defparam i1_4_lut_LC_18_8_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_LC_18_8_5.LUT_INIT=16'b1110111011100000;
    LogicCell40 i1_4_lut_LC_18_8_5 (
            .in0(N__46084),
            .in1(N__46438),
            .in2(N__46063),
            .in3(N__46398),
            .lcout(),
            .ltout(n4_adj_1483_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_adj_52_LC_18_8_6.C_ON=1'b0;
    defparam i2_4_lut_adj_52_LC_18_8_6.SEQ_MODE=4'b0000;
    defparam i2_4_lut_adj_52_LC_18_8_6.LUT_INIT=16'b1111000010110000;
    LogicCell40 i2_4_lut_adj_52_LC_18_8_6 (
            .in0(N__46467),
            .in1(N__49750),
            .in2(N__46510),
            .in3(N__46507),
            .lcout(n20510),
            .ltout(n20510_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_146_LC_18_8_7.C_ON=1'b0;
    defparam i1_4_lut_adj_146_LC_18_8_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_146_LC_18_8_7.LUT_INIT=16'b1010000010000000;
    LogicCell40 i1_4_lut_adj_146_LC_18_8_7 (
            .in0(N__46387),
            .in1(N__46483),
            .in2(N__46471),
            .in3(N__46468),
            .lcout(n20534),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_2_lut_3_lut_LC_18_9_0.C_ON=1'b0;
    defparam i3_2_lut_3_lut_LC_18_9_0.SEQ_MODE=4'b0000;
    defparam i3_2_lut_3_lut_LC_18_9_0.LUT_INIT=16'b1111111111111100;
    LogicCell40 i3_2_lut_3_lut_LC_18_9_0 (
            .in0(_gnd_net_),
            .in1(N__53474),
            .in2(N__49796),
            .in3(N__49626),
            .lcout(n11810),
            .ltout(n11810_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_LC_18_9_1.C_ON=1'b0;
    defparam i1_3_lut_LC_18_9_1.SEQ_MODE=4'b0000;
    defparam i1_3_lut_LC_18_9_1.LUT_INIT=16'b1111101010101010;
    LogicCell40 i1_3_lut_LC_18_9_1 (
            .in0(N__49140),
            .in1(_gnd_net_),
            .in2(N__46432),
            .in3(N__46399),
            .lcout(),
            .ltout(n20672_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_71_LC_18_9_2.C_ON=1'b0;
    defparam i1_4_lut_adj_71_LC_18_9_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_71_LC_18_9_2.LUT_INIT=16'b1110000000000000;
    LogicCell40 i1_4_lut_adj_71_LC_18_9_2 (
            .in0(N__46422),
            .in1(N__49126),
            .in2(N__46408),
            .in3(N__46405),
            .lcout(n20536),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_306_LC_18_9_4.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_306_LC_18_9_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_306_LC_18_9_4.LUT_INIT=16'b0011001111110011;
    LogicCell40 i1_2_lut_3_lut_adj_306_LC_18_9_4 (
            .in0(_gnd_net_),
            .in1(N__53475),
            .in2(N__49795),
            .in3(N__49625),
            .lcout(n20585),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_4_lut_adj_241_LC_18_9_5.C_ON=1'b0;
    defparam i1_4_lut_4_lut_adj_241_LC_18_9_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_4_lut_adj_241_LC_18_9_5.LUT_INIT=16'b1111010011111110;
    LogicCell40 i1_4_lut_4_lut_adj_241_LC_18_9_5 (
            .in0(N__49627),
            .in1(N__49774),
            .in2(N__49144),
            .in3(N__53438),
            .lcout(n11824),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_valid_85_LC_18_9_6 .C_ON=1'b0;
    defparam \comm_spi.data_valid_85_LC_18_9_6 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_valid_85_LC_18_9_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \comm_spi.data_valid_85_LC_18_9_6  (
            .in0(_gnd_net_),
            .in1(N__46381),
            .in2(_gnd_net_),
            .in3(N__46342),
            .lcout(comm_data_vld),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.data_valid_85C_net ),
            .ce(),
            .sr(N__55383));
    defparam i18843_2_lut_3_lut_LC_18_9_7.C_ON=1'b0;
    defparam i18843_2_lut_3_lut_LC_18_9_7.SEQ_MODE=4'b0000;
    defparam i18843_2_lut_3_lut_LC_18_9_7.LUT_INIT=16'b0001000100000000;
    LogicCell40 i18843_2_lut_3_lut_LC_18_9_7 (
            .in0(N__49628),
            .in1(N__49770),
            .in2(_gnd_net_),
            .in3(N__53900),
            .lcout(n21087),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_1__bdd_4_lut_19462_LC_18_10_0.C_ON=1'b0;
    defparam comm_index_1__bdd_4_lut_19462_LC_18_10_0.SEQ_MODE=4'b0000;
    defparam comm_index_1__bdd_4_lut_19462_LC_18_10_0.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_index_1__bdd_4_lut_19462_LC_18_10_0 (
            .in0(N__46753),
            .in1(N__49396),
            .in2(N__46717),
            .in3(N__50006),
            .lcout(),
            .ltout(n22063_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i4_LC_18_10_1.C_ON=1'b0;
    defparam comm_tx_buf_i4_LC_18_10_1.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i4_LC_18_10_1.LUT_INIT=16'b1111010010100100;
    LogicCell40 comm_tx_buf_i4_LC_18_10_1 (
            .in0(N__50007),
            .in1(N__46597),
            .in2(N__46741),
            .in3(N__46537),
            .lcout(comm_tx_buf_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55143),
            .ce(N__47104),
            .sr(N__47048));
    defparam i19042_2_lut_LC_18_10_2.C_ON=1'b0;
    defparam i19042_2_lut_LC_18_10_2.SEQ_MODE=4'b0000;
    defparam i19042_2_lut_LC_18_10_2.LUT_INIT=16'b0011001100000000;
    LogicCell40 i19042_2_lut_LC_18_10_2 (
            .in0(_gnd_net_),
            .in1(N__51516),
            .in2(_gnd_net_),
            .in3(N__46738),
            .lcout(n21081),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_137_Mux_4_i1_3_lut_LC_18_10_3.C_ON=1'b0;
    defparam mux_137_Mux_4_i1_3_lut_LC_18_10_3.SEQ_MODE=4'b0000;
    defparam mux_137_Mux_4_i1_3_lut_LC_18_10_3.LUT_INIT=16'b1110111001000100;
    LogicCell40 mux_137_Mux_4_i1_3_lut_LC_18_10_3 (
            .in0(N__51518),
            .in1(N__46707),
            .in2(_gnd_net_),
            .in3(N__46664),
            .lcout(n1_adj_1564),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_181_LC_18_10_5.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_181_LC_18_10_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_181_LC_18_10_5.LUT_INIT=16'b0001000100000000;
    LogicCell40 i1_2_lut_3_lut_adj_181_LC_18_10_5 (
            .in0(N__49781),
            .in1(N__49298),
            .in2(_gnd_net_),
            .in3(N__49624),
            .lcout(n18824),
            .ltout(n18824_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_LC_18_10_6.C_ON=1'b0;
    defparam i2_3_lut_LC_18_10_6.SEQ_MODE=4'b0000;
    defparam i2_3_lut_LC_18_10_6.LUT_INIT=16'b0011000000000000;
    LogicCell40 i2_3_lut_LC_18_10_6 (
            .in0(_gnd_net_),
            .in1(N__51515),
            .in2(N__46591),
            .in3(N__49395),
            .lcout(n20507),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_137_Mux_4_i2_3_lut_LC_18_10_7.C_ON=1'b0;
    defparam mux_137_Mux_4_i2_3_lut_LC_18_10_7.SEQ_MODE=4'b0000;
    defparam mux_137_Mux_4_i2_3_lut_LC_18_10_7.LUT_INIT=16'b1111101001010000;
    LogicCell40 mux_137_Mux_4_i2_3_lut_LC_18_10_7 (
            .in0(N__51517),
            .in1(_gnd_net_),
            .in2(N__46567),
            .in3(N__46552),
            .lcout(n2_adj_1565),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_137_Mux_1_i4_3_lut_LC_18_11_2.C_ON=1'b0;
    defparam mux_137_Mux_1_i4_3_lut_LC_18_11_2.SEQ_MODE=4'b0000;
    defparam mux_137_Mux_1_i4_3_lut_LC_18_11_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_137_Mux_1_i4_3_lut_LC_18_11_2 (
            .in0(N__46531),
            .in1(N__46522),
            .in2(_gnd_net_),
            .in3(N__51605),
            .lcout(),
            .ltout(n4_adj_1569_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18197_4_lut_LC_18_11_3.C_ON=1'b0;
    defparam i18197_4_lut_LC_18_11_3.SEQ_MODE=4'b0000;
    defparam i18197_4_lut_LC_18_11_3.LUT_INIT=16'b0111010000110000;
    LogicCell40 i18197_4_lut_LC_18_11_3 (
            .in0(N__51606),
            .in1(N__49467),
            .in2(N__47179),
            .in3(N__47176),
            .lcout(),
            .ltout(n20792_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i1_LC_18_11_4.C_ON=1'b0;
    defparam comm_tx_buf_i1_LC_18_11_4.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i1_LC_18_11_4.LUT_INIT=16'b1111010110100000;
    LogicCell40 comm_tx_buf_i1_LC_18_11_4 (
            .in0(N__50010),
            .in1(_gnd_net_),
            .in2(N__47158),
            .in3(N__47155),
            .lcout(comm_tx_buf_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55157),
            .ce(N__47135),
            .sr(N__47052));
    defparam i19037_3_lut_4_lut_LC_18_11_5.C_ON=1'b0;
    defparam i19037_3_lut_4_lut_LC_18_11_5.SEQ_MODE=4'b0000;
    defparam i19037_3_lut_4_lut_LC_18_11_5.LUT_INIT=16'b0000001000000000;
    LogicCell40 i19037_3_lut_4_lut_LC_18_11_5 (
            .in0(N__51604),
            .in1(N__50009),
            .in2(N__49514),
            .in3(N__49939),
            .lcout(n21069),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_cntvec_i0_i0_LC_18_12_0.C_ON=1'b1;
    defparam data_cntvec_i0_i0_LC_18_12_0.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i0_LC_18_12_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i0_LC_18_12_0 (
            .in0(_gnd_net_),
            .in1(N__46928),
            .in2(N__46987),
            .in3(_gnd_net_),
            .lcout(data_cntvec_0),
            .ltout(),
            .carryin(bfn_18_12_0_),
            .carryout(n19296),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__48662),
            .sr(N__48604));
    defparam data_cntvec_i0_i1_LC_18_12_1.C_ON=1'b1;
    defparam data_cntvec_i0_i1_LC_18_12_1.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i1_LC_18_12_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i1_LC_18_12_1 (
            .in0(_gnd_net_),
            .in1(N__46907),
            .in2(_gnd_net_),
            .in3(N__46885),
            .lcout(data_cntvec_1),
            .ltout(),
            .carryin(n19296),
            .carryout(n19297),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__48662),
            .sr(N__48604));
    defparam data_cntvec_i0_i2_LC_18_12_2.C_ON=1'b1;
    defparam data_cntvec_i0_i2_LC_18_12_2.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i2_LC_18_12_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i2_LC_18_12_2 (
            .in0(_gnd_net_),
            .in1(N__46871),
            .in2(_gnd_net_),
            .in3(N__46855),
            .lcout(data_cntvec_2),
            .ltout(),
            .carryin(n19297),
            .carryout(n19298),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__48662),
            .sr(N__48604));
    defparam data_cntvec_i0_i3_LC_18_12_3.C_ON=1'b1;
    defparam data_cntvec_i0_i3_LC_18_12_3.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i3_LC_18_12_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i3_LC_18_12_3 (
            .in0(_gnd_net_),
            .in1(N__46838),
            .in2(_gnd_net_),
            .in3(N__46816),
            .lcout(data_cntvec_3),
            .ltout(),
            .carryin(n19298),
            .carryout(n19299),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__48662),
            .sr(N__48604));
    defparam data_cntvec_i0_i4_LC_18_12_4.C_ON=1'b1;
    defparam data_cntvec_i0_i4_LC_18_12_4.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i4_LC_18_12_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i4_LC_18_12_4 (
            .in0(_gnd_net_),
            .in1(N__46802),
            .in2(_gnd_net_),
            .in3(N__46786),
            .lcout(data_cntvec_4),
            .ltout(),
            .carryin(n19299),
            .carryout(n19300),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__48662),
            .sr(N__48604));
    defparam data_cntvec_i0_i5_LC_18_12_5.C_ON=1'b1;
    defparam data_cntvec_i0_i5_LC_18_12_5.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i5_LC_18_12_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i5_LC_18_12_5 (
            .in0(_gnd_net_),
            .in1(N__46772),
            .in2(_gnd_net_),
            .in3(N__46756),
            .lcout(data_cntvec_5),
            .ltout(),
            .carryin(n19300),
            .carryout(n19301),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__48662),
            .sr(N__48604));
    defparam data_cntvec_i0_i6_LC_18_12_6.C_ON=1'b1;
    defparam data_cntvec_i0_i6_LC_18_12_6.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i6_LC_18_12_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i6_LC_18_12_6 (
            .in0(_gnd_net_),
            .in1(N__47402),
            .in2(_gnd_net_),
            .in3(N__47380),
            .lcout(data_cntvec_6),
            .ltout(),
            .carryin(n19301),
            .carryout(n19302),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__48662),
            .sr(N__48604));
    defparam data_cntvec_i0_i7_LC_18_12_7.C_ON=1'b1;
    defparam data_cntvec_i0_i7_LC_18_12_7.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i7_LC_18_12_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i7_LC_18_12_7 (
            .in0(_gnd_net_),
            .in1(N__47369),
            .in2(_gnd_net_),
            .in3(N__47347),
            .lcout(data_cntvec_7),
            .ltout(),
            .carryin(n19302),
            .carryout(n19303),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__48662),
            .sr(N__48604));
    defparam data_cntvec_i0_i8_LC_18_13_0.C_ON=1'b1;
    defparam data_cntvec_i0_i8_LC_18_13_0.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i8_LC_18_13_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i8_LC_18_13_0 (
            .in0(_gnd_net_),
            .in1(N__47336),
            .in2(_gnd_net_),
            .in3(N__47314),
            .lcout(data_cntvec_8),
            .ltout(),
            .carryin(bfn_18_13_0_),
            .carryout(n19304),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__48667),
            .sr(N__48603));
    defparam data_cntvec_i0_i9_LC_18_13_1.C_ON=1'b1;
    defparam data_cntvec_i0_i9_LC_18_13_1.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i9_LC_18_13_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i9_LC_18_13_1 (
            .in0(_gnd_net_),
            .in1(N__47297),
            .in2(_gnd_net_),
            .in3(N__47281),
            .lcout(data_cntvec_9),
            .ltout(),
            .carryin(n19304),
            .carryout(n19305),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__48667),
            .sr(N__48603));
    defparam data_cntvec_i0_i10_LC_18_13_2.C_ON=1'b1;
    defparam data_cntvec_i0_i10_LC_18_13_2.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i10_LC_18_13_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i10_LC_18_13_2 (
            .in0(_gnd_net_),
            .in1(N__47267),
            .in2(_gnd_net_),
            .in3(N__47245),
            .lcout(data_cntvec_10),
            .ltout(),
            .carryin(n19305),
            .carryout(n19306),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__48667),
            .sr(N__48603));
    defparam data_cntvec_i0_i11_LC_18_13_3.C_ON=1'b1;
    defparam data_cntvec_i0_i11_LC_18_13_3.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i11_LC_18_13_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i11_LC_18_13_3 (
            .in0(_gnd_net_),
            .in1(N__47242),
            .in2(_gnd_net_),
            .in3(N__47224),
            .lcout(data_cntvec_11),
            .ltout(),
            .carryin(n19306),
            .carryout(n19307),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__48667),
            .sr(N__48603));
    defparam data_cntvec_i0_i12_LC_18_13_4.C_ON=1'b1;
    defparam data_cntvec_i0_i12_LC_18_13_4.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i12_LC_18_13_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i12_LC_18_13_4 (
            .in0(_gnd_net_),
            .in1(N__47217),
            .in2(_gnd_net_),
            .in3(N__47203),
            .lcout(data_cntvec_12),
            .ltout(),
            .carryin(n19307),
            .carryout(n19308),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__48667),
            .sr(N__48603));
    defparam data_cntvec_i0_i13_LC_18_13_5.C_ON=1'b1;
    defparam data_cntvec_i0_i13_LC_18_13_5.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i13_LC_18_13_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i13_LC_18_13_5 (
            .in0(_gnd_net_),
            .in1(N__47196),
            .in2(_gnd_net_),
            .in3(N__47182),
            .lcout(data_cntvec_13),
            .ltout(),
            .carryin(n19308),
            .carryout(n19309),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__48667),
            .sr(N__48603));
    defparam data_cntvec_i0_i14_LC_18_13_6.C_ON=1'b1;
    defparam data_cntvec_i0_i14_LC_18_13_6.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i14_LC_18_13_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i14_LC_18_13_6 (
            .in0(_gnd_net_),
            .in1(N__48700),
            .in2(_gnd_net_),
            .in3(N__48688),
            .lcout(data_cntvec_14),
            .ltout(),
            .carryin(n19309),
            .carryout(n19310),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__48667),
            .sr(N__48603));
    defparam data_cntvec_i0_i15_LC_18_13_7.C_ON=1'b0;
    defparam data_cntvec_i0_i15_LC_18_13_7.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i15_LC_18_13_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i15_LC_18_13_7 (
            .in0(_gnd_net_),
            .in1(N__48681),
            .in2(_gnd_net_),
            .in3(N__48685),
            .lcout(data_cntvec_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__48667),
            .sr(N__48603));
    defparam i6956_2_lut_LC_18_14_0.C_ON=1'b0;
    defparam i6956_2_lut_LC_18_14_0.SEQ_MODE=4'b0000;
    defparam i6956_2_lut_LC_18_14_0.LUT_INIT=16'b1111111111001100;
    LogicCell40 i6956_2_lut_LC_18_14_0 (
            .in0(_gnd_net_),
            .in1(N__51221),
            .in2(_gnd_net_),
            .in3(N__53985),
            .lcout(n9273),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i6_LC_18_14_3 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i6_LC_18_14_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i6_LC_18_14_3 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i6_LC_18_14_3  (
            .in0(N__49009),
            .in1(N__50964),
            .in2(N__48799),
            .in3(N__48557),
            .lcout(buf_adcdata_iac_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55201),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i4_LC_18_14_4 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i4_LC_18_14_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i4_LC_18_14_4 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i4_LC_18_14_4  (
            .in0(N__48534),
            .in1(N__48348),
            .in2(N__47968),
            .in3(N__51330),
            .lcout(buf_adcdata_vac_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55201),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_7_i19_3_lut_LC_18_14_5.C_ON=1'b0;
    defparam mux_130_Mux_7_i19_3_lut_LC_18_14_5.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_7_i19_3_lut_LC_18_14_5.LUT_INIT=16'b1100110010101010;
    LogicCell40 mux_130_Mux_7_i19_3_lut_LC_18_14_5 (
            .in0(N__47924),
            .in1(N__47908),
            .in2(_gnd_net_),
            .in3(N__56988),
            .lcout(),
            .ltout(n19_adj_1589_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_7_i22_3_lut_LC_18_14_6.C_ON=1'b0;
    defparam mux_130_Mux_7_i22_3_lut_LC_18_14_6.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_7_i22_3_lut_LC_18_14_6.LUT_INIT=16'b1111000011001100;
    LogicCell40 mux_130_Mux_7_i22_3_lut_LC_18_14_6 (
            .in0(_gnd_net_),
            .in1(N__47873),
            .in2(N__47854),
            .in3(N__47846),
            .lcout(),
            .ltout(n22_adj_1590_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_7_i30_3_lut_LC_18_14_7.C_ON=1'b0;
    defparam mux_130_Mux_7_i30_3_lut_LC_18_14_7.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_7_i30_3_lut_LC_18_14_7.LUT_INIT=16'b1100110011110000;
    LogicCell40 mux_130_Mux_7_i30_3_lut_LC_18_14_7 (
            .in0(_gnd_net_),
            .in1(N__47443),
            .in2(N__47431),
            .in3(N__56316),
            .lcout(n30_adj_1591),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i5_LC_18_15_6 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i5_LC_18_15_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i5_LC_18_15_6 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i5_LC_18_15_6  (
            .in0(N__49000),
            .in1(N__50911),
            .in2(N__50323),
            .in3(N__49070),
            .lcout(buf_adcdata_iac_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55213),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i12_LC_18_16_0 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i12_LC_18_16_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i12_LC_18_16_0 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i12_LC_18_16_0  (
            .in0(N__50912),
            .in1(N__50540),
            .in2(N__49048),
            .in3(N__50527),
            .lcout(cmd_rdadctmp_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55224),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i4_LC_18_16_1 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i4_LC_18_16_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i4_LC_18_16_1 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i4_LC_18_16_1  (
            .in0(N__49004),
            .in1(N__50913),
            .in2(N__50547),
            .in3(N__48821),
            .lcout(buf_adcdata_iac_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55224),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.dds_state_i2_LC_18_16_3 .C_ON=1'b0;
    defparam \SIG_DDS.dds_state_i2_LC_18_16_3 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.dds_state_i2_LC_18_16_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \SIG_DDS.dds_state_i2_LC_18_16_3  (
            .in0(N__55613),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55795),
            .lcout(dds_state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55224),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i14_LC_18_17_2 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i14_LC_18_17_2 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i14_LC_18_17_2 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i14_LC_18_17_2  (
            .in0(N__48785),
            .in1(N__50914),
            .in2(N__50322),
            .in3(N__50526),
            .lcout(cmd_rdadctmp_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55233),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.iclk_40_12179_12180_set_LC_19_4_0 .C_ON=1'b0;
    defparam \comm_spi.iclk_40_12179_12180_set_LC_19_4_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.iclk_40_12179_12180_set_LC_19_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \comm_spi.iclk_40_12179_12180_set_LC_19_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52952),
            .lcout(\comm_spi.n14581 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55091),
            .ce(),
            .sr(N__48760));
    defparam \comm_spi.RESET_I_0_90_2_lut_LC_19_5_3 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_90_2_lut_LC_19_5_3 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_90_2_lut_LC_19_5_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \comm_spi.RESET_I_0_90_2_lut_LC_19_5_3  (
            .in0(N__52953),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55405),
            .lcout(\comm_spi.iclk_N_754 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_94_2_lut_LC_19_5_7 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_94_2_lut_LC_19_5_7 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_94_2_lut_LC_19_5_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \comm_spi.RESET_I_0_94_2_lut_LC_19_5_7  (
            .in0(_gnd_net_),
            .in1(N__48748),
            .in2(_gnd_net_),
            .in3(N__55406),
            .lcout(\comm_spi.data_tx_7__N_760 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i0_12175_12176_set_LC_19_6_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i0_12175_12176_set_LC_19_6_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i0_12175_12176_set_LC_19_6_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \comm_spi.data_tx_i0_12175_12176_set_LC_19_6_0  (
            .in0(N__52795),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\comm_spi.n14577 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52375),
            .ce(),
            .sr(N__52897));
    defparam comm_response_302_LC_19_7_0.C_ON=1'b0;
    defparam comm_response_302_LC_19_7_0.SEQ_MODE=4'b1000;
    defparam comm_response_302_LC_19_7_0.LUT_INIT=16'b0000010000100110;
    LogicCell40 comm_response_302_LC_19_7_0 (
            .in0(N__53742),
            .in1(N__54244),
            .in2(N__51264),
            .in3(N__53450),
            .lcout(ICE_GPMI_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55122),
            .ce(N__49249),
            .sr(_gnd_net_));
    defparam i1_3_lut_4_lut_adj_258_LC_19_7_1.C_ON=1'b0;
    defparam i1_3_lut_4_lut_adj_258_LC_19_7_1.SEQ_MODE=4'b0000;
    defparam i1_3_lut_4_lut_adj_258_LC_19_7_1.LUT_INIT=16'b1111001110100010;
    LogicCell40 i1_3_lut_4_lut_adj_258_LC_19_7_1 (
            .in0(N__53449),
            .in1(N__51234),
            .in2(N__54368),
            .in3(N__49186),
            .lcout(n11406),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i17_4_lut_3_lut_LC_19_7_2.C_ON=1'b0;
    defparam i17_4_lut_3_lut_LC_19_7_2.SEQ_MODE=4'b0000;
    defparam i17_4_lut_3_lut_LC_19_7_2.LUT_INIT=16'b0000010110100000;
    LogicCell40 i17_4_lut_3_lut_LC_19_7_2 (
            .in0(N__53741),
            .in1(_gnd_net_),
            .in2(N__51263),
            .in3(N__53448),
            .lcout(),
            .ltout(n10_adj_1572_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_285_LC_19_7_3.C_ON=1'b0;
    defparam i1_3_lut_adj_285_LC_19_7_3.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_285_LC_19_7_3.LUT_INIT=16'b1100100011001000;
    LogicCell40 i1_3_lut_adj_285_LC_19_7_3 (
            .in0(N__54240),
            .in1(N__49185),
            .in2(N__49147),
            .in3(_gnd_net_),
            .lcout(n11836),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_292_LC_19_7_7.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_292_LC_19_7_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_292_LC_19_7_7.LUT_INIT=16'b1110111011111111;
    LogicCell40 i1_2_lut_3_lut_adj_292_LC_19_7_7 (
            .in0(N__54239),
            .in1(N__51230),
            .in2(_gnd_net_),
            .in3(N__53740),
            .lcout(n20643),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_286_LC_19_8_2.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_286_LC_19_8_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_286_LC_19_8_2.LUT_INIT=16'b1011101111111111;
    LogicCell40 i1_2_lut_3_lut_adj_286_LC_19_8_2 (
            .in0(N__49699),
            .in1(N__53437),
            .in2(_gnd_net_),
            .in3(N__49635),
            .lcout(n4_adj_1596),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_i1_LC_19_9_0.C_ON=1'b0;
    defparam comm_index_i1_LC_19_9_0.SEQ_MODE=4'b1000;
    defparam comm_index_i1_LC_19_9_0.LUT_INIT=16'b1101111100100000;
    LogicCell40 comm_index_i1_LC_19_9_0 (
            .in0(N__49640),
            .in1(N__49769),
            .in2(N__51577),
            .in3(N__49462),
            .lcout(comm_index_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55144),
            .ce(N__49102),
            .sr(N__49093));
    defparam comm_index_i0_LC_19_9_1.C_ON=1'b0;
    defparam comm_index_i0_LC_19_9_1.SEQ_MODE=4'b1000;
    defparam comm_index_i0_LC_19_9_1.LUT_INIT=16'b1001100111001100;
    LogicCell40 comm_index_i0_LC_19_9_1 (
            .in0(N__49768),
            .in1(N__51533),
            .in2(_gnd_net_),
            .in3(N__49639),
            .lcout(comm_index_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55144),
            .ce(N__49102),
            .sr(N__49093));
    defparam comm_index_i2_LC_19_9_2.C_ON=1'b0;
    defparam comm_index_i2_LC_19_9_2.SEQ_MODE=4'b1000;
    defparam comm_index_i2_LC_19_9_2.LUT_INIT=16'b0110110011001100;
    LogicCell40 comm_index_i2_LC_19_9_2 (
            .in0(N__51537),
            .in1(N__50008),
            .in2(N__49513),
            .in3(N__49120),
            .lcout(comm_index_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55144),
            .ce(N__49102),
            .sr(N__49093));
    defparam \comm_spi.i19169_4_lut_3_lut_LC_19_10_0 .C_ON=1'b0;
    defparam \comm_spi.i19169_4_lut_3_lut_LC_19_10_0 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19169_4_lut_3_lut_LC_19_10_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.i19169_4_lut_3_lut_LC_19_10_0  (
            .in0(N__53193),
            .in1(N__50205),
            .in2(_gnd_net_),
            .in3(N__55382),
            .lcout(\comm_spi.n22647 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15191_2_lut_3_lut_LC_19_10_1.C_ON=1'b0;
    defparam i15191_2_lut_3_lut_LC_19_10_1.SEQ_MODE=4'b0000;
    defparam i15191_2_lut_3_lut_LC_19_10_1.LUT_INIT=16'b0000000001000100;
    LogicCell40 i15191_2_lut_3_lut_LC_19_10_1 (
            .in0(N__51225),
            .in1(N__50194),
            .in2(_gnd_net_),
            .in3(N__53884),
            .lcout(n14_adj_1557),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_297_LC_19_10_2.C_ON=1'b0;
    defparam i1_4_lut_adj_297_LC_19_10_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_297_LC_19_10_2.LUT_INIT=16'b0000001000000000;
    LogicCell40 i1_4_lut_adj_297_LC_19_10_2 (
            .in0(N__50002),
            .in1(N__53361),
            .in2(N__49429),
            .in3(N__49940),
            .lcout(n20563),
            .ltout(n20563_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19_4_lut_adj_295_LC_19_10_3.C_ON=1'b0;
    defparam i19_4_lut_adj_295_LC_19_10_3.SEQ_MODE=4'b0000;
    defparam i19_4_lut_adj_295_LC_19_10_3.LUT_INIT=16'b0100000001110011;
    LogicCell40 i19_4_lut_adj_295_LC_19_10_3 (
            .in0(N__51529),
            .in1(N__53883),
            .in2(N__49918),
            .in3(N__51684),
            .lcout(),
            .ltout(n12_adj_1539_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_296_LC_19_10_4.C_ON=1'b0;
    defparam i1_3_lut_adj_296_LC_19_10_4.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_296_LC_19_10_4.LUT_INIT=16'b1111110000000000;
    LogicCell40 i1_3_lut_adj_296_LC_19_10_4 (
            .in0(_gnd_net_),
            .in1(N__49915),
            .in2(N__49873),
            .in3(N__49846),
            .lcout(n12164),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_4_lut_LC_19_10_5.C_ON=1'b0;
    defparam i1_4_lut_4_lut_LC_19_10_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_4_lut_LC_19_10_5.LUT_INIT=16'b0100011000000000;
    LogicCell40 i1_4_lut_4_lut_LC_19_10_5 (
            .in0(N__51226),
            .in1(N__53885),
            .in2(N__49797),
            .in3(N__49634),
            .lcout(),
            .ltout(n21_adj_1573_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19127_4_lut_LC_19_10_6.C_ON=1'b0;
    defparam i19127_4_lut_LC_19_10_6.SEQ_MODE=4'b0000;
    defparam i19127_4_lut_LC_19_10_6.LUT_INIT=16'b0011111100110111;
    LogicCell40 i19127_4_lut_LC_19_10_6 (
            .in0(N__49573),
            .in1(N__56362),
            .in2(N__49558),
            .in3(N__51227),
            .lcout(n18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_adj_318_LC_19_11_0.C_ON=1'b0;
    defparam i2_3_lut_adj_318_LC_19_11_0.SEQ_MODE=4'b0000;
    defparam i2_3_lut_adj_318_LC_19_11_0.LUT_INIT=16'b1111111101100110;
    LogicCell40 i2_3_lut_adj_318_LC_19_11_0 (
            .in0(N__49463),
            .in1(N__49344),
            .in2(_gnd_net_),
            .in3(N__49323),
            .lcout(),
            .ltout(n5_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19063_3_lut_LC_19_11_1.C_ON=1'b0;
    defparam i19063_3_lut_LC_19_11_1.SEQ_MODE=4'b0000;
    defparam i19063_3_lut_LC_19_11_1.LUT_INIT=16'b1111101000000000;
    LogicCell40 i19063_3_lut_LC_19_11_1 (
            .in0(N__49303),
            .in1(_gnd_net_),
            .in2(N__49270),
            .in3(N__53882),
            .lcout(),
            .ltout(n21658_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18270_4_lut_LC_19_11_2.C_ON=1'b0;
    defparam i18270_4_lut_LC_19_11_2.SEQ_MODE=4'b0000;
    defparam i18270_4_lut_LC_19_11_2.LUT_INIT=16'b1111110010101010;
    LogicCell40 i18270_4_lut_LC_19_11_2 (
            .in0(N__52246),
            .in1(N__52234),
            .in2(N__52198),
            .in3(N__51229),
            .lcout(),
            .ltout(n20865_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_i0_LC_19_11_3.C_ON=1'b0;
    defparam comm_state_i0_LC_19_11_3.SEQ_MODE=4'b1000;
    defparam comm_state_i0_LC_19_11_3.LUT_INIT=16'b0011001111110000;
    LogicCell40 comm_state_i0_LC_19_11_3 (
            .in0(_gnd_net_),
            .in1(N__51881),
            .in2(N__51703),
            .in3(N__54536),
            .lcout(comm_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55173),
            .ce(N__51700),
            .sr(_gnd_net_));
    defparam i19_4_lut_adj_298_LC_19_11_6.C_ON=1'b0;
    defparam i19_4_lut_adj_298_LC_19_11_6.SEQ_MODE=4'b0000;
    defparam i19_4_lut_adj_298_LC_19_11_6.LUT_INIT=16'b1011000100010001;
    LogicCell40 i19_4_lut_adj_298_LC_19_11_6 (
            .in0(N__53881),
            .in1(N__51677),
            .in2(N__51619),
            .in3(N__51460),
            .lcout(n12_adj_1585),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15206_2_lut_3_lut_LC_19_12_5.C_ON=1'b0;
    defparam i15206_2_lut_3_lut_LC_19_12_5.SEQ_MODE=4'b0000;
    defparam i15206_2_lut_3_lut_LC_19_12_5.LUT_INIT=16'b0000000001000100;
    LogicCell40 i15206_2_lut_3_lut_LC_19_12_5 (
            .in0(N__51228),
            .in1(N__51442),
            .in2(_gnd_net_),
            .in3(N__53984),
            .lcout(n14_adj_1526),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_4_i19_3_lut_LC_19_13_3.C_ON=1'b0;
    defparam mux_130_Mux_4_i19_3_lut_LC_19_13_3.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_4_i19_3_lut_LC_19_13_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_130_Mux_4_i19_3_lut_LC_19_13_3 (
            .in0(N__51358),
            .in1(N__51326),
            .in2(_gnd_net_),
            .in3(N__56941),
            .lcout(n19_adj_1605),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18139_2_lut_3_lut_LC_19_14_1.C_ON=1'b0;
    defparam i18139_2_lut_3_lut_LC_19_14_1.SEQ_MODE=4'b0000;
    defparam i18139_2_lut_3_lut_LC_19_14_1.LUT_INIT=16'b1111111111101110;
    LogicCell40 i18139_2_lut_3_lut_LC_19_14_1 (
            .in0(N__51262),
            .in1(N__53983),
            .in2(_gnd_net_),
            .in3(N__53417),
            .lcout(n20734),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i13_LC_19_16_5 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i13_LC_19_16_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i13_LC_19_16_5 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i13_LC_19_16_5  (
            .in0(N__50315),
            .in1(N__50915),
            .in2(N__50548),
            .in3(N__50517),
            .lcout(cmd_rdadctmp_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55234),
            .ce(),
            .sr(_gnd_net_));
    defparam i14972_2_lut_2_lut_LC_19_17_2.C_ON=1'b0;
    defparam i14972_2_lut_2_lut_LC_19_17_2.SEQ_MODE=4'b0000;
    defparam i14972_2_lut_2_lut_LC_19_17_2.LUT_INIT=16'b0000000010101010;
    LogicCell40 i14972_2_lut_2_lut_LC_19_17_2 (
            .in0(N__50292),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50266),
            .lcout(CONT_SD),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.i23_4_lut_LC_19_18_7 .C_ON=1'b0;
    defparam \SIG_DDS.i23_4_lut_LC_19_18_7 .SEQ_MODE=4'b0000;
    defparam \SIG_DDS.i23_4_lut_LC_19_18_7 .LUT_INIT=16'b1010101010011101;
    LogicCell40 \SIG_DDS.i23_4_lut_LC_19_18_7  (
            .in0(N__55832),
            .in1(N__55738),
            .in2(N__53026),
            .in3(N__55585),
            .lcout(\SIG_DDS.n9_adj_1385 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.iclk_40_12179_12180_reset_LC_20_4_0 .C_ON=1'b0;
    defparam \comm_spi.iclk_40_12179_12180_reset_LC_20_4_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.iclk_40_12179_12180_reset_LC_20_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \comm_spi.iclk_40_12179_12180_reset_LC_20_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52941),
            .lcout(\comm_spi.n14582 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55102),
            .ce(),
            .sr(N__52906));
    defparam \comm_spi.RESET_I_0_91_2_lut_LC_20_5_0 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_91_2_lut_LC_20_5_0 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_91_2_lut_LC_20_5_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \comm_spi.RESET_I_0_91_2_lut_LC_20_5_0  (
            .in0(N__52942),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55407),
            .lcout(\comm_spi.iclk_N_755 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_2_lut_LC_20_6_2 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_2_lut_LC_20_6_2 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_2_lut_LC_20_6_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \comm_spi.RESET_I_0_2_lut_LC_20_6_2  (
            .in0(N__55377),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53258),
            .lcout(\comm_spi.data_tx_7__N_787 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_99_2_lut_LC_20_6_6 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_99_2_lut_LC_20_6_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_99_2_lut_LC_20_6_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \comm_spi.RESET_I_0_99_2_lut_LC_20_6_6  (
            .in0(N__55378),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53259),
            .lcout(\comm_spi.data_tx_7__N_765 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i0_12175_12176_reset_LC_20_7_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i0_12175_12176_reset_LC_20_7_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i0_12175_12176_reset_LC_20_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \comm_spi.data_tx_i0_12175_12176_reset_LC_20_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52724),
            .lcout(\comm_spi.n14578 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52437),
            .ce(),
            .sr(N__52534));
    defparam \comm_spi.data_tx_i1_12201_12202_reset_LC_20_8_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i1_12201_12202_reset_LC_20_8_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i1_12201_12202_reset_LC_20_8_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i1_12201_12202_reset_LC_20_8_0  (
            .in0(N__53233),
            .in1(N__52482),
            .in2(_gnd_net_),
            .in3(N__52497),
            .lcout(\comm_spi.n14604 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52415),
            .ce(),
            .sr(N__53176));
    defparam \comm_spi.data_tx_i1_12201_12202_set_LC_20_9_7 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i1_12201_12202_set_LC_20_9_7 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i1_12201_12202_set_LC_20_9_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \comm_spi.data_tx_i1_12201_12202_set_LC_20_9_7  (
            .in0(N__53229),
            .in1(N__52501),
            .in2(_gnd_net_),
            .in3(N__52486),
            .lcout(\comm_spi.n14603 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__52444),
            .ce(),
            .sr(N__53212));
    defparam \comm_spi.i19204_4_lut_3_lut_LC_20_10_0 .C_ON=1'b0;
    defparam \comm_spi.i19204_4_lut_3_lut_LC_20_10_0 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19204_4_lut_3_lut_LC_20_10_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.i19204_4_lut_3_lut_LC_20_10_0  (
            .in0(N__53260),
            .in1(N__53228),
            .in2(_gnd_net_),
            .in3(N__55404),
            .lcout(\comm_spi.n22650 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_98_2_lut_LC_20_10_2 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_98_2_lut_LC_20_10_2 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_98_2_lut_LC_20_10_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \comm_spi.RESET_I_0_98_2_lut_LC_20_10_2  (
            .in0(N__53200),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55403),
            .lcout(\comm_spi.data_tx_7__N_764 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_106_2_lut_LC_20_10_3 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_106_2_lut_LC_20_10_3 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_106_2_lut_LC_20_10_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \comm_spi.RESET_I_0_106_2_lut_LC_20_10_3  (
            .in0(N__55402),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53199),
            .lcout(\comm_spi.data_tx_7__N_784 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_103_2_lut_LC_20_10_6 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_103_2_lut_LC_20_10_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_103_2_lut_LC_20_10_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \comm_spi.RESET_I_0_103_2_lut_LC_20_10_6  (
            .in0(N__53148),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55401),
            .lcout(\comm_spi.data_tx_7__N_775 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6_4_lut_adj_231_LC_20_11_0.C_ON=1'b0;
    defparam i6_4_lut_adj_231_LC_20_11_0.SEQ_MODE=4'b0000;
    defparam i6_4_lut_adj_231_LC_20_11_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i6_4_lut_adj_231_LC_20_11_0 (
            .in0(N__57715),
            .in1(N__57568),
            .in2(N__57673),
            .in3(N__53116),
            .lcout(n20502),
            .ltout(n20502_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15112_2_lut_LC_20_11_1.C_ON=1'b0;
    defparam i15112_2_lut_LC_20_11_1.SEQ_MODE=4'b0000;
    defparam i15112_2_lut_LC_20_11_1.LUT_INIT=16'b1111000000000000;
    LogicCell40 i15112_2_lut_LC_20_11_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__53119),
            .in3(N__57588),
            .lcout(n10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i5_4_lut_adj_224_LC_20_11_2.C_ON=1'b0;
    defparam i5_4_lut_adj_224_LC_20_11_2.SEQ_MODE=4'b0000;
    defparam i5_4_lut_adj_224_LC_20_11_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i5_4_lut_adj_224_LC_20_11_2 (
            .in0(N__57652),
            .in1(N__57616),
            .in2(N__57697),
            .in3(N__57634),
            .lcout(n12_adj_1583),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclk_294_LC_20_11_3.C_ON=1'b0;
    defparam dds0_mclk_294_LC_20_11_3.SEQ_MODE=4'b1000;
    defparam dds0_mclk_294_LC_20_11_3.LUT_INIT=16'b1010101001100110;
    LogicCell40 dds0_mclk_294_LC_20_11_3 (
            .in0(N__55977),
            .in1(N__57589),
            .in2(_gnd_net_),
            .in3(N__53110),
            .lcout(dds0_mclk),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVdds0_mclk_294C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam i6_4_lut_adj_226_LC_20_11_6.C_ON=1'b0;
    defparam i6_4_lut_adj_226_LC_20_11_6.SEQ_MODE=4'b0000;
    defparam i6_4_lut_adj_226_LC_20_11_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 i6_4_lut_adj_226_LC_20_11_6 (
            .in0(N__53104),
            .in1(N__53089),
            .in2(N__53074),
            .in3(N__53053),
            .lcout(n14_adj_1578),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18214_4_lut_LC_20_11_7.C_ON=1'b0;
    defparam i18214_4_lut_LC_20_11_7.SEQ_MODE=4'b0000;
    defparam i18214_4_lut_LC_20_11_7.LUT_INIT=16'b0111001001010000;
    LogicCell40 i18214_4_lut_LC_20_11_7 (
            .in0(N__57553),
            .in1(N__56978),
            .in2(N__56416),
            .in3(N__56401),
            .lcout(n20809),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15033_2_lut_LC_20_12_2.C_ON=1'b0;
    defparam i15033_2_lut_LC_20_12_2.SEQ_MODE=4'b0000;
    defparam i15033_2_lut_LC_20_12_2.LUT_INIT=16'b0011001100000000;
    LogicCell40 i15033_2_lut_LC_20_12_2 (
            .in0(_gnd_net_),
            .in1(N__54535),
            .in2(_gnd_net_),
            .in3(N__53371),
            .lcout(n17415),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_4_i30_3_lut_LC_20_13_2.C_ON=1'b0;
    defparam mux_130_Mux_4_i30_3_lut_LC_20_13_2.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_4_i30_3_lut_LC_20_13_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_130_Mux_4_i30_3_lut_LC_20_13_2 (
            .in0(N__56353),
            .in1(N__56310),
            .in2(_gnd_net_),
            .in3(N__56065),
            .lcout(n30_adj_1608),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_16MHz_I_0_3_lut_LC_20_14_1.C_ON=1'b0;
    defparam clk_16MHz_I_0_3_lut_LC_20_14_1.SEQ_MODE=4'b0000;
    defparam clk_16MHz_I_0_3_lut_LC_20_14_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 clk_16MHz_I_0_3_lut_LC_20_14_1 (
            .in0(N__56041),
            .in1(N__55981),
            .in2(_gnd_net_),
            .in3(N__55966),
            .lcout(DDS_MCLK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.SCLK_27_LC_20_17_0 .C_ON=1'b0;
    defparam \SIG_DDS.SCLK_27_LC_20_17_0 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.SCLK_27_LC_20_17_0 .LUT_INIT=16'b0011001010110001;
    LogicCell40 \SIG_DDS.SCLK_27_LC_20_17_0  (
            .in0(N__55744),
            .in1(N__55860),
            .in2(N__55905),
            .in3(N__55627),
            .lcout(DDS_SCK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55241),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.CS_28_LC_20_18_2 .C_ON=1'b0;
    defparam \SIG_DDS.CS_28_LC_20_18_2 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.CS_28_LC_20_18_2 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \SIG_DDS.CS_28_LC_20_18_2  (
            .in0(N__55861),
            .in1(N__55740),
            .in2(_gnd_net_),
            .in3(N__55626),
            .lcout(DDS_CS),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55244),
            .ce(N__55483),
            .sr(_gnd_net_));
    defparam comm_clear_301_LC_22_9_0.C_ON=1'b0;
    defparam comm_clear_301_LC_22_9_0.SEQ_MODE=4'b1000;
    defparam comm_clear_301_LC_22_9_0.LUT_INIT=16'b0111011100110011;
    LogicCell40 comm_clear_301_LC_22_9_0 (
            .in0(N__54561),
            .in1(N__54035),
            .in2(_gnd_net_),
            .in3(N__53486),
            .lcout(comm_clear),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55187),
            .ce(N__53266),
            .sr(_gnd_net_));
    defparam i2_2_lut_3_lut_adj_220_LC_22_10_2.C_ON=1'b0;
    defparam i2_2_lut_3_lut_adj_220_LC_22_10_2.SEQ_MODE=4'b0000;
    defparam i2_2_lut_3_lut_adj_220_LC_22_10_2.LUT_INIT=16'b1111111111011101;
    LogicCell40 i2_2_lut_3_lut_adj_220_LC_22_10_2 (
            .in0(N__54544),
            .in1(N__54034),
            .in2(_gnd_net_),
            .in3(N__53485),
            .lcout(n11347),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3772__i0_LC_22_11_0.C_ON=1'b1;
    defparam dds0_mclkcnt_i7_3772__i0_LC_22_11_0.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3772__i0_LC_22_11_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3772__i0_LC_22_11_0 (
            .in0(_gnd_net_),
            .in1(N__57714),
            .in2(_gnd_net_),
            .in3(N__57700),
            .lcout(dds0_mclkcnt_0),
            .ltout(),
            .carryin(bfn_22_11_0_),
            .carryout(n19440),
            .clk(INVdds0_mclkcnt_i7_3772__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3772__i1_LC_22_11_1.C_ON=1'b1;
    defparam dds0_mclkcnt_i7_3772__i1_LC_22_11_1.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3772__i1_LC_22_11_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3772__i1_LC_22_11_1 (
            .in0(_gnd_net_),
            .in1(N__57693),
            .in2(_gnd_net_),
            .in3(N__57676),
            .lcout(dds0_mclkcnt_1),
            .ltout(),
            .carryin(n19440),
            .carryout(n19441),
            .clk(INVdds0_mclkcnt_i7_3772__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3772__i2_LC_22_11_2.C_ON=1'b1;
    defparam dds0_mclkcnt_i7_3772__i2_LC_22_11_2.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3772__i2_LC_22_11_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3772__i2_LC_22_11_2 (
            .in0(_gnd_net_),
            .in1(N__57669),
            .in2(_gnd_net_),
            .in3(N__57655),
            .lcout(dds0_mclkcnt_2),
            .ltout(),
            .carryin(n19441),
            .carryout(n19442),
            .clk(INVdds0_mclkcnt_i7_3772__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3772__i3_LC_22_11_3.C_ON=1'b1;
    defparam dds0_mclkcnt_i7_3772__i3_LC_22_11_3.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3772__i3_LC_22_11_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3772__i3_LC_22_11_3 (
            .in0(_gnd_net_),
            .in1(N__57651),
            .in2(_gnd_net_),
            .in3(N__57637),
            .lcout(dds0_mclkcnt_3),
            .ltout(),
            .carryin(n19442),
            .carryout(n19443),
            .clk(INVdds0_mclkcnt_i7_3772__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3772__i4_LC_22_11_4.C_ON=1'b1;
    defparam dds0_mclkcnt_i7_3772__i4_LC_22_11_4.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3772__i4_LC_22_11_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3772__i4_LC_22_11_4 (
            .in0(_gnd_net_),
            .in1(N__57633),
            .in2(_gnd_net_),
            .in3(N__57619),
            .lcout(dds0_mclkcnt_4),
            .ltout(),
            .carryin(n19443),
            .carryout(n19444),
            .clk(INVdds0_mclkcnt_i7_3772__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3772__i5_LC_22_11_5.C_ON=1'b1;
    defparam dds0_mclkcnt_i7_3772__i5_LC_22_11_5.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3772__i5_LC_22_11_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3772__i5_LC_22_11_5 (
            .in0(_gnd_net_),
            .in1(N__57615),
            .in2(_gnd_net_),
            .in3(N__57601),
            .lcout(dds0_mclkcnt_5),
            .ltout(),
            .carryin(n19444),
            .carryout(n19445),
            .clk(INVdds0_mclkcnt_i7_3772__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3772__i6_LC_22_11_6.C_ON=1'b1;
    defparam dds0_mclkcnt_i7_3772__i6_LC_22_11_6.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3772__i6_LC_22_11_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3772__i6_LC_22_11_6 (
            .in0(_gnd_net_),
            .in1(N__57598),
            .in2(_gnd_net_),
            .in3(N__57574),
            .lcout(dds0_mclkcnt_6),
            .ltout(),
            .carryin(n19445),
            .carryout(n19446),
            .clk(INVdds0_mclkcnt_i7_3772__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3772__i7_LC_22_11_7.C_ON=1'b0;
    defparam dds0_mclkcnt_i7_3772__i7_LC_22_11_7.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3772__i7_LC_22_11_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3772__i7_LC_22_11_7 (
            .in0(_gnd_net_),
            .in1(N__57567),
            .in2(_gnd_net_),
            .in3(N__57571),
            .lcout(dds0_mclkcnt_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVdds0_mclkcnt_i7_3772__i0C_net),
            .ce(),
            .sr(_gnd_net_));
endmodule // zim
