-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jun 28 2024 10:36:39

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "vdc_gen_clk" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of vdc_gen_clk
entity vdc_gen_clk is
port (
    DIVIDE : in std_logic_vector(15 downto 0);
    ICLK : in std_logic;
    OCLK : out std_logic);
end vdc_gen_clk;

-- Architecture of vdc_gen_clk
-- View name is \INTERFACE\
architecture \INTERFACE\ of vdc_gen_clk is

signal \N__4245\ : std_logic;
signal \N__4244\ : std_logic;
signal \N__4243\ : std_logic;
signal \N__4236\ : std_logic;
signal \N__4235\ : std_logic;
signal \N__4234\ : std_logic;
signal \N__4227\ : std_logic;
signal \N__4226\ : std_logic;
signal \N__4225\ : std_logic;
signal \N__4218\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4216\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4208\ : std_logic;
signal \N__4207\ : std_logic;
signal \N__4200\ : std_logic;
signal \N__4199\ : std_logic;
signal \N__4198\ : std_logic;
signal \N__4191\ : std_logic;
signal \N__4190\ : std_logic;
signal \N__4189\ : std_logic;
signal \N__4182\ : std_logic;
signal \N__4181\ : std_logic;
signal \N__4180\ : std_logic;
signal \N__4173\ : std_logic;
signal \N__4172\ : std_logic;
signal \N__4171\ : std_logic;
signal \N__4164\ : std_logic;
signal \N__4163\ : std_logic;
signal \N__4162\ : std_logic;
signal \N__4155\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4153\ : std_logic;
signal \N__4146\ : std_logic;
signal \N__4145\ : std_logic;
signal \N__4144\ : std_logic;
signal \N__4137\ : std_logic;
signal \N__4136\ : std_logic;
signal \N__4135\ : std_logic;
signal \N__4128\ : std_logic;
signal \N__4127\ : std_logic;
signal \N__4126\ : std_logic;
signal \N__4119\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4117\ : std_logic;
signal \N__4110\ : std_logic;
signal \N__4109\ : std_logic;
signal \N__4108\ : std_logic;
signal \N__4101\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4099\ : std_logic;
signal \N__4092\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4090\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4072\ : std_logic;
signal \N__4069\ : std_logic;
signal \N__4066\ : std_logic;
signal \N__4063\ : std_logic;
signal \N__4060\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4054\ : std_logic;
signal \N__4051\ : std_logic;
signal \N__4048\ : std_logic;
signal \N__4043\ : std_logic;
signal \N__4040\ : std_logic;
signal \N__4039\ : std_logic;
signal \N__4036\ : std_logic;
signal \N__4033\ : std_logic;
signal \N__4030\ : std_logic;
signal \N__4025\ : std_logic;
signal \N__4022\ : std_logic;
signal \N__4019\ : std_logic;
signal \N__4018\ : std_logic;
signal \N__4015\ : std_logic;
signal \N__4012\ : std_logic;
signal \N__4009\ : std_logic;
signal \N__4004\ : std_logic;
signal \N__4001\ : std_logic;
signal \N__4000\ : std_logic;
signal \N__3997\ : std_logic;
signal \N__3994\ : std_logic;
signal \N__3991\ : std_logic;
signal \N__3986\ : std_logic;
signal \N__3985\ : std_logic;
signal \N__3982\ : std_logic;
signal \N__3979\ : std_logic;
signal \N__3974\ : std_logic;
signal \N__3971\ : std_logic;
signal \N__3968\ : std_logic;
signal \N__3965\ : std_logic;
signal \N__3964\ : std_logic;
signal \N__3961\ : std_logic;
signal \N__3958\ : std_logic;
signal \N__3955\ : std_logic;
signal \N__3950\ : std_logic;
signal \N__3947\ : std_logic;
signal \N__3946\ : std_logic;
signal \N__3943\ : std_logic;
signal \N__3940\ : std_logic;
signal \N__3937\ : std_logic;
signal \N__3932\ : std_logic;
signal \N__3931\ : std_logic;
signal \N__3928\ : std_logic;
signal \N__3925\ : std_logic;
signal \N__3922\ : std_logic;
signal \N__3917\ : std_logic;
signal \N__3914\ : std_logic;
signal \N__3911\ : std_logic;
signal \N__3908\ : std_logic;
signal \N__3905\ : std_logic;
signal \N__3902\ : std_logic;
signal \N__3899\ : std_logic;
signal \N__3896\ : std_logic;
signal \N__3893\ : std_logic;
signal \N__3890\ : std_logic;
signal \N__3889\ : std_logic;
signal \N__3886\ : std_logic;
signal \N__3883\ : std_logic;
signal \N__3880\ : std_logic;
signal \N__3877\ : std_logic;
signal \N__3872\ : std_logic;
signal \N__3869\ : std_logic;
signal \N__3866\ : std_logic;
signal \N__3863\ : std_logic;
signal \N__3860\ : std_logic;
signal \N__3857\ : std_logic;
signal \N__3854\ : std_logic;
signal \N__3851\ : std_logic;
signal \N__3848\ : std_logic;
signal \N__3847\ : std_logic;
signal \N__3844\ : std_logic;
signal \N__3841\ : std_logic;
signal \N__3836\ : std_logic;
signal \N__3833\ : std_logic;
signal \N__3830\ : std_logic;
signal \N__3827\ : std_logic;
signal \N__3824\ : std_logic;
signal \N__3823\ : std_logic;
signal \N__3822\ : std_logic;
signal \N__3821\ : std_logic;
signal \N__3820\ : std_logic;
signal \N__3819\ : std_logic;
signal \N__3818\ : std_logic;
signal \N__3817\ : std_logic;
signal \N__3816\ : std_logic;
signal \N__3815\ : std_logic;
signal \N__3814\ : std_logic;
signal \N__3813\ : std_logic;
signal \N__3812\ : std_logic;
signal \N__3811\ : std_logic;
signal \N__3798\ : std_logic;
signal \N__3795\ : std_logic;
signal \N__3782\ : std_logic;
signal \N__3781\ : std_logic;
signal \N__3780\ : std_logic;
signal \N__3777\ : std_logic;
signal \N__3774\ : std_logic;
signal \N__3771\ : std_logic;
signal \N__3768\ : std_logic;
signal \N__3763\ : std_logic;
signal \N__3762\ : std_logic;
signal \N__3759\ : std_logic;
signal \N__3758\ : std_logic;
signal \N__3757\ : std_logic;
signal \N__3756\ : std_logic;
signal \N__3755\ : std_logic;
signal \N__3754\ : std_logic;
signal \N__3751\ : std_logic;
signal \N__3744\ : std_logic;
signal \N__3741\ : std_logic;
signal \N__3738\ : std_logic;
signal \N__3727\ : std_logic;
signal \N__3716\ : std_logic;
signal \N__3713\ : std_logic;
signal \N__3710\ : std_logic;
signal \N__3707\ : std_logic;
signal \N__3704\ : std_logic;
signal \N__3703\ : std_logic;
signal \N__3700\ : std_logic;
signal \N__3697\ : std_logic;
signal \N__3692\ : std_logic;
signal \N__3691\ : std_logic;
signal \N__3690\ : std_logic;
signal \N__3689\ : std_logic;
signal \N__3688\ : std_logic;
signal \N__3685\ : std_logic;
signal \N__3682\ : std_logic;
signal \N__3681\ : std_logic;
signal \N__3680\ : std_logic;
signal \N__3679\ : std_logic;
signal \N__3678\ : std_logic;
signal \N__3677\ : std_logic;
signal \N__3676\ : std_logic;
signal \N__3675\ : std_logic;
signal \N__3672\ : std_logic;
signal \N__3669\ : std_logic;
signal \N__3666\ : std_logic;
signal \N__3661\ : std_logic;
signal \N__3658\ : std_logic;
signal \N__3655\ : std_logic;
signal \N__3652\ : std_logic;
signal \N__3649\ : std_logic;
signal \N__3648\ : std_logic;
signal \N__3645\ : std_logic;
signal \N__3642\ : std_logic;
signal \N__3639\ : std_logic;
signal \N__3636\ : std_logic;
signal \N__3631\ : std_logic;
signal \N__3626\ : std_logic;
signal \N__3623\ : std_logic;
signal \N__3618\ : std_logic;
signal \N__3615\ : std_logic;
signal \N__3614\ : std_logic;
signal \N__3611\ : std_logic;
signal \N__3606\ : std_logic;
signal \N__3603\ : std_logic;
signal \N__3600\ : std_logic;
signal \N__3597\ : std_logic;
signal \N__3594\ : std_logic;
signal \N__3589\ : std_logic;
signal \N__3586\ : std_logic;
signal \N__3581\ : std_logic;
signal \N__3568\ : std_logic;
signal \N__3565\ : std_logic;
signal \N__3562\ : std_logic;
signal \N__3559\ : std_logic;
signal \N__3556\ : std_logic;
signal \N__3553\ : std_logic;
signal \N__3550\ : std_logic;
signal \N__3545\ : std_logic;
signal \N__3542\ : std_logic;
signal \N__3541\ : std_logic;
signal \N__3540\ : std_logic;
signal \N__3537\ : std_logic;
signal \N__3534\ : std_logic;
signal \N__3533\ : std_logic;
signal \N__3530\ : std_logic;
signal \N__3529\ : std_logic;
signal \N__3524\ : std_logic;
signal \N__3521\ : std_logic;
signal \N__3518\ : std_logic;
signal \N__3515\ : std_logic;
signal \N__3510\ : std_logic;
signal \N__3505\ : std_logic;
signal \N__3502\ : std_logic;
signal \N__3499\ : std_logic;
signal \N__3494\ : std_logic;
signal \N__3491\ : std_logic;
signal \N__3488\ : std_logic;
signal \N__3485\ : std_logic;
signal \N__3482\ : std_logic;
signal \N__3479\ : std_logic;
signal \N__3476\ : std_logic;
signal \N__3473\ : std_logic;
signal \N__3470\ : std_logic;
signal \N__3467\ : std_logic;
signal \N__3464\ : std_logic;
signal \N__3461\ : std_logic;
signal \N__3458\ : std_logic;
signal \N__3455\ : std_logic;
signal \N__3452\ : std_logic;
signal \N__3449\ : std_logic;
signal \N__3446\ : std_logic;
signal \N__3443\ : std_logic;
signal \N__3440\ : std_logic;
signal \N__3437\ : std_logic;
signal \N__3434\ : std_logic;
signal \N__3431\ : std_logic;
signal \N__3428\ : std_logic;
signal \N__3425\ : std_logic;
signal \N__3422\ : std_logic;
signal \N__3419\ : std_logic;
signal \N__3416\ : std_logic;
signal \N__3413\ : std_logic;
signal \N__3412\ : std_logic;
signal \N__3411\ : std_logic;
signal \N__3408\ : std_logic;
signal \N__3407\ : std_logic;
signal \N__3406\ : std_logic;
signal \N__3403\ : std_logic;
signal \N__3402\ : std_logic;
signal \N__3399\ : std_logic;
signal \N__3398\ : std_logic;
signal \N__3395\ : std_logic;
signal \N__3392\ : std_logic;
signal \N__3389\ : std_logic;
signal \N__3386\ : std_logic;
signal \N__3383\ : std_logic;
signal \N__3380\ : std_logic;
signal \N__3377\ : std_logic;
signal \N__3372\ : std_logic;
signal \N__3369\ : std_logic;
signal \N__3364\ : std_logic;
signal \N__3359\ : std_logic;
signal \N__3356\ : std_logic;
signal \N__3351\ : std_logic;
signal \N__3344\ : std_logic;
signal \N__3343\ : std_logic;
signal \N__3342\ : std_logic;
signal \N__3341\ : std_logic;
signal \N__3340\ : std_logic;
signal \N__3339\ : std_logic;
signal \N__3338\ : std_logic;
signal \N__3337\ : std_logic;
signal \N__3336\ : std_logic;
signal \N__3335\ : std_logic;
signal \N__3334\ : std_logic;
signal \N__3333\ : std_logic;
signal \N__3330\ : std_logic;
signal \N__3325\ : std_logic;
signal \N__3324\ : std_logic;
signal \N__3313\ : std_logic;
signal \N__3304\ : std_logic;
signal \N__3299\ : std_logic;
signal \N__3298\ : std_logic;
signal \N__3297\ : std_logic;
signal \N__3294\ : std_logic;
signal \N__3293\ : std_logic;
signal \N__3288\ : std_logic;
signal \N__3285\ : std_logic;
signal \N__3278\ : std_logic;
signal \N__3277\ : std_logic;
signal \N__3276\ : std_logic;
signal \N__3273\ : std_logic;
signal \N__3272\ : std_logic;
signal \N__3271\ : std_logic;
signal \N__3268\ : std_logic;
signal \N__3263\ : std_logic;
signal \N__3260\ : std_logic;
signal \N__3257\ : std_logic;
signal \N__3250\ : std_logic;
signal \N__3239\ : std_logic;
signal \N__3236\ : std_logic;
signal \N__3235\ : std_logic;
signal \N__3232\ : std_logic;
signal \N__3229\ : std_logic;
signal \N__3226\ : std_logic;
signal \N__3221\ : std_logic;
signal \N__3220\ : std_logic;
signal \N__3217\ : std_logic;
signal \N__3214\ : std_logic;
signal \N__3211\ : std_logic;
signal \N__3206\ : std_logic;
signal \N__3203\ : std_logic;
signal \N__3202\ : std_logic;
signal \N__3199\ : std_logic;
signal \N__3196\ : std_logic;
signal \N__3193\ : std_logic;
signal \N__3188\ : std_logic;
signal \N__3187\ : std_logic;
signal \N__3184\ : std_logic;
signal \N__3181\ : std_logic;
signal \N__3178\ : std_logic;
signal \N__3173\ : std_logic;
signal \N__3170\ : std_logic;
signal \N__3169\ : std_logic;
signal \N__3164\ : std_logic;
signal \N__3161\ : std_logic;
signal \N__3158\ : std_logic;
signal \N__3155\ : std_logic;
signal \N__3152\ : std_logic;
signal \N__3149\ : std_logic;
signal \N__3146\ : std_logic;
signal \N__3143\ : std_logic;
signal \N__3140\ : std_logic;
signal \N__3137\ : std_logic;
signal \N__3134\ : std_logic;
signal \N__3131\ : std_logic;
signal \N__3128\ : std_logic;
signal \N__3125\ : std_logic;
signal \N__3122\ : std_logic;
signal \N__3119\ : std_logic;
signal \N__3116\ : std_logic;
signal \N__3113\ : std_logic;
signal \N__3110\ : std_logic;
signal \N__3107\ : std_logic;
signal \N__3104\ : std_logic;
signal \N__3101\ : std_logic;
signal \N__3098\ : std_logic;
signal \N__3095\ : std_logic;
signal \N__3092\ : std_logic;
signal \N__3089\ : std_logic;
signal \N__3086\ : std_logic;
signal \N__3083\ : std_logic;
signal \N__3080\ : std_logic;
signal \N__3077\ : std_logic;
signal \N__3074\ : std_logic;
signal \N__3071\ : std_logic;
signal \N__3068\ : std_logic;
signal \N__3065\ : std_logic;
signal \N__3062\ : std_logic;
signal \N__3059\ : std_logic;
signal \N__3056\ : std_logic;
signal \N__3053\ : std_logic;
signal \N__3050\ : std_logic;
signal \N__3047\ : std_logic;
signal \N__3044\ : std_logic;
signal \N__3041\ : std_logic;
signal \N__3038\ : std_logic;
signal \N__3035\ : std_logic;
signal \N__3032\ : std_logic;
signal \N__3029\ : std_logic;
signal \N__3026\ : std_logic;
signal \N__3023\ : std_logic;
signal \N__3020\ : std_logic;
signal \N__3019\ : std_logic;
signal \N__3016\ : std_logic;
signal \N__3013\ : std_logic;
signal \N__3008\ : std_logic;
signal \N__3007\ : std_logic;
signal \N__3004\ : std_logic;
signal \N__3001\ : std_logic;
signal \N__2998\ : std_logic;
signal \N__2995\ : std_logic;
signal \N__2994\ : std_logic;
signal \N__2991\ : std_logic;
signal \N__2988\ : std_logic;
signal \N__2985\ : std_logic;
signal \N__2978\ : std_logic;
signal \N__2975\ : std_logic;
signal \N__2972\ : std_logic;
signal \N__2969\ : std_logic;
signal \N__2968\ : std_logic;
signal \N__2965\ : std_logic;
signal \N__2962\ : std_logic;
signal \N__2957\ : std_logic;
signal \N__2956\ : std_logic;
signal \N__2953\ : std_logic;
signal \N__2950\ : std_logic;
signal \N__2945\ : std_logic;
signal \N__2944\ : std_logic;
signal \N__2941\ : std_logic;
signal \N__2938\ : std_logic;
signal \N__2933\ : std_logic;
signal \N__2930\ : std_logic;
signal \N__2927\ : std_logic;
signal \N__2924\ : std_logic;
signal \N__2921\ : std_logic;
signal \N__2918\ : std_logic;
signal \N__2917\ : std_logic;
signal \N__2912\ : std_logic;
signal \N__2909\ : std_logic;
signal \N__2908\ : std_logic;
signal \N__2905\ : std_logic;
signal \N__2902\ : std_logic;
signal \N__2897\ : std_logic;
signal \N__2894\ : std_logic;
signal \N__2891\ : std_logic;
signal \N__2888\ : std_logic;
signal \N__2885\ : std_logic;
signal \N__2882\ : std_logic;
signal \N__2879\ : std_logic;
signal \N__2876\ : std_logic;
signal \N__2873\ : std_logic;
signal \N__2870\ : std_logic;
signal \N__2867\ : std_logic;
signal \N__2864\ : std_logic;
signal \N__2861\ : std_logic;
signal \N__2858\ : std_logic;
signal \N__2855\ : std_logic;
signal \N__2852\ : std_logic;
signal \N__2849\ : std_logic;
signal \N__2846\ : std_logic;
signal \N__2843\ : std_logic;
signal \N__2840\ : std_logic;
signal \N__2837\ : std_logic;
signal \N__2834\ : std_logic;
signal \N__2831\ : std_logic;
signal \N__2828\ : std_logic;
signal \N__2825\ : std_logic;
signal \N__2822\ : std_logic;
signal \N__2819\ : std_logic;
signal \N__2816\ : std_logic;
signal \N__2813\ : std_logic;
signal \N__2810\ : std_logic;
signal \N__2809\ : std_logic;
signal \N__2808\ : std_logic;
signal \N__2807\ : std_logic;
signal \N__2806\ : std_logic;
signal \N__2805\ : std_logic;
signal \N__2804\ : std_logic;
signal \N__2801\ : std_logic;
signal \N__2798\ : std_logic;
signal \N__2795\ : std_logic;
signal \N__2794\ : std_logic;
signal \N__2791\ : std_logic;
signal \N__2788\ : std_logic;
signal \N__2785\ : std_logic;
signal \N__2784\ : std_logic;
signal \N__2783\ : std_logic;
signal \N__2782\ : std_logic;
signal \N__2781\ : std_logic;
signal \N__2780\ : std_logic;
signal \N__2779\ : std_logic;
signal \N__2778\ : std_logic;
signal \N__2777\ : std_logic;
signal \N__2776\ : std_logic;
signal \N__2775\ : std_logic;
signal \N__2774\ : std_logic;
signal \N__2773\ : std_logic;
signal \N__2772\ : std_logic;
signal \N__2771\ : std_logic;
signal \N__2770\ : std_logic;
signal \N__2769\ : std_logic;
signal \N__2768\ : std_logic;
signal \N__2761\ : std_logic;
signal \N__2750\ : std_logic;
signal \N__2747\ : std_logic;
signal \N__2744\ : std_logic;
signal \N__2741\ : std_logic;
signal \N__2738\ : std_logic;
signal \N__2735\ : std_logic;
signal \N__2732\ : std_logic;
signal \N__2729\ : std_logic;
signal \N__2728\ : std_logic;
signal \N__2725\ : std_logic;
signal \N__2724\ : std_logic;
signal \N__2721\ : std_logic;
signal \N__2720\ : std_logic;
signal \N__2717\ : std_logic;
signal \N__2716\ : std_logic;
signal \N__2713\ : std_logic;
signal \N__2710\ : std_logic;
signal \N__2709\ : std_logic;
signal \N__2706\ : std_logic;
signal \N__2703\ : std_logic;
signal \N__2700\ : std_logic;
signal \N__2697\ : std_logic;
signal \N__2694\ : std_logic;
signal \N__2689\ : std_logic;
signal \N__2682\ : std_logic;
signal \N__2673\ : std_logic;
signal \N__2656\ : std_logic;
signal \N__2647\ : std_logic;
signal \N__2640\ : std_logic;
signal \N__2627\ : std_logic;
signal \N__2624\ : std_logic;
signal \N__2621\ : std_logic;
signal \N__2618\ : std_logic;
signal \N__2615\ : std_logic;
signal \N__2612\ : std_logic;
signal \N__2609\ : std_logic;
signal \N__2608\ : std_logic;
signal \N__2607\ : std_logic;
signal \N__2604\ : std_logic;
signal \N__2601\ : std_logic;
signal \N__2598\ : std_logic;
signal \N__2595\ : std_logic;
signal \N__2592\ : std_logic;
signal \N__2587\ : std_logic;
signal \N__2584\ : std_logic;
signal \N__2581\ : std_logic;
signal \N__2578\ : std_logic;
signal \N__2575\ : std_logic;
signal \N__2572\ : std_logic;
signal \N__2567\ : std_logic;
signal \N__2564\ : std_logic;
signal \N__2561\ : std_logic;
signal \N__2560\ : std_logic;
signal \N__2557\ : std_logic;
signal \N__2554\ : std_logic;
signal \N__2549\ : std_logic;
signal \N__2548\ : std_logic;
signal \N__2545\ : std_logic;
signal \N__2544\ : std_logic;
signal \N__2541\ : std_logic;
signal \N__2538\ : std_logic;
signal \N__2535\ : std_logic;
signal \N__2532\ : std_logic;
signal \N__2527\ : std_logic;
signal \N__2524\ : std_logic;
signal \N__2521\ : std_logic;
signal \N__2516\ : std_logic;
signal \N__2513\ : std_logic;
signal \N__2510\ : std_logic;
signal \N__2507\ : std_logic;
signal \N__2506\ : std_logic;
signal \N__2503\ : std_logic;
signal \N__2500\ : std_logic;
signal \N__2495\ : std_logic;
signal \N__2492\ : std_logic;
signal \N__2491\ : std_logic;
signal \N__2490\ : std_logic;
signal \N__2487\ : std_logic;
signal \N__2484\ : std_logic;
signal \N__2481\ : std_logic;
signal \N__2476\ : std_logic;
signal \N__2473\ : std_logic;
signal \N__2470\ : std_logic;
signal \N__2467\ : std_logic;
signal \N__2464\ : std_logic;
signal \N__2461\ : std_logic;
signal \N__2458\ : std_logic;
signal \N__2453\ : std_logic;
signal \N__2450\ : std_logic;
signal \N__2447\ : std_logic;
signal \N__2446\ : std_logic;
signal \N__2443\ : std_logic;
signal \N__2440\ : std_logic;
signal \N__2435\ : std_logic;
signal \N__2434\ : std_logic;
signal \N__2433\ : std_logic;
signal \N__2430\ : std_logic;
signal \N__2427\ : std_logic;
signal \N__2424\ : std_logic;
signal \N__2421\ : std_logic;
signal \N__2416\ : std_logic;
signal \N__2413\ : std_logic;
signal \N__2410\ : std_logic;
signal \N__2407\ : std_logic;
signal \N__2404\ : std_logic;
signal \N__2401\ : std_logic;
signal \N__2398\ : std_logic;
signal \N__2393\ : std_logic;
signal \N__2390\ : std_logic;
signal \N__2387\ : std_logic;
signal \N__2386\ : std_logic;
signal \N__2383\ : std_logic;
signal \N__2380\ : std_logic;
signal \N__2377\ : std_logic;
signal \N__2372\ : std_logic;
signal \N__2371\ : std_logic;
signal \N__2368\ : std_logic;
signal \N__2365\ : std_logic;
signal \N__2362\ : std_logic;
signal \N__2357\ : std_logic;
signal \N__2354\ : std_logic;
signal \N__2351\ : std_logic;
signal \N__2348\ : std_logic;
signal \N__2345\ : std_logic;
signal \N__2344\ : std_logic;
signal \N__2341\ : std_logic;
signal \N__2338\ : std_logic;
signal \N__2333\ : std_logic;
signal \N__2330\ : std_logic;
signal \N__2327\ : std_logic;
signal \N__2324\ : std_logic;
signal \N__2321\ : std_logic;
signal \N__2318\ : std_logic;
signal \N__2315\ : std_logic;
signal \N__2312\ : std_logic;
signal \N__2309\ : std_logic;
signal \N__2306\ : std_logic;
signal \N__2303\ : std_logic;
signal \N__2300\ : std_logic;
signal \N__2297\ : std_logic;
signal \N__2296\ : std_logic;
signal \N__2293\ : std_logic;
signal \N__2290\ : std_logic;
signal \N__2285\ : std_logic;
signal \N__2282\ : std_logic;
signal \N__2279\ : std_logic;
signal \N__2276\ : std_logic;
signal \N__2273\ : std_logic;
signal \N__2270\ : std_logic;
signal \N__2267\ : std_logic;
signal \N__2264\ : std_logic;
signal \N__2261\ : std_logic;
signal \N__2258\ : std_logic;
signal \N__2255\ : std_logic;
signal \N__2254\ : std_logic;
signal \N__2251\ : std_logic;
signal \N__2248\ : std_logic;
signal \N__2245\ : std_logic;
signal \N__2240\ : std_logic;
signal \N__2237\ : std_logic;
signal \N__2234\ : std_logic;
signal \N__2231\ : std_logic;
signal \N__2230\ : std_logic;
signal \N__2227\ : std_logic;
signal \N__2224\ : std_logic;
signal \N__2221\ : std_logic;
signal \N__2218\ : std_logic;
signal \N__2213\ : std_logic;
signal \N__2210\ : std_logic;
signal \N__2207\ : std_logic;
signal \N__2204\ : std_logic;
signal \N__2203\ : std_logic;
signal \N__2200\ : std_logic;
signal \N__2197\ : std_logic;
signal \N__2192\ : std_logic;
signal \N__2189\ : std_logic;
signal \N__2186\ : std_logic;
signal \N__2183\ : std_logic;
signal \N__2180\ : std_logic;
signal \N__2179\ : std_logic;
signal \N__2176\ : std_logic;
signal \N__2173\ : std_logic;
signal \N__2168\ : std_logic;
signal \N__2165\ : std_logic;
signal \N__2162\ : std_logic;
signal \N__2159\ : std_logic;
signal \N__2156\ : std_logic;
signal \N__2153\ : std_logic;
signal \N__2150\ : std_logic;
signal \N__2147\ : std_logic;
signal \N__2144\ : std_logic;
signal \N__2143\ : std_logic;
signal \N__2140\ : std_logic;
signal \N__2137\ : std_logic;
signal \N__2136\ : std_logic;
signal \N__2133\ : std_logic;
signal \N__2130\ : std_logic;
signal \N__2127\ : std_logic;
signal \N__2122\ : std_logic;
signal \N__2119\ : std_logic;
signal \N__2116\ : std_logic;
signal \N__2113\ : std_logic;
signal \N__2108\ : std_logic;
signal \N__2105\ : std_logic;
signal \N__2102\ : std_logic;
signal \N__2099\ : std_logic;
signal \N__2096\ : std_logic;
signal \N__2093\ : std_logic;
signal \N__2090\ : std_logic;
signal \N__2089\ : std_logic;
signal \N__2086\ : std_logic;
signal \N__2083\ : std_logic;
signal \N__2082\ : std_logic;
signal \N__2079\ : std_logic;
signal \N__2076\ : std_logic;
signal \N__2073\ : std_logic;
signal \N__2070\ : std_logic;
signal \N__2065\ : std_logic;
signal \N__2060\ : std_logic;
signal \N__2057\ : std_logic;
signal \N__2056\ : std_logic;
signal \N__2053\ : std_logic;
signal \N__2050\ : std_logic;
signal \N__2049\ : std_logic;
signal \N__2046\ : std_logic;
signal \N__2043\ : std_logic;
signal \N__2040\ : std_logic;
signal \N__2033\ : std_logic;
signal \N__2030\ : std_logic;
signal \N__2027\ : std_logic;
signal \N__2026\ : std_logic;
signal \N__2023\ : std_logic;
signal \N__2020\ : std_logic;
signal \N__2015\ : std_logic;
signal \N__2012\ : std_logic;
signal \N__2009\ : std_logic;
signal \N__2006\ : std_logic;
signal \N__2005\ : std_logic;
signal \N__2002\ : std_logic;
signal \N__1999\ : std_logic;
signal \N__1994\ : std_logic;
signal \N__1991\ : std_logic;
signal \N__1988\ : std_logic;
signal \N__1985\ : std_logic;
signal \N__1982\ : std_logic;
signal \N__1981\ : std_logic;
signal \N__1978\ : std_logic;
signal \N__1975\ : std_logic;
signal \N__1970\ : std_logic;
signal \N__1967\ : std_logic;
signal \N__1964\ : std_logic;
signal \N__1961\ : std_logic;
signal \N__1958\ : std_logic;
signal \N__1955\ : std_logic;
signal \N__1952\ : std_logic;
signal \N__1949\ : std_logic;
signal \N__1946\ : std_logic;
signal \N__1943\ : std_logic;
signal \N__1940\ : std_logic;
signal \N__1937\ : std_logic;
signal \N__1934\ : std_logic;
signal \N__1931\ : std_logic;
signal \N__1928\ : std_logic;
signal \N__1927\ : std_logic;
signal \N__1926\ : std_logic;
signal \N__1923\ : std_logic;
signal \N__1920\ : std_logic;
signal \N__1917\ : std_logic;
signal \N__1910\ : std_logic;
signal \N__1907\ : std_logic;
signal \N__1904\ : std_logic;
signal \N__1901\ : std_logic;
signal \N__1898\ : std_logic;
signal \N__1895\ : std_logic;
signal \N__1892\ : std_logic;
signal \N__1889\ : std_logic;
signal \N__1886\ : std_logic;
signal \N__1883\ : std_logic;
signal \N__1880\ : std_logic;
signal \N__1877\ : std_logic;
signal \N__1874\ : std_logic;
signal \N__1871\ : std_logic;
signal \N__1868\ : std_logic;
signal \N__1865\ : std_logic;
signal \N__1862\ : std_logic;
signal \N__1859\ : std_logic;
signal \N__1858\ : std_logic;
signal \N__1855\ : std_logic;
signal \N__1852\ : std_logic;
signal \N__1851\ : std_logic;
signal \N__1846\ : std_logic;
signal \N__1843\ : std_logic;
signal \N__1838\ : std_logic;
signal \N__1835\ : std_logic;
signal \N__1832\ : std_logic;
signal \N__1829\ : std_logic;
signal \N__1826\ : std_logic;
signal \N__1823\ : std_logic;
signal \N__1820\ : std_logic;
signal \N__1817\ : std_logic;
signal \N__1814\ : std_logic;
signal \N__1811\ : std_logic;
signal \N__1808\ : std_logic;
signal \N__1805\ : std_logic;
signal \N__1802\ : std_logic;
signal \N__1799\ : std_logic;
signal \N__1798\ : std_logic;
signal \N__1797\ : std_logic;
signal \N__1794\ : std_logic;
signal \N__1791\ : std_logic;
signal \N__1788\ : std_logic;
signal \N__1781\ : std_logic;
signal \N__1778\ : std_logic;
signal \N__1775\ : std_logic;
signal \N__1772\ : std_logic;
signal \N__1769\ : std_logic;
signal \N__1766\ : std_logic;
signal \N__1763\ : std_logic;
signal \N__1762\ : std_logic;
signal \N__1759\ : std_logic;
signal \N__1756\ : std_logic;
signal \N__1751\ : std_logic;
signal \N__1750\ : std_logic;
signal \N__1747\ : std_logic;
signal \N__1744\ : std_logic;
signal \N__1739\ : std_logic;
signal \N__1736\ : std_logic;
signal \N__1733\ : std_logic;
signal \N__1730\ : std_logic;
signal \N__1727\ : std_logic;
signal \N__1724\ : std_logic;
signal \N__1721\ : std_logic;
signal \N__1718\ : std_logic;
signal \N__1715\ : std_logic;
signal \N__1712\ : std_logic;
signal \N__1709\ : std_logic;
signal \N__1706\ : std_logic;
signal \N__1703\ : std_logic;
signal \N__1700\ : std_logic;
signal \N__1699\ : std_logic;
signal \N__1698\ : std_logic;
signal \N__1695\ : std_logic;
signal \N__1692\ : std_logic;
signal \N__1689\ : std_logic;
signal \N__1686\ : std_logic;
signal \N__1681\ : std_logic;
signal \N__1678\ : std_logic;
signal \N__1675\ : std_logic;
signal \N__1670\ : std_logic;
signal \N__1667\ : std_logic;
signal \N__1664\ : std_logic;
signal \N__1661\ : std_logic;
signal \N__1658\ : std_logic;
signal \N__1655\ : std_logic;
signal \N__1652\ : std_logic;
signal \N__1649\ : std_logic;
signal \N__1646\ : std_logic;
signal \N__1643\ : std_logic;
signal \N__1640\ : std_logic;
signal \N__1637\ : std_logic;
signal \N__1634\ : std_logic;
signal \N__1631\ : std_logic;
signal \N__1628\ : std_logic;
signal \N__1625\ : std_logic;
signal \N__1622\ : std_logic;
signal \N__1619\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \DIVIDE_0_\ : std_logic;
signal \bfn_1_9_0_\ : std_logic;
signal n16 : std_logic;
signal n418 : std_logic;
signal n15 : std_logic;
signal n419 : std_logic;
signal n14 : std_logic;
signal n420 : std_logic;
signal n13 : std_logic;
signal \DIVIDE_4_\ : std_logic;
signal n421 : std_logic;
signal \DIVIDE_5_\ : std_logic;
signal n422 : std_logic;
signal n11 : std_logic;
signal n423 : std_logic;
signal n424 : std_logic;
signal n425 : std_logic;
signal n9 : std_logic;
signal \bfn_1_10_0_\ : std_logic;
signal \DIVIDE_9_\ : std_logic;
signal n426 : std_logic;
signal n427 : std_logic;
signal n428 : std_logic;
signal n5 : std_logic;
signal n429 : std_logic;
signal n4 : std_logic;
signal n430 : std_logic;
signal \DIVIDE_14_\ : std_logic;
signal n431 : std_logic;
signal n432 : std_logic;
signal n7 : std_logic;
signal \OCLK\ : std_logic;
signal n10 : std_logic;
signal \DIVIDE_6_\ : std_logic;
signal n12 : std_logic;
signal n3 : std_logic;
signal \DIVIDE_1_\ : std_logic;
signal n17 : std_logic;
signal \DIVIDE_7_\ : std_logic;
signal \DIVIDE_2_\ : std_logic;
signal t0on_0 : std_logic;
signal \t0on_15_N_35_0\ : std_logic;
signal \bfn_2_7_0_\ : std_logic;
signal t0on_1 : std_logic;
signal \t0on_15_N_35_1\ : std_logic;
signal n403 : std_logic;
signal n404 : std_logic;
signal t0on_3 : std_logic;
signal \t0on_15_N_35_3\ : std_logic;
signal n405 : std_logic;
signal t0on_4 : std_logic;
signal \t0on_15_N_35_4\ : std_logic;
signal n406 : std_logic;
signal t0on_5 : std_logic;
signal \t0on_15_N_35_5\ : std_logic;
signal n407 : std_logic;
signal t0on_6 : std_logic;
signal \t0on_15_N_35_6\ : std_logic;
signal n408 : std_logic;
signal n409 : std_logic;
signal n410 : std_logic;
signal t0on_8 : std_logic;
signal \t0on_15_N_35_8\ : std_logic;
signal \bfn_2_8_0_\ : std_logic;
signal n411 : std_logic;
signal n412 : std_logic;
signal n413 : std_logic;
signal n414 : std_logic;
signal t0on_13 : std_logic;
signal \t0on_15_N_35_13\ : std_logic;
signal n415 : std_logic;
signal n416 : std_logic;
signal n417 : std_logic;
signal \bfn_2_9_0_\ : std_logic;
signal n388 : std_logic;
signal n389 : std_logic;
signal n390 : std_logic;
signal n391 : std_logic;
signal n392 : std_logic;
signal n393 : std_logic;
signal n394 : std_logic;
signal n395 : std_logic;
signal \bfn_2_10_0_\ : std_logic;
signal n396 : std_logic;
signal n397 : std_logic;
signal n398 : std_logic;
signal n399 : std_logic;
signal n400 : std_logic;
signal n401 : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal n402 : std_logic;
signal \t0off_15_N_51_15\ : std_logic;
signal \DIVIDE_11_\ : std_logic;
signal \t0on_15_N_35_10\ : std_logic;
signal t0on_10 : std_logic;
signal \DIVIDE_3_\ : std_logic;
signal \t0on_15_N_35_2\ : std_logic;
signal t0on_2 : std_logic;
signal \DIVIDE_13_\ : std_logic;
signal \t0on_15_N_35_12\ : std_logic;
signal t0on_12 : std_logic;
signal \DIVIDE_8_\ : std_logic;
signal \t0on_15_N_35_7\ : std_logic;
signal t0on_7 : std_logic;
signal t0on_15 : std_logic;
signal \t0on_15_N_35_11\ : std_logic;
signal t0on_11 : std_logic;
signal \t0on_15_N_35_9\ : std_logic;
signal t0on_9 : std_logic;
signal \DIVIDE_15_\ : std_logic;
signal \t0on_15_N_35_14\ : std_logic;
signal t0on_14 : std_logic;
signal \DIVIDE_12_\ : std_logic;
signal n6 : std_logic;
signal \DIVIDE_10_\ : std_logic;
signal n8 : std_logic;
signal \t0off_15_N_67_3\ : std_logic;
signal \t0off_15_N_51_3\ : std_logic;
signal \t0off_15_N_67_8\ : std_logic;
signal \t0off_15_N_51_8\ : std_logic;
signal \t0off_15_N_67_2\ : std_logic;
signal \t0off_15_N_51_2\ : std_logic;
signal \t0off_15_N_67_10\ : std_logic;
signal \t0off_15_N_51_10\ : std_logic;
signal \t0off_15_N_67_13\ : std_logic;
signal \t0off_15_N_51_13\ : std_logic;
signal \t0off_15_N_67_7\ : std_logic;
signal \t0off_15_N_51_7\ : std_logic;
signal \t0off_15_N_67_12\ : std_logic;
signal \t0off_15_N_51_12\ : std_logic;
signal \t0off_15_N_51_9\ : std_logic;
signal \t0off_15_N_67_9\ : std_logic;
signal \t0off_15_N_67_14\ : std_logic;
signal \t0off_15_N_51_14\ : std_logic;
signal \t0off_15_N_67_4\ : std_logic;
signal \t0off_15_N_51_4\ : std_logic;
signal \t0off_15_N_67_1\ : std_logic;
signal \t0off_15_N_51_1\ : std_logic;
signal \t0off_15_N_67_0\ : std_logic;
signal \t0off_15_N_51_0\ : std_logic;
signal n26_adj_2 : std_logic;
signal n27_adj_18 : std_logic;
signal n28_adj_1 : std_logic;
signal n447 : std_logic;
signal \n441_cascade_\ : std_logic;
signal n6_adj_3 : std_logic;
signal n441 : std_logic;
signal n386 : std_logic;
signal \div_state_1__N_88\ : std_logic;
signal div_state_0 : std_logic;
signal t0off_12 : std_logic;
signal t0off_2 : std_logic;
signal t0off_7 : std_logic;
signal t0off_10 : std_logic;
signal \n27_cascade_\ : std_logic;
signal n442 : std_logic;
signal t0off_13 : std_logic;
signal t0off_3 : std_logic;
signal t0off_8 : std_logic;
signal n26 : std_logic;
signal t0off_14 : std_logic;
signal t0off_15 : std_logic;
signal t0off_9 : std_logic;
signal n28 : std_logic;
signal t0off_1 : std_logic;
signal t0off_4 : std_logic;
signal t0off_0 : std_logic;
signal n444 : std_logic;
signal \t0off_15_N_67_5\ : std_logic;
signal \t0off_15_N_51_5\ : std_logic;
signal t0off_5 : std_logic;
signal \t0off_15_N_67_6\ : std_logic;
signal \t0off_15_N_51_6\ : std_logic;
signal t0off_6 : std_logic;
signal \t0off_15_N_67_11\ : std_logic;
signal div_state_1 : std_logic;
signal \t0off_15_N_51_11\ : std_logic;
signal t0off_11 : std_logic;
signal \ICLK\ : std_logic;
signal n307 : std_logic;
signal \_gnd_net_\ : std_logic;

signal \DIVIDE_wire\ : std_logic_vector(15 downto 0);
signal \ICLK_wire\ : std_logic;
signal \OCLK_wire\ : std_logic;

begin
    \DIVIDE_wire\ <= DIVIDE;
    \ICLK_wire\ <= ICLK;
    OCLK <= \OCLK_wire\;

    \ipInertedIOPad_DIVIDE_c_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4245\,
            DIN => \N__4244\,
            DOUT => \N__4243\,
            PACKAGEPIN => \DIVIDE_wire\(2)
        );

    \ipInertedIOPad_DIVIDE_c_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__4245\,
            PADOUT => \N__4244\,
            PADIN => \N__4243\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \DIVIDE_2_\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DIVIDE_c_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4236\,
            DIN => \N__4235\,
            DOUT => \N__4234\,
            PACKAGEPIN => \DIVIDE_wire\(10)
        );

    \ipInertedIOPad_DIVIDE_c_10_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__4236\,
            PADOUT => \N__4235\,
            PADIN => \N__4234\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \DIVIDE_10_\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DIVIDE_c_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4227\,
            DIN => \N__4226\,
            DOUT => \N__4225\,
            PACKAGEPIN => \DIVIDE_wire\(9)
        );

    \ipInertedIOPad_DIVIDE_c_9_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__4227\,
            PADOUT => \N__4226\,
            PADIN => \N__4225\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \DIVIDE_9_\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DIVIDE_c_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4218\,
            DIN => \N__4217\,
            DOUT => \N__4216\,
            PACKAGEPIN => \DIVIDE_wire\(5)
        );

    \ipInertedIOPad_DIVIDE_c_5_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__4218\,
            PADOUT => \N__4217\,
            PADIN => \N__4216\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \DIVIDE_5_\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DIVIDE_c_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4209\,
            DIN => \N__4208\,
            DOUT => \N__4207\,
            PACKAGEPIN => \DIVIDE_wire\(15)
        );

    \ipInertedIOPad_DIVIDE_c_15_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__4209\,
            PADOUT => \N__4208\,
            PADIN => \N__4207\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \DIVIDE_15_\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DIVIDE_c_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4200\,
            DIN => \N__4199\,
            DOUT => \N__4198\,
            PACKAGEPIN => \DIVIDE_wire\(11)
        );

    \ipInertedIOPad_DIVIDE_c_11_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__4200\,
            PADOUT => \N__4199\,
            PADIN => \N__4198\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \DIVIDE_11_\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DIVIDE_c_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4191\,
            DIN => \N__4190\,
            DOUT => \N__4189\,
            PACKAGEPIN => \DIVIDE_wire\(1)
        );

    \ipInertedIOPad_DIVIDE_c_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__4191\,
            PADOUT => \N__4190\,
            PADIN => \N__4189\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \DIVIDE_1_\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_ICLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4182\,
            DIN => \N__4181\,
            DOUT => \N__4180\,
            PACKAGEPIN => \ICLK_wire\
        );

    \ipInertedIOPad_ICLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__4182\,
            PADOUT => \N__4181\,
            PADIN => \N__4180\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \ICLK\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DIVIDE_c_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4173\,
            DIN => \N__4172\,
            DOUT => \N__4171\,
            PACKAGEPIN => \DIVIDE_wire\(8)
        );

    \ipInertedIOPad_DIVIDE_c_8_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__4173\,
            PADOUT => \N__4172\,
            PADIN => \N__4171\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \DIVIDE_8_\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DIVIDE_c_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4164\,
            DIN => \N__4163\,
            DOUT => \N__4162\,
            PACKAGEPIN => \DIVIDE_wire\(4)
        );

    \ipInertedIOPad_DIVIDE_c_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__4164\,
            PADOUT => \N__4163\,
            PADIN => \N__4162\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \DIVIDE_4_\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DIVIDE_c_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4155\,
            DIN => \N__4154\,
            DOUT => \N__4153\,
            PACKAGEPIN => \DIVIDE_wire\(12)
        );

    \ipInertedIOPad_DIVIDE_c_12_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__4155\,
            PADOUT => \N__4154\,
            PADIN => \N__4153\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \DIVIDE_12_\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DIVIDE_c_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4146\,
            DIN => \N__4145\,
            DOUT => \N__4144\,
            PACKAGEPIN => \DIVIDE_wire\(0)
        );

    \ipInertedIOPad_DIVIDE_c_0_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__4146\,
            PADOUT => \N__4145\,
            PADIN => \N__4144\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \DIVIDE_0_\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_OCLK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4137\,
            DIN => \N__4136\,
            DOUT => \N__4135\,
            PACKAGEPIN => \OCLK_wire\
        );

    \ipInertedIOPad_OCLK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__4137\,
            PADOUT => \N__4136\,
            PADIN => \N__4135\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__1880\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DIVIDE_c_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4128\,
            DIN => \N__4127\,
            DOUT => \N__4126\,
            PACKAGEPIN => \DIVIDE_wire\(7)
        );

    \ipInertedIOPad_DIVIDE_c_7_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__4128\,
            PADOUT => \N__4127\,
            PADIN => \N__4126\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \DIVIDE_7_\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DIVIDE_c_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4119\,
            DIN => \N__4118\,
            DOUT => \N__4117\,
            PACKAGEPIN => \DIVIDE_wire\(3)
        );

    \ipInertedIOPad_DIVIDE_c_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__4119\,
            PADOUT => \N__4118\,
            PADIN => \N__4117\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \DIVIDE_3_\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DIVIDE_c_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4110\,
            DIN => \N__4109\,
            DOUT => \N__4108\,
            PACKAGEPIN => \DIVIDE_wire\(13)
        );

    \ipInertedIOPad_DIVIDE_c_13_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__4110\,
            PADOUT => \N__4109\,
            PADIN => \N__4108\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \DIVIDE_13_\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DIVIDE_c_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4101\,
            DIN => \N__4100\,
            DOUT => \N__4099\,
            PACKAGEPIN => \DIVIDE_wire\(6)
        );

    \ipInertedIOPad_DIVIDE_c_6_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__4101\,
            PADOUT => \N__4100\,
            PADIN => \N__4099\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \DIVIDE_6_\,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DIVIDE_c_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__4092\,
            DIN => \N__4091\,
            DOUT => \N__4090\,
            PACKAGEPIN => \DIVIDE_wire\(14)
        );

    \ipInertedIOPad_DIVIDE_c_14_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__4092\,
            PADOUT => \N__4091\,
            PADIN => \N__4090\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => \DIVIDE_14_\,
            DIN1 => OPEN
        );

    \I__956\ : CascadeMux
    port map (
            O => \N__4073\,
            I => \N__4069\
        );

    \I__955\ : InMux
    port map (
            O => \N__4072\,
            I => \N__4066\
        );

    \I__954\ : InMux
    port map (
            O => \N__4069\,
            I => \N__4063\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__4066\,
            I => \N__4060\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__4063\,
            I => t0off_13
        );

    \I__951\ : Odrv4
    port map (
            O => \N__4060\,
            I => t0off_13
        );

    \I__950\ : InMux
    port map (
            O => \N__4055\,
            I => \N__4051\
        );

    \I__949\ : InMux
    port map (
            O => \N__4054\,
            I => \N__4048\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__4051\,
            I => \N__4043\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__4048\,
            I => \N__4043\
        );

    \I__946\ : Odrv4
    port map (
            O => \N__4043\,
            I => t0off_3
        );

    \I__945\ : InMux
    port map (
            O => \N__4040\,
            I => \N__4036\
        );

    \I__944\ : InMux
    port map (
            O => \N__4039\,
            I => \N__4033\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__4036\,
            I => \N__4030\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__4033\,
            I => t0off_8
        );

    \I__941\ : Odrv4
    port map (
            O => \N__4030\,
            I => t0off_8
        );

    \I__940\ : InMux
    port map (
            O => \N__4025\,
            I => \N__4022\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__4022\,
            I => n26
        );

    \I__938\ : InMux
    port map (
            O => \N__4019\,
            I => \N__4015\
        );

    \I__937\ : InMux
    port map (
            O => \N__4018\,
            I => \N__4012\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__4015\,
            I => \N__4009\
        );

    \I__935\ : LocalMux
    port map (
            O => \N__4012\,
            I => t0off_14
        );

    \I__934\ : Odrv12
    port map (
            O => \N__4009\,
            I => t0off_14
        );

    \I__933\ : CascadeMux
    port map (
            O => \N__4004\,
            I => \N__4001\
        );

    \I__932\ : InMux
    port map (
            O => \N__4001\,
            I => \N__3997\
        );

    \I__931\ : InMux
    port map (
            O => \N__4000\,
            I => \N__3994\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__3997\,
            I => \N__3991\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__3994\,
            I => t0off_15
        );

    \I__928\ : Odrv12
    port map (
            O => \N__3991\,
            I => t0off_15
        );

    \I__927\ : InMux
    port map (
            O => \N__3986\,
            I => \N__3982\
        );

    \I__926\ : InMux
    port map (
            O => \N__3985\,
            I => \N__3979\
        );

    \I__925\ : LocalMux
    port map (
            O => \N__3982\,
            I => \N__3974\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__3979\,
            I => \N__3974\
        );

    \I__923\ : Odrv4
    port map (
            O => \N__3974\,
            I => t0off_9
        );

    \I__922\ : InMux
    port map (
            O => \N__3971\,
            I => \N__3968\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__3968\,
            I => n28
        );

    \I__920\ : InMux
    port map (
            O => \N__3965\,
            I => \N__3961\
        );

    \I__919\ : InMux
    port map (
            O => \N__3964\,
            I => \N__3958\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__3961\,
            I => \N__3955\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__3958\,
            I => t0off_1
        );

    \I__916\ : Odrv4
    port map (
            O => \N__3955\,
            I => t0off_1
        );

    \I__915\ : CascadeMux
    port map (
            O => \N__3950\,
            I => \N__3947\
        );

    \I__914\ : InMux
    port map (
            O => \N__3947\,
            I => \N__3943\
        );

    \I__913\ : InMux
    port map (
            O => \N__3946\,
            I => \N__3940\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__3943\,
            I => \N__3937\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__3940\,
            I => t0off_4
        );

    \I__910\ : Odrv4
    port map (
            O => \N__3937\,
            I => t0off_4
        );

    \I__909\ : InMux
    port map (
            O => \N__3932\,
            I => \N__3928\
        );

    \I__908\ : InMux
    port map (
            O => \N__3931\,
            I => \N__3925\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__3928\,
            I => \N__3922\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__3925\,
            I => t0off_0
        );

    \I__905\ : Odrv4
    port map (
            O => \N__3922\,
            I => t0off_0
        );

    \I__904\ : InMux
    port map (
            O => \N__3917\,
            I => \N__3914\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__3914\,
            I => n444
        );

    \I__902\ : InMux
    port map (
            O => \N__3911\,
            I => \N__3908\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__3908\,
            I => \N__3905\
        );

    \I__900\ : Odrv12
    port map (
            O => \N__3905\,
            I => \t0off_15_N_67_5\
        );

    \I__899\ : InMux
    port map (
            O => \N__3902\,
            I => \N__3899\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__3899\,
            I => \N__3896\
        );

    \I__897\ : Span4Mux_h
    port map (
            O => \N__3896\,
            I => \N__3893\
        );

    \I__896\ : Odrv4
    port map (
            O => \N__3893\,
            I => \t0off_15_N_51_5\
        );

    \I__895\ : InMux
    port map (
            O => \N__3890\,
            I => \N__3886\
        );

    \I__894\ : CascadeMux
    port map (
            O => \N__3889\,
            I => \N__3883\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__3886\,
            I => \N__3880\
        );

    \I__892\ : InMux
    port map (
            O => \N__3883\,
            I => \N__3877\
        );

    \I__891\ : Span4Mux_h
    port map (
            O => \N__3880\,
            I => \N__3872\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__3877\,
            I => \N__3872\
        );

    \I__889\ : Odrv4
    port map (
            O => \N__3872\,
            I => t0off_5
        );

    \I__888\ : InMux
    port map (
            O => \N__3869\,
            I => \N__3866\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__3866\,
            I => \N__3863\
        );

    \I__886\ : Odrv12
    port map (
            O => \N__3863\,
            I => \t0off_15_N_67_6\
        );

    \I__885\ : InMux
    port map (
            O => \N__3860\,
            I => \N__3857\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__3857\,
            I => \N__3854\
        );

    \I__883\ : Odrv12
    port map (
            O => \N__3854\,
            I => \t0off_15_N_51_6\
        );

    \I__882\ : InMux
    port map (
            O => \N__3851\,
            I => \N__3848\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__3848\,
            I => \N__3844\
        );

    \I__880\ : InMux
    port map (
            O => \N__3847\,
            I => \N__3841\
        );

    \I__879\ : Odrv12
    port map (
            O => \N__3844\,
            I => t0off_6
        );

    \I__878\ : LocalMux
    port map (
            O => \N__3841\,
            I => t0off_6
        );

    \I__877\ : InMux
    port map (
            O => \N__3836\,
            I => \N__3833\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__3833\,
            I => \N__3830\
        );

    \I__875\ : Span4Mux_h
    port map (
            O => \N__3830\,
            I => \N__3827\
        );

    \I__874\ : Odrv4
    port map (
            O => \N__3827\,
            I => \t0off_15_N_67_11\
        );

    \I__873\ : InMux
    port map (
            O => \N__3824\,
            I => \N__3798\
        );

    \I__872\ : InMux
    port map (
            O => \N__3823\,
            I => \N__3798\
        );

    \I__871\ : InMux
    port map (
            O => \N__3822\,
            I => \N__3798\
        );

    \I__870\ : InMux
    port map (
            O => \N__3821\,
            I => \N__3798\
        );

    \I__869\ : InMux
    port map (
            O => \N__3820\,
            I => \N__3798\
        );

    \I__868\ : InMux
    port map (
            O => \N__3819\,
            I => \N__3798\
        );

    \I__867\ : InMux
    port map (
            O => \N__3818\,
            I => \N__3795\
        );

    \I__866\ : InMux
    port map (
            O => \N__3817\,
            I => \N__3782\
        );

    \I__865\ : InMux
    port map (
            O => \N__3816\,
            I => \N__3782\
        );

    \I__864\ : InMux
    port map (
            O => \N__3815\,
            I => \N__3782\
        );

    \I__863\ : InMux
    port map (
            O => \N__3814\,
            I => \N__3782\
        );

    \I__862\ : InMux
    port map (
            O => \N__3813\,
            I => \N__3782\
        );

    \I__861\ : InMux
    port map (
            O => \N__3812\,
            I => \N__3782\
        );

    \I__860\ : InMux
    port map (
            O => \N__3811\,
            I => \N__3777\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__3798\,
            I => \N__3774\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__3795\,
            I => \N__3771\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__3782\,
            I => \N__3768\
        );

    \I__856\ : InMux
    port map (
            O => \N__3781\,
            I => \N__3763\
        );

    \I__855\ : InMux
    port map (
            O => \N__3780\,
            I => \N__3763\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__3777\,
            I => \N__3759\
        );

    \I__853\ : Span4Mux_v
    port map (
            O => \N__3774\,
            I => \N__3751\
        );

    \I__852\ : Span4Mux_v
    port map (
            O => \N__3771\,
            I => \N__3744\
        );

    \I__851\ : Span4Mux_h
    port map (
            O => \N__3768\,
            I => \N__3744\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__3763\,
            I => \N__3744\
        );

    \I__849\ : InMux
    port map (
            O => \N__3762\,
            I => \N__3741\
        );

    \I__848\ : Span12Mux_v
    port map (
            O => \N__3759\,
            I => \N__3738\
        );

    \I__847\ : InMux
    port map (
            O => \N__3758\,
            I => \N__3727\
        );

    \I__846\ : InMux
    port map (
            O => \N__3757\,
            I => \N__3727\
        );

    \I__845\ : InMux
    port map (
            O => \N__3756\,
            I => \N__3727\
        );

    \I__844\ : InMux
    port map (
            O => \N__3755\,
            I => \N__3727\
        );

    \I__843\ : InMux
    port map (
            O => \N__3754\,
            I => \N__3727\
        );

    \I__842\ : Odrv4
    port map (
            O => \N__3751\,
            I => div_state_1
        );

    \I__841\ : Odrv4
    port map (
            O => \N__3744\,
            I => div_state_1
        );

    \I__840\ : LocalMux
    port map (
            O => \N__3741\,
            I => div_state_1
        );

    \I__839\ : Odrv12
    port map (
            O => \N__3738\,
            I => div_state_1
        );

    \I__838\ : LocalMux
    port map (
            O => \N__3727\,
            I => div_state_1
        );

    \I__837\ : InMux
    port map (
            O => \N__3716\,
            I => \N__3713\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__3713\,
            I => \N__3710\
        );

    \I__835\ : Odrv12
    port map (
            O => \N__3710\,
            I => \t0off_15_N_51_11\
        );

    \I__834\ : InMux
    port map (
            O => \N__3707\,
            I => \N__3704\
        );

    \I__833\ : LocalMux
    port map (
            O => \N__3704\,
            I => \N__3700\
        );

    \I__832\ : InMux
    port map (
            O => \N__3703\,
            I => \N__3697\
        );

    \I__831\ : Odrv12
    port map (
            O => \N__3700\,
            I => t0off_11
        );

    \I__830\ : LocalMux
    port map (
            O => \N__3697\,
            I => t0off_11
        );

    \I__829\ : ClkMux
    port map (
            O => \N__3692\,
            I => \N__3685\
        );

    \I__828\ : ClkMux
    port map (
            O => \N__3691\,
            I => \N__3682\
        );

    \I__827\ : ClkMux
    port map (
            O => \N__3690\,
            I => \N__3672\
        );

    \I__826\ : ClkMux
    port map (
            O => \N__3689\,
            I => \N__3669\
        );

    \I__825\ : ClkMux
    port map (
            O => \N__3688\,
            I => \N__3666\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__3685\,
            I => \N__3661\
        );

    \I__823\ : LocalMux
    port map (
            O => \N__3682\,
            I => \N__3661\
        );

    \I__822\ : ClkMux
    port map (
            O => \N__3681\,
            I => \N__3658\
        );

    \I__821\ : ClkMux
    port map (
            O => \N__3680\,
            I => \N__3655\
        );

    \I__820\ : ClkMux
    port map (
            O => \N__3679\,
            I => \N__3652\
        );

    \I__819\ : ClkMux
    port map (
            O => \N__3678\,
            I => \N__3649\
        );

    \I__818\ : ClkMux
    port map (
            O => \N__3677\,
            I => \N__3645\
        );

    \I__817\ : ClkMux
    port map (
            O => \N__3676\,
            I => \N__3642\
        );

    \I__816\ : ClkMux
    port map (
            O => \N__3675\,
            I => \N__3639\
        );

    \I__815\ : LocalMux
    port map (
            O => \N__3672\,
            I => \N__3636\
        );

    \I__814\ : LocalMux
    port map (
            O => \N__3669\,
            I => \N__3631\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__3666\,
            I => \N__3631\
        );

    \I__812\ : Span4Mux_h
    port map (
            O => \N__3661\,
            I => \N__3626\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__3658\,
            I => \N__3626\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__3655\,
            I => \N__3623\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__3652\,
            I => \N__3618\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__3649\,
            I => \N__3618\
        );

    \I__807\ : ClkMux
    port map (
            O => \N__3648\,
            I => \N__3615\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__3645\,
            I => \N__3611\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__3642\,
            I => \N__3606\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__3639\,
            I => \N__3606\
        );

    \I__803\ : Span4Mux_v
    port map (
            O => \N__3636\,
            I => \N__3603\
        );

    \I__802\ : Span4Mux_v
    port map (
            O => \N__3631\,
            I => \N__3600\
        );

    \I__801\ : Span4Mux_v
    port map (
            O => \N__3626\,
            I => \N__3597\
        );

    \I__800\ : Span4Mux_v
    port map (
            O => \N__3623\,
            I => \N__3594\
        );

    \I__799\ : Span4Mux_v
    port map (
            O => \N__3618\,
            I => \N__3589\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__3615\,
            I => \N__3589\
        );

    \I__797\ : ClkMux
    port map (
            O => \N__3614\,
            I => \N__3586\
        );

    \I__796\ : Span4Mux_v
    port map (
            O => \N__3611\,
            I => \N__3581\
        );

    \I__795\ : Span4Mux_v
    port map (
            O => \N__3606\,
            I => \N__3581\
        );

    \I__794\ : Span4Mux_h
    port map (
            O => \N__3603\,
            I => \N__3568\
        );

    \I__793\ : Span4Mux_h
    port map (
            O => \N__3600\,
            I => \N__3568\
        );

    \I__792\ : Span4Mux_v
    port map (
            O => \N__3597\,
            I => \N__3568\
        );

    \I__791\ : Span4Mux_v
    port map (
            O => \N__3594\,
            I => \N__3568\
        );

    \I__790\ : Span4Mux_v
    port map (
            O => \N__3589\,
            I => \N__3568\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__3586\,
            I => \N__3568\
        );

    \I__788\ : Span4Mux_v
    port map (
            O => \N__3581\,
            I => \N__3565\
        );

    \I__787\ : Span4Mux_h
    port map (
            O => \N__3568\,
            I => \N__3562\
        );

    \I__786\ : Span4Mux_v
    port map (
            O => \N__3565\,
            I => \N__3559\
        );

    \I__785\ : Span4Mux_v
    port map (
            O => \N__3562\,
            I => \N__3556\
        );

    \I__784\ : Sp12to4
    port map (
            O => \N__3559\,
            I => \N__3553\
        );

    \I__783\ : Span4Mux_v
    port map (
            O => \N__3556\,
            I => \N__3550\
        );

    \I__782\ : Odrv12
    port map (
            O => \N__3553\,
            I => \ICLK\
        );

    \I__781\ : Odrv4
    port map (
            O => \N__3550\,
            I => \ICLK\
        );

    \I__780\ : CEMux
    port map (
            O => \N__3545\,
            I => \N__3542\
        );

    \I__779\ : LocalMux
    port map (
            O => \N__3542\,
            I => \N__3537\
        );

    \I__778\ : CEMux
    port map (
            O => \N__3541\,
            I => \N__3534\
        );

    \I__777\ : CEMux
    port map (
            O => \N__3540\,
            I => \N__3530\
        );

    \I__776\ : Span4Mux_h
    port map (
            O => \N__3537\,
            I => \N__3524\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__3534\,
            I => \N__3524\
        );

    \I__774\ : CEMux
    port map (
            O => \N__3533\,
            I => \N__3521\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__3530\,
            I => \N__3518\
        );

    \I__772\ : CEMux
    port map (
            O => \N__3529\,
            I => \N__3515\
        );

    \I__771\ : Span4Mux_h
    port map (
            O => \N__3524\,
            I => \N__3510\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__3521\,
            I => \N__3510\
        );

    \I__769\ : Span4Mux_h
    port map (
            O => \N__3518\,
            I => \N__3505\
        );

    \I__768\ : LocalMux
    port map (
            O => \N__3515\,
            I => \N__3505\
        );

    \I__767\ : Span4Mux_h
    port map (
            O => \N__3510\,
            I => \N__3502\
        );

    \I__766\ : Span4Mux_h
    port map (
            O => \N__3505\,
            I => \N__3499\
        );

    \I__765\ : Odrv4
    port map (
            O => \N__3502\,
            I => n307
        );

    \I__764\ : Odrv4
    port map (
            O => \N__3499\,
            I => n307
        );

    \I__763\ : InMux
    port map (
            O => \N__3494\,
            I => \N__3491\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__3491\,
            I => \N__3488\
        );

    \I__761\ : Span4Mux_h
    port map (
            O => \N__3488\,
            I => \N__3485\
        );

    \I__760\ : Odrv4
    port map (
            O => \N__3485\,
            I => n26_adj_2
        );

    \I__759\ : InMux
    port map (
            O => \N__3482\,
            I => \N__3479\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__3479\,
            I => \N__3476\
        );

    \I__757\ : Span4Mux_h
    port map (
            O => \N__3476\,
            I => \N__3473\
        );

    \I__756\ : Odrv4
    port map (
            O => \N__3473\,
            I => n27_adj_18
        );

    \I__755\ : CascadeMux
    port map (
            O => \N__3470\,
            I => \N__3467\
        );

    \I__754\ : InMux
    port map (
            O => \N__3467\,
            I => \N__3464\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__3464\,
            I => \N__3461\
        );

    \I__752\ : Odrv4
    port map (
            O => \N__3461\,
            I => n28_adj_1
        );

    \I__751\ : InMux
    port map (
            O => \N__3458\,
            I => \N__3455\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__3455\,
            I => \N__3452\
        );

    \I__749\ : Span4Mux_h
    port map (
            O => \N__3452\,
            I => \N__3449\
        );

    \I__748\ : Odrv4
    port map (
            O => \N__3449\,
            I => n447
        );

    \I__747\ : CascadeMux
    port map (
            O => \N__3446\,
            I => \n441_cascade_\
        );

    \I__746\ : CEMux
    port map (
            O => \N__3443\,
            I => \N__3440\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__3440\,
            I => \N__3437\
        );

    \I__744\ : Span4Mux_v
    port map (
            O => \N__3437\,
            I => \N__3434\
        );

    \I__743\ : Odrv4
    port map (
            O => \N__3434\,
            I => n6_adj_3
        );

    \I__742\ : InMux
    port map (
            O => \N__3431\,
            I => \N__3428\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__3428\,
            I => n441
        );

    \I__740\ : SRMux
    port map (
            O => \N__3425\,
            I => \N__3422\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__3422\,
            I => \N__3419\
        );

    \I__738\ : Span4Mux_h
    port map (
            O => \N__3419\,
            I => \N__3416\
        );

    \I__737\ : Odrv4
    port map (
            O => \N__3416\,
            I => n386
        );

    \I__736\ : CEMux
    port map (
            O => \N__3413\,
            I => \N__3408\
        );

    \I__735\ : CEMux
    port map (
            O => \N__3412\,
            I => \N__3403\
        );

    \I__734\ : CEMux
    port map (
            O => \N__3411\,
            I => \N__3399\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__3408\,
            I => \N__3395\
        );

    \I__732\ : CEMux
    port map (
            O => \N__3407\,
            I => \N__3392\
        );

    \I__731\ : CEMux
    port map (
            O => \N__3406\,
            I => \N__3389\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__3403\,
            I => \N__3386\
        );

    \I__729\ : InMux
    port map (
            O => \N__3402\,
            I => \N__3383\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__3399\,
            I => \N__3380\
        );

    \I__727\ : CEMux
    port map (
            O => \N__3398\,
            I => \N__3377\
        );

    \I__726\ : Span4Mux_v
    port map (
            O => \N__3395\,
            I => \N__3372\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__3392\,
            I => \N__3372\
        );

    \I__724\ : LocalMux
    port map (
            O => \N__3389\,
            I => \N__3369\
        );

    \I__723\ : Span4Mux_v
    port map (
            O => \N__3386\,
            I => \N__3364\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__3383\,
            I => \N__3364\
        );

    \I__721\ : Span4Mux_v
    port map (
            O => \N__3380\,
            I => \N__3359\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__3377\,
            I => \N__3359\
        );

    \I__719\ : Span4Mux_h
    port map (
            O => \N__3372\,
            I => \N__3356\
        );

    \I__718\ : Span4Mux_h
    port map (
            O => \N__3369\,
            I => \N__3351\
        );

    \I__717\ : Span4Mux_h
    port map (
            O => \N__3364\,
            I => \N__3351\
        );

    \I__716\ : Odrv4
    port map (
            O => \N__3359\,
            I => \div_state_1__N_88\
        );

    \I__715\ : Odrv4
    port map (
            O => \N__3356\,
            I => \div_state_1__N_88\
        );

    \I__714\ : Odrv4
    port map (
            O => \N__3351\,
            I => \div_state_1__N_88\
        );

    \I__713\ : InMux
    port map (
            O => \N__3344\,
            I => \N__3330\
        );

    \I__712\ : InMux
    port map (
            O => \N__3343\,
            I => \N__3325\
        );

    \I__711\ : InMux
    port map (
            O => \N__3342\,
            I => \N__3325\
        );

    \I__710\ : InMux
    port map (
            O => \N__3341\,
            I => \N__3313\
        );

    \I__709\ : InMux
    port map (
            O => \N__3340\,
            I => \N__3313\
        );

    \I__708\ : InMux
    port map (
            O => \N__3339\,
            I => \N__3313\
        );

    \I__707\ : InMux
    port map (
            O => \N__3338\,
            I => \N__3313\
        );

    \I__706\ : InMux
    port map (
            O => \N__3337\,
            I => \N__3313\
        );

    \I__705\ : InMux
    port map (
            O => \N__3336\,
            I => \N__3304\
        );

    \I__704\ : InMux
    port map (
            O => \N__3335\,
            I => \N__3304\
        );

    \I__703\ : InMux
    port map (
            O => \N__3334\,
            I => \N__3304\
        );

    \I__702\ : InMux
    port map (
            O => \N__3333\,
            I => \N__3304\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__3330\,
            I => \N__3299\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__3325\,
            I => \N__3299\
        );

    \I__699\ : CascadeMux
    port map (
            O => \N__3324\,
            I => \N__3294\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__3313\,
            I => \N__3288\
        );

    \I__697\ : LocalMux
    port map (
            O => \N__3304\,
            I => \N__3288\
        );

    \I__696\ : Span4Mux_v
    port map (
            O => \N__3299\,
            I => \N__3285\
        );

    \I__695\ : InMux
    port map (
            O => \N__3298\,
            I => \N__3278\
        );

    \I__694\ : InMux
    port map (
            O => \N__3297\,
            I => \N__3278\
        );

    \I__693\ : InMux
    port map (
            O => \N__3294\,
            I => \N__3278\
        );

    \I__692\ : CascadeMux
    port map (
            O => \N__3293\,
            I => \N__3273\
        );

    \I__691\ : Span4Mux_h
    port map (
            O => \N__3288\,
            I => \N__3268\
        );

    \I__690\ : Sp12to4
    port map (
            O => \N__3285\,
            I => \N__3263\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__3278\,
            I => \N__3263\
        );

    \I__688\ : InMux
    port map (
            O => \N__3277\,
            I => \N__3260\
        );

    \I__687\ : InMux
    port map (
            O => \N__3276\,
            I => \N__3257\
        );

    \I__686\ : InMux
    port map (
            O => \N__3273\,
            I => \N__3250\
        );

    \I__685\ : InMux
    port map (
            O => \N__3272\,
            I => \N__3250\
        );

    \I__684\ : InMux
    port map (
            O => \N__3271\,
            I => \N__3250\
        );

    \I__683\ : Odrv4
    port map (
            O => \N__3268\,
            I => div_state_0
        );

    \I__682\ : Odrv12
    port map (
            O => \N__3263\,
            I => div_state_0
        );

    \I__681\ : LocalMux
    port map (
            O => \N__3260\,
            I => div_state_0
        );

    \I__680\ : LocalMux
    port map (
            O => \N__3257\,
            I => div_state_0
        );

    \I__679\ : LocalMux
    port map (
            O => \N__3250\,
            I => div_state_0
        );

    \I__678\ : InMux
    port map (
            O => \N__3239\,
            I => \N__3236\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__3236\,
            I => \N__3232\
        );

    \I__676\ : InMux
    port map (
            O => \N__3235\,
            I => \N__3229\
        );

    \I__675\ : Span4Mux_v
    port map (
            O => \N__3232\,
            I => \N__3226\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__3229\,
            I => t0off_12
        );

    \I__673\ : Odrv4
    port map (
            O => \N__3226\,
            I => t0off_12
        );

    \I__672\ : InMux
    port map (
            O => \N__3221\,
            I => \N__3217\
        );

    \I__671\ : InMux
    port map (
            O => \N__3220\,
            I => \N__3214\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__3217\,
            I => \N__3211\
        );

    \I__669\ : LocalMux
    port map (
            O => \N__3214\,
            I => t0off_2
        );

    \I__668\ : Odrv4
    port map (
            O => \N__3211\,
            I => t0off_2
        );

    \I__667\ : CascadeMux
    port map (
            O => \N__3206\,
            I => \N__3203\
        );

    \I__666\ : InMux
    port map (
            O => \N__3203\,
            I => \N__3199\
        );

    \I__665\ : InMux
    port map (
            O => \N__3202\,
            I => \N__3196\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__3199\,
            I => \N__3193\
        );

    \I__663\ : LocalMux
    port map (
            O => \N__3196\,
            I => t0off_7
        );

    \I__662\ : Odrv4
    port map (
            O => \N__3193\,
            I => t0off_7
        );

    \I__661\ : InMux
    port map (
            O => \N__3188\,
            I => \N__3184\
        );

    \I__660\ : InMux
    port map (
            O => \N__3187\,
            I => \N__3181\
        );

    \I__659\ : LocalMux
    port map (
            O => \N__3184\,
            I => \N__3178\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__3181\,
            I => t0off_10
        );

    \I__657\ : Odrv4
    port map (
            O => \N__3178\,
            I => t0off_10
        );

    \I__656\ : CascadeMux
    port map (
            O => \N__3173\,
            I => \n27_cascade_\
        );

    \I__655\ : InMux
    port map (
            O => \N__3170\,
            I => \N__3164\
        );

    \I__654\ : InMux
    port map (
            O => \N__3169\,
            I => \N__3164\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__3164\,
            I => n442
        );

    \I__652\ : InMux
    port map (
            O => \N__3161\,
            I => \N__3158\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__3158\,
            I => \N__3155\
        );

    \I__650\ : Span4Mux_h
    port map (
            O => \N__3155\,
            I => \N__3152\
        );

    \I__649\ : Odrv4
    port map (
            O => \N__3152\,
            I => \t0off_15_N_67_13\
        );

    \I__648\ : InMux
    port map (
            O => \N__3149\,
            I => \N__3146\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__3146\,
            I => \t0off_15_N_51_13\
        );

    \I__646\ : InMux
    port map (
            O => \N__3143\,
            I => \N__3140\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__3140\,
            I => \N__3137\
        );

    \I__644\ : Odrv4
    port map (
            O => \N__3137\,
            I => \t0off_15_N_67_7\
        );

    \I__643\ : InMux
    port map (
            O => \N__3134\,
            I => \N__3131\
        );

    \I__642\ : LocalMux
    port map (
            O => \N__3131\,
            I => \t0off_15_N_51_7\
        );

    \I__641\ : InMux
    port map (
            O => \N__3128\,
            I => \N__3125\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__3125\,
            I => \N__3122\
        );

    \I__639\ : Odrv12
    port map (
            O => \N__3122\,
            I => \t0off_15_N_67_12\
        );

    \I__638\ : InMux
    port map (
            O => \N__3119\,
            I => \N__3116\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__3116\,
            I => \t0off_15_N_51_12\
        );

    \I__636\ : InMux
    port map (
            O => \N__3113\,
            I => \N__3110\
        );

    \I__635\ : LocalMux
    port map (
            O => \N__3110\,
            I => \t0off_15_N_51_9\
        );

    \I__634\ : InMux
    port map (
            O => \N__3107\,
            I => \N__3104\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__3104\,
            I => \N__3101\
        );

    \I__632\ : Odrv4
    port map (
            O => \N__3101\,
            I => \t0off_15_N_67_9\
        );

    \I__631\ : InMux
    port map (
            O => \N__3098\,
            I => \N__3095\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__3095\,
            I => \N__3092\
        );

    \I__629\ : Odrv12
    port map (
            O => \N__3092\,
            I => \t0off_15_N_67_14\
        );

    \I__628\ : InMux
    port map (
            O => \N__3089\,
            I => \N__3086\
        );

    \I__627\ : LocalMux
    port map (
            O => \N__3086\,
            I => \t0off_15_N_51_14\
        );

    \I__626\ : InMux
    port map (
            O => \N__3083\,
            I => \N__3080\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__3080\,
            I => \N__3077\
        );

    \I__624\ : Span4Mux_v
    port map (
            O => \N__3077\,
            I => \N__3074\
        );

    \I__623\ : Odrv4
    port map (
            O => \N__3074\,
            I => \t0off_15_N_67_4\
        );

    \I__622\ : InMux
    port map (
            O => \N__3071\,
            I => \N__3068\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__3068\,
            I => \t0off_15_N_51_4\
        );

    \I__620\ : InMux
    port map (
            O => \N__3065\,
            I => \N__3062\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__3062\,
            I => \N__3059\
        );

    \I__618\ : Span4Mux_v
    port map (
            O => \N__3059\,
            I => \N__3056\
        );

    \I__617\ : Odrv4
    port map (
            O => \N__3056\,
            I => \t0off_15_N_67_1\
        );

    \I__616\ : InMux
    port map (
            O => \N__3053\,
            I => \N__3050\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__3050\,
            I => \t0off_15_N_51_1\
        );

    \I__614\ : InMux
    port map (
            O => \N__3047\,
            I => \N__3044\
        );

    \I__613\ : LocalMux
    port map (
            O => \N__3044\,
            I => \N__3041\
        );

    \I__612\ : Span4Mux_h
    port map (
            O => \N__3041\,
            I => \N__3038\
        );

    \I__611\ : Odrv4
    port map (
            O => \N__3038\,
            I => \t0off_15_N_67_0\
        );

    \I__610\ : InMux
    port map (
            O => \N__3035\,
            I => \N__3032\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__3032\,
            I => \t0off_15_N_51_0\
        );

    \I__608\ : InMux
    port map (
            O => \N__3029\,
            I => \N__3026\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__3026\,
            I => \t0on_15_N_35_9\
        );

    \I__606\ : CascadeMux
    port map (
            O => \N__3023\,
            I => \N__3020\
        );

    \I__605\ : InMux
    port map (
            O => \N__3020\,
            I => \N__3016\
        );

    \I__604\ : InMux
    port map (
            O => \N__3019\,
            I => \N__3013\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__3016\,
            I => t0on_9
        );

    \I__602\ : LocalMux
    port map (
            O => \N__3013\,
            I => t0on_9
        );

    \I__601\ : InMux
    port map (
            O => \N__3008\,
            I => \N__3004\
        );

    \I__600\ : InMux
    port map (
            O => \N__3007\,
            I => \N__3001\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__3004\,
            I => \N__2998\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__3001\,
            I => \N__2995\
        );

    \I__597\ : Span4Mux_v
    port map (
            O => \N__2998\,
            I => \N__2991\
        );

    \I__596\ : Span4Mux_v
    port map (
            O => \N__2995\,
            I => \N__2988\
        );

    \I__595\ : InMux
    port map (
            O => \N__2994\,
            I => \N__2985\
        );

    \I__594\ : Sp12to4
    port map (
            O => \N__2991\,
            I => \N__2978\
        );

    \I__593\ : Sp12to4
    port map (
            O => \N__2988\,
            I => \N__2978\
        );

    \I__592\ : LocalMux
    port map (
            O => \N__2985\,
            I => \N__2978\
        );

    \I__591\ : Odrv12
    port map (
            O => \N__2978\,
            I => \DIVIDE_15_\
        );

    \I__590\ : InMux
    port map (
            O => \N__2975\,
            I => \N__2972\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__2972\,
            I => \t0on_15_N_35_14\
        );

    \I__588\ : InMux
    port map (
            O => \N__2969\,
            I => \N__2965\
        );

    \I__587\ : InMux
    port map (
            O => \N__2968\,
            I => \N__2962\
        );

    \I__586\ : LocalMux
    port map (
            O => \N__2965\,
            I => t0on_14
        );

    \I__585\ : LocalMux
    port map (
            O => \N__2962\,
            I => t0on_14
        );

    \I__584\ : InMux
    port map (
            O => \N__2957\,
            I => \N__2953\
        );

    \I__583\ : InMux
    port map (
            O => \N__2956\,
            I => \N__2950\
        );

    \I__582\ : LocalMux
    port map (
            O => \N__2953\,
            I => \N__2945\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__2950\,
            I => \N__2945\
        );

    \I__580\ : Span4Mux_v
    port map (
            O => \N__2945\,
            I => \N__2941\
        );

    \I__579\ : InMux
    port map (
            O => \N__2944\,
            I => \N__2938\
        );

    \I__578\ : Sp12to4
    port map (
            O => \N__2941\,
            I => \N__2933\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__2938\,
            I => \N__2933\
        );

    \I__576\ : Odrv12
    port map (
            O => \N__2933\,
            I => \DIVIDE_12_\
        );

    \I__575\ : InMux
    port map (
            O => \N__2930\,
            I => \N__2927\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__2927\,
            I => \N__2924\
        );

    \I__573\ : Span4Mux_v
    port map (
            O => \N__2924\,
            I => \N__2921\
        );

    \I__572\ : Odrv4
    port map (
            O => \N__2921\,
            I => n6
        );

    \I__571\ : InMux
    port map (
            O => \N__2918\,
            I => \N__2912\
        );

    \I__570\ : InMux
    port map (
            O => \N__2917\,
            I => \N__2912\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__2912\,
            I => \N__2909\
        );

    \I__568\ : Span4Mux_v
    port map (
            O => \N__2909\,
            I => \N__2905\
        );

    \I__567\ : InMux
    port map (
            O => \N__2908\,
            I => \N__2902\
        );

    \I__566\ : Sp12to4
    port map (
            O => \N__2905\,
            I => \N__2897\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__2902\,
            I => \N__2897\
        );

    \I__564\ : Odrv12
    port map (
            O => \N__2897\,
            I => \DIVIDE_10_\
        );

    \I__563\ : CascadeMux
    port map (
            O => \N__2894\,
            I => \N__2891\
        );

    \I__562\ : InMux
    port map (
            O => \N__2891\,
            I => \N__2888\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__2888\,
            I => \N__2885\
        );

    \I__560\ : Span4Mux_v
    port map (
            O => \N__2885\,
            I => \N__2882\
        );

    \I__559\ : Odrv4
    port map (
            O => \N__2882\,
            I => n8
        );

    \I__558\ : InMux
    port map (
            O => \N__2879\,
            I => \N__2876\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__2876\,
            I => \N__2873\
        );

    \I__556\ : Odrv12
    port map (
            O => \N__2873\,
            I => \t0off_15_N_67_3\
        );

    \I__555\ : InMux
    port map (
            O => \N__2870\,
            I => \N__2867\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__2867\,
            I => \t0off_15_N_51_3\
        );

    \I__553\ : InMux
    port map (
            O => \N__2864\,
            I => \N__2861\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__2861\,
            I => \N__2858\
        );

    \I__551\ : Span4Mux_v
    port map (
            O => \N__2858\,
            I => \N__2855\
        );

    \I__550\ : Odrv4
    port map (
            O => \N__2855\,
            I => \t0off_15_N_67_8\
        );

    \I__549\ : InMux
    port map (
            O => \N__2852\,
            I => \N__2849\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__2849\,
            I => \t0off_15_N_51_8\
        );

    \I__547\ : InMux
    port map (
            O => \N__2846\,
            I => \N__2843\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__2843\,
            I => \N__2840\
        );

    \I__545\ : Odrv4
    port map (
            O => \N__2840\,
            I => \t0off_15_N_67_2\
        );

    \I__544\ : InMux
    port map (
            O => \N__2837\,
            I => \N__2834\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__2834\,
            I => \t0off_15_N_51_2\
        );

    \I__542\ : CascadeMux
    port map (
            O => \N__2831\,
            I => \N__2828\
        );

    \I__541\ : InMux
    port map (
            O => \N__2828\,
            I => \N__2825\
        );

    \I__540\ : LocalMux
    port map (
            O => \N__2825\,
            I => \N__2822\
        );

    \I__539\ : Span4Mux_v
    port map (
            O => \N__2822\,
            I => \N__2819\
        );

    \I__538\ : Odrv4
    port map (
            O => \N__2819\,
            I => \t0off_15_N_67_10\
        );

    \I__537\ : InMux
    port map (
            O => \N__2816\,
            I => \N__2813\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__2813\,
            I => \t0off_15_N_51_10\
        );

    \I__535\ : CascadeMux
    port map (
            O => \N__2810\,
            I => \N__2801\
        );

    \I__534\ : CascadeMux
    port map (
            O => \N__2809\,
            I => \N__2798\
        );

    \I__533\ : CascadeMux
    port map (
            O => \N__2808\,
            I => \N__2795\
        );

    \I__532\ : CascadeMux
    port map (
            O => \N__2807\,
            I => \N__2791\
        );

    \I__531\ : CascadeMux
    port map (
            O => \N__2806\,
            I => \N__2788\
        );

    \I__530\ : CascadeMux
    port map (
            O => \N__2805\,
            I => \N__2785\
        );

    \I__529\ : InMux
    port map (
            O => \N__2804\,
            I => \N__2761\
        );

    \I__528\ : InMux
    port map (
            O => \N__2801\,
            I => \N__2761\
        );

    \I__527\ : InMux
    port map (
            O => \N__2798\,
            I => \N__2761\
        );

    \I__526\ : InMux
    port map (
            O => \N__2795\,
            I => \N__2750\
        );

    \I__525\ : InMux
    port map (
            O => \N__2794\,
            I => \N__2750\
        );

    \I__524\ : InMux
    port map (
            O => \N__2791\,
            I => \N__2750\
        );

    \I__523\ : InMux
    port map (
            O => \N__2788\,
            I => \N__2750\
        );

    \I__522\ : InMux
    port map (
            O => \N__2785\,
            I => \N__2750\
        );

    \I__521\ : CascadeMux
    port map (
            O => \N__2784\,
            I => \N__2747\
        );

    \I__520\ : CascadeMux
    port map (
            O => \N__2783\,
            I => \N__2744\
        );

    \I__519\ : CascadeMux
    port map (
            O => \N__2782\,
            I => \N__2741\
        );

    \I__518\ : CascadeMux
    port map (
            O => \N__2781\,
            I => \N__2738\
        );

    \I__517\ : CascadeMux
    port map (
            O => \N__2780\,
            I => \N__2735\
        );

    \I__516\ : CascadeMux
    port map (
            O => \N__2779\,
            I => \N__2732\
        );

    \I__515\ : CascadeMux
    port map (
            O => \N__2778\,
            I => \N__2729\
        );

    \I__514\ : CascadeMux
    port map (
            O => \N__2777\,
            I => \N__2725\
        );

    \I__513\ : CascadeMux
    port map (
            O => \N__2776\,
            I => \N__2721\
        );

    \I__512\ : CascadeMux
    port map (
            O => \N__2775\,
            I => \N__2717\
        );

    \I__511\ : CascadeMux
    port map (
            O => \N__2774\,
            I => \N__2713\
        );

    \I__510\ : CascadeMux
    port map (
            O => \N__2773\,
            I => \N__2710\
        );

    \I__509\ : CascadeMux
    port map (
            O => \N__2772\,
            I => \N__2706\
        );

    \I__508\ : CascadeMux
    port map (
            O => \N__2771\,
            I => \N__2703\
        );

    \I__507\ : CascadeMux
    port map (
            O => \N__2770\,
            I => \N__2700\
        );

    \I__506\ : CascadeMux
    port map (
            O => \N__2769\,
            I => \N__2697\
        );

    \I__505\ : CascadeMux
    port map (
            O => \N__2768\,
            I => \N__2694\
        );

    \I__504\ : LocalMux
    port map (
            O => \N__2761\,
            I => \N__2689\
        );

    \I__503\ : LocalMux
    port map (
            O => \N__2750\,
            I => \N__2689\
        );

    \I__502\ : InMux
    port map (
            O => \N__2747\,
            I => \N__2682\
        );

    \I__501\ : InMux
    port map (
            O => \N__2744\,
            I => \N__2682\
        );

    \I__500\ : InMux
    port map (
            O => \N__2741\,
            I => \N__2682\
        );

    \I__499\ : InMux
    port map (
            O => \N__2738\,
            I => \N__2673\
        );

    \I__498\ : InMux
    port map (
            O => \N__2735\,
            I => \N__2673\
        );

    \I__497\ : InMux
    port map (
            O => \N__2732\,
            I => \N__2673\
        );

    \I__496\ : InMux
    port map (
            O => \N__2729\,
            I => \N__2673\
        );

    \I__495\ : InMux
    port map (
            O => \N__2728\,
            I => \N__2656\
        );

    \I__494\ : InMux
    port map (
            O => \N__2725\,
            I => \N__2656\
        );

    \I__493\ : InMux
    port map (
            O => \N__2724\,
            I => \N__2656\
        );

    \I__492\ : InMux
    port map (
            O => \N__2721\,
            I => \N__2656\
        );

    \I__491\ : InMux
    port map (
            O => \N__2720\,
            I => \N__2656\
        );

    \I__490\ : InMux
    port map (
            O => \N__2717\,
            I => \N__2656\
        );

    \I__489\ : InMux
    port map (
            O => \N__2716\,
            I => \N__2656\
        );

    \I__488\ : InMux
    port map (
            O => \N__2713\,
            I => \N__2656\
        );

    \I__487\ : InMux
    port map (
            O => \N__2710\,
            I => \N__2647\
        );

    \I__486\ : InMux
    port map (
            O => \N__2709\,
            I => \N__2647\
        );

    \I__485\ : InMux
    port map (
            O => \N__2706\,
            I => \N__2647\
        );

    \I__484\ : InMux
    port map (
            O => \N__2703\,
            I => \N__2647\
        );

    \I__483\ : InMux
    port map (
            O => \N__2700\,
            I => \N__2640\
        );

    \I__482\ : InMux
    port map (
            O => \N__2697\,
            I => \N__2640\
        );

    \I__481\ : InMux
    port map (
            O => \N__2694\,
            I => \N__2640\
        );

    \I__480\ : Span4Mux_v
    port map (
            O => \N__2689\,
            I => \N__2627\
        );

    \I__479\ : LocalMux
    port map (
            O => \N__2682\,
            I => \N__2627\
        );

    \I__478\ : LocalMux
    port map (
            O => \N__2673\,
            I => \N__2627\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__2656\,
            I => \N__2627\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__2647\,
            I => \N__2627\
        );

    \I__475\ : LocalMux
    port map (
            O => \N__2640\,
            I => \N__2627\
        );

    \I__474\ : Span4Mux_v
    port map (
            O => \N__2627\,
            I => \N__2624\
        );

    \I__473\ : Odrv4
    port map (
            O => \N__2624\,
            I => \CONSTANT_ONE_NET\
        );

    \I__472\ : InMux
    port map (
            O => \N__2621\,
            I => n402
        );

    \I__471\ : CascadeMux
    port map (
            O => \N__2618\,
            I => \N__2615\
        );

    \I__470\ : InMux
    port map (
            O => \N__2615\,
            I => \N__2612\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__2612\,
            I => \t0off_15_N_51_15\
        );

    \I__468\ : CascadeMux
    port map (
            O => \N__2609\,
            I => \N__2604\
        );

    \I__467\ : InMux
    port map (
            O => \N__2608\,
            I => \N__2601\
        );

    \I__466\ : InMux
    port map (
            O => \N__2607\,
            I => \N__2598\
        );

    \I__465\ : InMux
    port map (
            O => \N__2604\,
            I => \N__2595\
        );

    \I__464\ : LocalMux
    port map (
            O => \N__2601\,
            I => \N__2592\
        );

    \I__463\ : LocalMux
    port map (
            O => \N__2598\,
            I => \N__2587\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__2595\,
            I => \N__2587\
        );

    \I__461\ : Span4Mux_v
    port map (
            O => \N__2592\,
            I => \N__2584\
        );

    \I__460\ : Sp12to4
    port map (
            O => \N__2587\,
            I => \N__2581\
        );

    \I__459\ : Span4Mux_h
    port map (
            O => \N__2584\,
            I => \N__2578\
        );

    \I__458\ : Span12Mux_v
    port map (
            O => \N__2581\,
            I => \N__2575\
        );

    \I__457\ : Span4Mux_v
    port map (
            O => \N__2578\,
            I => \N__2572\
        );

    \I__456\ : Odrv12
    port map (
            O => \N__2575\,
            I => \DIVIDE_11_\
        );

    \I__455\ : Odrv4
    port map (
            O => \N__2572\,
            I => \DIVIDE_11_\
        );

    \I__454\ : InMux
    port map (
            O => \N__2567\,
            I => \N__2564\
        );

    \I__453\ : LocalMux
    port map (
            O => \N__2564\,
            I => \t0on_15_N_35_10\
        );

    \I__452\ : InMux
    port map (
            O => \N__2561\,
            I => \N__2557\
        );

    \I__451\ : InMux
    port map (
            O => \N__2560\,
            I => \N__2554\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__2557\,
            I => t0on_10
        );

    \I__449\ : LocalMux
    port map (
            O => \N__2554\,
            I => t0on_10
        );

    \I__448\ : CascadeMux
    port map (
            O => \N__2549\,
            I => \N__2545\
        );

    \I__447\ : InMux
    port map (
            O => \N__2548\,
            I => \N__2541\
        );

    \I__446\ : InMux
    port map (
            O => \N__2545\,
            I => \N__2538\
        );

    \I__445\ : InMux
    port map (
            O => \N__2544\,
            I => \N__2535\
        );

    \I__444\ : LocalMux
    port map (
            O => \N__2541\,
            I => \N__2532\
        );

    \I__443\ : LocalMux
    port map (
            O => \N__2538\,
            I => \N__2527\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__2535\,
            I => \N__2527\
        );

    \I__441\ : Sp12to4
    port map (
            O => \N__2532\,
            I => \N__2524\
        );

    \I__440\ : Span4Mux_v
    port map (
            O => \N__2527\,
            I => \N__2521\
        );

    \I__439\ : Span12Mux_v
    port map (
            O => \N__2524\,
            I => \N__2516\
        );

    \I__438\ : Sp12to4
    port map (
            O => \N__2521\,
            I => \N__2516\
        );

    \I__437\ : Odrv12
    port map (
            O => \N__2516\,
            I => \DIVIDE_3_\
        );

    \I__436\ : InMux
    port map (
            O => \N__2513\,
            I => \N__2510\
        );

    \I__435\ : LocalMux
    port map (
            O => \N__2510\,
            I => \t0on_15_N_35_2\
        );

    \I__434\ : InMux
    port map (
            O => \N__2507\,
            I => \N__2503\
        );

    \I__433\ : InMux
    port map (
            O => \N__2506\,
            I => \N__2500\
        );

    \I__432\ : LocalMux
    port map (
            O => \N__2503\,
            I => t0on_2
        );

    \I__431\ : LocalMux
    port map (
            O => \N__2500\,
            I => t0on_2
        );

    \I__430\ : InMux
    port map (
            O => \N__2495\,
            I => \N__2492\
        );

    \I__429\ : LocalMux
    port map (
            O => \N__2492\,
            I => \N__2487\
        );

    \I__428\ : InMux
    port map (
            O => \N__2491\,
            I => \N__2484\
        );

    \I__427\ : InMux
    port map (
            O => \N__2490\,
            I => \N__2481\
        );

    \I__426\ : Span4Mux_v
    port map (
            O => \N__2487\,
            I => \N__2476\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__2484\,
            I => \N__2476\
        );

    \I__424\ : LocalMux
    port map (
            O => \N__2481\,
            I => \N__2473\
        );

    \I__423\ : Span4Mux_v
    port map (
            O => \N__2476\,
            I => \N__2470\
        );

    \I__422\ : Sp12to4
    port map (
            O => \N__2473\,
            I => \N__2467\
        );

    \I__421\ : Span4Mux_h
    port map (
            O => \N__2470\,
            I => \N__2464\
        );

    \I__420\ : Span12Mux_v
    port map (
            O => \N__2467\,
            I => \N__2461\
        );

    \I__419\ : Span4Mux_v
    port map (
            O => \N__2464\,
            I => \N__2458\
        );

    \I__418\ : Odrv12
    port map (
            O => \N__2461\,
            I => \DIVIDE_13_\
        );

    \I__417\ : Odrv4
    port map (
            O => \N__2458\,
            I => \DIVIDE_13_\
        );

    \I__416\ : InMux
    port map (
            O => \N__2453\,
            I => \N__2450\
        );

    \I__415\ : LocalMux
    port map (
            O => \N__2450\,
            I => \t0on_15_N_35_12\
        );

    \I__414\ : InMux
    port map (
            O => \N__2447\,
            I => \N__2443\
        );

    \I__413\ : InMux
    port map (
            O => \N__2446\,
            I => \N__2440\
        );

    \I__412\ : LocalMux
    port map (
            O => \N__2443\,
            I => t0on_12
        );

    \I__411\ : LocalMux
    port map (
            O => \N__2440\,
            I => t0on_12
        );

    \I__410\ : InMux
    port map (
            O => \N__2435\,
            I => \N__2430\
        );

    \I__409\ : InMux
    port map (
            O => \N__2434\,
            I => \N__2427\
        );

    \I__408\ : InMux
    port map (
            O => \N__2433\,
            I => \N__2424\
        );

    \I__407\ : LocalMux
    port map (
            O => \N__2430\,
            I => \N__2421\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__2427\,
            I => \N__2416\
        );

    \I__405\ : LocalMux
    port map (
            O => \N__2424\,
            I => \N__2416\
        );

    \I__404\ : Span4Mux_v
    port map (
            O => \N__2421\,
            I => \N__2413\
        );

    \I__403\ : Span4Mux_v
    port map (
            O => \N__2416\,
            I => \N__2410\
        );

    \I__402\ : Sp12to4
    port map (
            O => \N__2413\,
            I => \N__2407\
        );

    \I__401\ : Span4Mux_v
    port map (
            O => \N__2410\,
            I => \N__2404\
        );

    \I__400\ : Span12Mux_v
    port map (
            O => \N__2407\,
            I => \N__2401\
        );

    \I__399\ : Span4Mux_h
    port map (
            O => \N__2404\,
            I => \N__2398\
        );

    \I__398\ : Odrv12
    port map (
            O => \N__2401\,
            I => \DIVIDE_8_\
        );

    \I__397\ : Odrv4
    port map (
            O => \N__2398\,
            I => \DIVIDE_8_\
        );

    \I__396\ : InMux
    port map (
            O => \N__2393\,
            I => \N__2390\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__2390\,
            I => \t0on_15_N_35_7\
        );

    \I__394\ : CascadeMux
    port map (
            O => \N__2387\,
            I => \N__2383\
        );

    \I__393\ : InMux
    port map (
            O => \N__2386\,
            I => \N__2380\
        );

    \I__392\ : InMux
    port map (
            O => \N__2383\,
            I => \N__2377\
        );

    \I__391\ : LocalMux
    port map (
            O => \N__2380\,
            I => t0on_7
        );

    \I__390\ : LocalMux
    port map (
            O => \N__2377\,
            I => t0on_7
        );

    \I__389\ : CascadeMux
    port map (
            O => \N__2372\,
            I => \N__2368\
        );

    \I__388\ : InMux
    port map (
            O => \N__2371\,
            I => \N__2365\
        );

    \I__387\ : InMux
    port map (
            O => \N__2368\,
            I => \N__2362\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__2365\,
            I => t0on_15
        );

    \I__385\ : LocalMux
    port map (
            O => \N__2362\,
            I => t0on_15
        );

    \I__384\ : InMux
    port map (
            O => \N__2357\,
            I => \N__2354\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__2354\,
            I => \t0on_15_N_35_11\
        );

    \I__382\ : CascadeMux
    port map (
            O => \N__2351\,
            I => \N__2348\
        );

    \I__381\ : InMux
    port map (
            O => \N__2348\,
            I => \N__2345\
        );

    \I__380\ : LocalMux
    port map (
            O => \N__2345\,
            I => \N__2341\
        );

    \I__379\ : InMux
    port map (
            O => \N__2344\,
            I => \N__2338\
        );

    \I__378\ : Odrv4
    port map (
            O => \N__2341\,
            I => t0on_11
        );

    \I__377\ : LocalMux
    port map (
            O => \N__2338\,
            I => t0on_11
        );

    \I__376\ : InMux
    port map (
            O => \N__2333\,
            I => n392
        );

    \I__375\ : InMux
    port map (
            O => \N__2330\,
            I => n393
        );

    \I__374\ : InMux
    port map (
            O => \N__2327\,
            I => n394
        );

    \I__373\ : InMux
    port map (
            O => \N__2324\,
            I => \bfn_2_10_0_\
        );

    \I__372\ : InMux
    port map (
            O => \N__2321\,
            I => n396
        );

    \I__371\ : InMux
    port map (
            O => \N__2318\,
            I => n397
        );

    \I__370\ : InMux
    port map (
            O => \N__2315\,
            I => n398
        );

    \I__369\ : InMux
    port map (
            O => \N__2312\,
            I => n399
        );

    \I__368\ : InMux
    port map (
            O => \N__2309\,
            I => n400
        );

    \I__367\ : InMux
    port map (
            O => \N__2306\,
            I => n401
        );

    \I__366\ : InMux
    port map (
            O => \N__2303\,
            I => n414
        );

    \I__365\ : CascadeMux
    port map (
            O => \N__2300\,
            I => \N__2297\
        );

    \I__364\ : InMux
    port map (
            O => \N__2297\,
            I => \N__2293\
        );

    \I__363\ : InMux
    port map (
            O => \N__2296\,
            I => \N__2290\
        );

    \I__362\ : LocalMux
    port map (
            O => \N__2293\,
            I => t0on_13
        );

    \I__361\ : LocalMux
    port map (
            O => \N__2290\,
            I => t0on_13
        );

    \I__360\ : InMux
    port map (
            O => \N__2285\,
            I => \N__2282\
        );

    \I__359\ : LocalMux
    port map (
            O => \N__2282\,
            I => \t0on_15_N_35_13\
        );

    \I__358\ : InMux
    port map (
            O => \N__2279\,
            I => n415
        );

    \I__357\ : InMux
    port map (
            O => \N__2276\,
            I => n416
        );

    \I__356\ : InMux
    port map (
            O => \N__2273\,
            I => n417
        );

    \I__355\ : InMux
    port map (
            O => \N__2270\,
            I => \bfn_2_9_0_\
        );

    \I__354\ : InMux
    port map (
            O => \N__2267\,
            I => n388
        );

    \I__353\ : InMux
    port map (
            O => \N__2264\,
            I => n389
        );

    \I__352\ : InMux
    port map (
            O => \N__2261\,
            I => n390
        );

    \I__351\ : InMux
    port map (
            O => \N__2258\,
            I => n391
        );

    \I__350\ : CascadeMux
    port map (
            O => \N__2255\,
            I => \N__2251\
        );

    \I__349\ : InMux
    port map (
            O => \N__2254\,
            I => \N__2248\
        );

    \I__348\ : InMux
    port map (
            O => \N__2251\,
            I => \N__2245\
        );

    \I__347\ : LocalMux
    port map (
            O => \N__2248\,
            I => t0on_4
        );

    \I__346\ : LocalMux
    port map (
            O => \N__2245\,
            I => t0on_4
        );

    \I__345\ : InMux
    port map (
            O => \N__2240\,
            I => \N__2237\
        );

    \I__344\ : LocalMux
    port map (
            O => \N__2237\,
            I => \t0on_15_N_35_4\
        );

    \I__343\ : InMux
    port map (
            O => \N__2234\,
            I => n406
        );

    \I__342\ : CascadeMux
    port map (
            O => \N__2231\,
            I => \N__2227\
        );

    \I__341\ : CascadeMux
    port map (
            O => \N__2230\,
            I => \N__2224\
        );

    \I__340\ : InMux
    port map (
            O => \N__2227\,
            I => \N__2221\
        );

    \I__339\ : InMux
    port map (
            O => \N__2224\,
            I => \N__2218\
        );

    \I__338\ : LocalMux
    port map (
            O => \N__2221\,
            I => t0on_5
        );

    \I__337\ : LocalMux
    port map (
            O => \N__2218\,
            I => t0on_5
        );

    \I__336\ : InMux
    port map (
            O => \N__2213\,
            I => \N__2210\
        );

    \I__335\ : LocalMux
    port map (
            O => \N__2210\,
            I => \t0on_15_N_35_5\
        );

    \I__334\ : InMux
    port map (
            O => \N__2207\,
            I => n407
        );

    \I__333\ : InMux
    port map (
            O => \N__2204\,
            I => \N__2200\
        );

    \I__332\ : InMux
    port map (
            O => \N__2203\,
            I => \N__2197\
        );

    \I__331\ : LocalMux
    port map (
            O => \N__2200\,
            I => t0on_6
        );

    \I__330\ : LocalMux
    port map (
            O => \N__2197\,
            I => t0on_6
        );

    \I__329\ : InMux
    port map (
            O => \N__2192\,
            I => \N__2189\
        );

    \I__328\ : LocalMux
    port map (
            O => \N__2189\,
            I => \t0on_15_N_35_6\
        );

    \I__327\ : InMux
    port map (
            O => \N__2186\,
            I => n408
        );

    \I__326\ : InMux
    port map (
            O => \N__2183\,
            I => n409
        );

    \I__325\ : InMux
    port map (
            O => \N__2180\,
            I => \N__2176\
        );

    \I__324\ : InMux
    port map (
            O => \N__2179\,
            I => \N__2173\
        );

    \I__323\ : LocalMux
    port map (
            O => \N__2176\,
            I => t0on_8
        );

    \I__322\ : LocalMux
    port map (
            O => \N__2173\,
            I => t0on_8
        );

    \I__321\ : InMux
    port map (
            O => \N__2168\,
            I => \N__2165\
        );

    \I__320\ : LocalMux
    port map (
            O => \N__2165\,
            I => \t0on_15_N_35_8\
        );

    \I__319\ : InMux
    port map (
            O => \N__2162\,
            I => \bfn_2_8_0_\
        );

    \I__318\ : InMux
    port map (
            O => \N__2159\,
            I => n411
        );

    \I__317\ : InMux
    port map (
            O => \N__2156\,
            I => n412
        );

    \I__316\ : InMux
    port map (
            O => \N__2153\,
            I => n413
        );

    \I__315\ : InMux
    port map (
            O => \N__2150\,
            I => \N__2147\
        );

    \I__314\ : LocalMux
    port map (
            O => \N__2147\,
            I => n3
        );

    \I__313\ : InMux
    port map (
            O => \N__2144\,
            I => \N__2140\
        );

    \I__312\ : CascadeMux
    port map (
            O => \N__2143\,
            I => \N__2137\
        );

    \I__311\ : LocalMux
    port map (
            O => \N__2140\,
            I => \N__2133\
        );

    \I__310\ : InMux
    port map (
            O => \N__2137\,
            I => \N__2130\
        );

    \I__309\ : InMux
    port map (
            O => \N__2136\,
            I => \N__2127\
        );

    \I__308\ : Span4Mux_v
    port map (
            O => \N__2133\,
            I => \N__2122\
        );

    \I__307\ : LocalMux
    port map (
            O => \N__2130\,
            I => \N__2122\
        );

    \I__306\ : LocalMux
    port map (
            O => \N__2127\,
            I => \N__2119\
        );

    \I__305\ : Span4Mux_v
    port map (
            O => \N__2122\,
            I => \N__2116\
        );

    \I__304\ : Span4Mux_v
    port map (
            O => \N__2119\,
            I => \N__2113\
        );

    \I__303\ : Span4Mux_h
    port map (
            O => \N__2116\,
            I => \N__2108\
        );

    \I__302\ : Span4Mux_h
    port map (
            O => \N__2113\,
            I => \N__2108\
        );

    \I__301\ : Odrv4
    port map (
            O => \N__2108\,
            I => \DIVIDE_1_\
        );

    \I__300\ : InMux
    port map (
            O => \N__2105\,
            I => \N__2102\
        );

    \I__299\ : LocalMux
    port map (
            O => \N__2102\,
            I => \N__2099\
        );

    \I__298\ : Odrv4
    port map (
            O => \N__2099\,
            I => n17
        );

    \I__297\ : CascadeMux
    port map (
            O => \N__2096\,
            I => \N__2093\
        );

    \I__296\ : InMux
    port map (
            O => \N__2093\,
            I => \N__2090\
        );

    \I__295\ : LocalMux
    port map (
            O => \N__2090\,
            I => \N__2086\
        );

    \I__294\ : InMux
    port map (
            O => \N__2089\,
            I => \N__2083\
        );

    \I__293\ : Span4Mux_v
    port map (
            O => \N__2086\,
            I => \N__2079\
        );

    \I__292\ : LocalMux
    port map (
            O => \N__2083\,
            I => \N__2076\
        );

    \I__291\ : InMux
    port map (
            O => \N__2082\,
            I => \N__2073\
        );

    \I__290\ : Span4Mux_h
    port map (
            O => \N__2079\,
            I => \N__2070\
        );

    \I__289\ : Sp12to4
    port map (
            O => \N__2076\,
            I => \N__2065\
        );

    \I__288\ : LocalMux
    port map (
            O => \N__2073\,
            I => \N__2065\
        );

    \I__287\ : Odrv4
    port map (
            O => \N__2070\,
            I => \DIVIDE_7_\
        );

    \I__286\ : Odrv12
    port map (
            O => \N__2065\,
            I => \DIVIDE_7_\
        );

    \I__285\ : CascadeMux
    port map (
            O => \N__2060\,
            I => \N__2057\
        );

    \I__284\ : InMux
    port map (
            O => \N__2057\,
            I => \N__2053\
        );

    \I__283\ : InMux
    port map (
            O => \N__2056\,
            I => \N__2050\
        );

    \I__282\ : LocalMux
    port map (
            O => \N__2053\,
            I => \N__2046\
        );

    \I__281\ : LocalMux
    port map (
            O => \N__2050\,
            I => \N__2043\
        );

    \I__280\ : InMux
    port map (
            O => \N__2049\,
            I => \N__2040\
        );

    \I__279\ : Sp12to4
    port map (
            O => \N__2046\,
            I => \N__2033\
        );

    \I__278\ : Sp12to4
    port map (
            O => \N__2043\,
            I => \N__2033\
        );

    \I__277\ : LocalMux
    port map (
            O => \N__2040\,
            I => \N__2033\
        );

    \I__276\ : Span12Mux_v
    port map (
            O => \N__2033\,
            I => \N__2030\
        );

    \I__275\ : Odrv12
    port map (
            O => \N__2030\,
            I => \DIVIDE_2_\
        );

    \I__274\ : InMux
    port map (
            O => \N__2027\,
            I => \N__2023\
        );

    \I__273\ : InMux
    port map (
            O => \N__2026\,
            I => \N__2020\
        );

    \I__272\ : LocalMux
    port map (
            O => \N__2023\,
            I => t0on_0
        );

    \I__271\ : LocalMux
    port map (
            O => \N__2020\,
            I => t0on_0
        );

    \I__270\ : InMux
    port map (
            O => \N__2015\,
            I => \N__2012\
        );

    \I__269\ : LocalMux
    port map (
            O => \N__2012\,
            I => \t0on_15_N_35_0\
        );

    \I__268\ : InMux
    port map (
            O => \N__2009\,
            I => \bfn_2_7_0_\
        );

    \I__267\ : InMux
    port map (
            O => \N__2006\,
            I => \N__2002\
        );

    \I__266\ : InMux
    port map (
            O => \N__2005\,
            I => \N__1999\
        );

    \I__265\ : LocalMux
    port map (
            O => \N__2002\,
            I => t0on_1
        );

    \I__264\ : LocalMux
    port map (
            O => \N__1999\,
            I => t0on_1
        );

    \I__263\ : InMux
    port map (
            O => \N__1994\,
            I => \N__1991\
        );

    \I__262\ : LocalMux
    port map (
            O => \N__1991\,
            I => \t0on_15_N_35_1\
        );

    \I__261\ : InMux
    port map (
            O => \N__1988\,
            I => n403
        );

    \I__260\ : InMux
    port map (
            O => \N__1985\,
            I => n404
        );

    \I__259\ : InMux
    port map (
            O => \N__1982\,
            I => \N__1978\
        );

    \I__258\ : InMux
    port map (
            O => \N__1981\,
            I => \N__1975\
        );

    \I__257\ : LocalMux
    port map (
            O => \N__1978\,
            I => t0on_3
        );

    \I__256\ : LocalMux
    port map (
            O => \N__1975\,
            I => t0on_3
        );

    \I__255\ : InMux
    port map (
            O => \N__1970\,
            I => \N__1967\
        );

    \I__254\ : LocalMux
    port map (
            O => \N__1967\,
            I => \t0on_15_N_35_3\
        );

    \I__253\ : InMux
    port map (
            O => \N__1964\,
            I => n405
        );

    \I__252\ : CascadeMux
    port map (
            O => \N__1961\,
            I => \N__1958\
        );

    \I__251\ : InMux
    port map (
            O => \N__1958\,
            I => \N__1955\
        );

    \I__250\ : LocalMux
    port map (
            O => \N__1955\,
            I => \N__1952\
        );

    \I__249\ : Odrv4
    port map (
            O => \N__1952\,
            I => n5
        );

    \I__248\ : InMux
    port map (
            O => \N__1949\,
            I => n429
        );

    \I__247\ : CascadeMux
    port map (
            O => \N__1946\,
            I => \N__1943\
        );

    \I__246\ : InMux
    port map (
            O => \N__1943\,
            I => \N__1940\
        );

    \I__245\ : LocalMux
    port map (
            O => \N__1940\,
            I => \N__1937\
        );

    \I__244\ : Odrv4
    port map (
            O => \N__1937\,
            I => n4
        );

    \I__243\ : InMux
    port map (
            O => \N__1934\,
            I => n430
        );

    \I__242\ : CascadeMux
    port map (
            O => \N__1931\,
            I => \N__1928\
        );

    \I__241\ : InMux
    port map (
            O => \N__1928\,
            I => \N__1923\
        );

    \I__240\ : InMux
    port map (
            O => \N__1927\,
            I => \N__1920\
        );

    \I__239\ : InMux
    port map (
            O => \N__1926\,
            I => \N__1917\
        );

    \I__238\ : LocalMux
    port map (
            O => \N__1923\,
            I => \N__1910\
        );

    \I__237\ : LocalMux
    port map (
            O => \N__1920\,
            I => \N__1910\
        );

    \I__236\ : LocalMux
    port map (
            O => \N__1917\,
            I => \N__1910\
        );

    \I__235\ : Span4Mux_v
    port map (
            O => \N__1910\,
            I => \N__1907\
        );

    \I__234\ : Span4Mux_v
    port map (
            O => \N__1907\,
            I => \N__1904\
        );

    \I__233\ : Span4Mux_v
    port map (
            O => \N__1904\,
            I => \N__1901\
        );

    \I__232\ : Sp12to4
    port map (
            O => \N__1901\,
            I => \N__1898\
        );

    \I__231\ : Odrv12
    port map (
            O => \N__1898\,
            I => \DIVIDE_14_\
        );

    \I__230\ : InMux
    port map (
            O => \N__1895\,
            I => n431
        );

    \I__229\ : InMux
    port map (
            O => \N__1892\,
            I => n432
        );

    \I__228\ : CascadeMux
    port map (
            O => \N__1889\,
            I => \N__1886\
        );

    \I__227\ : InMux
    port map (
            O => \N__1886\,
            I => \N__1883\
        );

    \I__226\ : LocalMux
    port map (
            O => \N__1883\,
            I => n7
        );

    \I__225\ : IoInMux
    port map (
            O => \N__1880\,
            I => \N__1877\
        );

    \I__224\ : LocalMux
    port map (
            O => \N__1877\,
            I => \N__1874\
        );

    \I__223\ : Span12Mux_s4_h
    port map (
            O => \N__1874\,
            I => \N__1871\
        );

    \I__222\ : Odrv12
    port map (
            O => \N__1871\,
            I => \OCLK\
        );

    \I__221\ : InMux
    port map (
            O => \N__1868\,
            I => \N__1865\
        );

    \I__220\ : LocalMux
    port map (
            O => \N__1865\,
            I => \N__1862\
        );

    \I__219\ : Odrv4
    port map (
            O => \N__1862\,
            I => n10
        );

    \I__218\ : InMux
    port map (
            O => \N__1859\,
            I => \N__1855\
        );

    \I__217\ : InMux
    port map (
            O => \N__1858\,
            I => \N__1852\
        );

    \I__216\ : LocalMux
    port map (
            O => \N__1855\,
            I => \N__1846\
        );

    \I__215\ : LocalMux
    port map (
            O => \N__1852\,
            I => \N__1846\
        );

    \I__214\ : InMux
    port map (
            O => \N__1851\,
            I => \N__1843\
        );

    \I__213\ : Span4Mux_v
    port map (
            O => \N__1846\,
            I => \N__1838\
        );

    \I__212\ : LocalMux
    port map (
            O => \N__1843\,
            I => \N__1838\
        );

    \I__211\ : Span4Mux_v
    port map (
            O => \N__1838\,
            I => \N__1835\
        );

    \I__210\ : Span4Mux_h
    port map (
            O => \N__1835\,
            I => \N__1832\
        );

    \I__209\ : Odrv4
    port map (
            O => \N__1832\,
            I => \DIVIDE_6_\
        );

    \I__208\ : InMux
    port map (
            O => \N__1829\,
            I => \N__1826\
        );

    \I__207\ : LocalMux
    port map (
            O => \N__1826\,
            I => \N__1823\
        );

    \I__206\ : Odrv4
    port map (
            O => \N__1823\,
            I => n12
        );

    \I__205\ : InMux
    port map (
            O => \N__1820\,
            I => \N__1817\
        );

    \I__204\ : LocalMux
    port map (
            O => \N__1817\,
            I => n14
        );

    \I__203\ : InMux
    port map (
            O => \N__1814\,
            I => n420
        );

    \I__202\ : InMux
    port map (
            O => \N__1811\,
            I => \N__1808\
        );

    \I__201\ : LocalMux
    port map (
            O => \N__1808\,
            I => n13
        );

    \I__200\ : CascadeMux
    port map (
            O => \N__1805\,
            I => \N__1802\
        );

    \I__199\ : InMux
    port map (
            O => \N__1802\,
            I => \N__1799\
        );

    \I__198\ : LocalMux
    port map (
            O => \N__1799\,
            I => \N__1794\
        );

    \I__197\ : InMux
    port map (
            O => \N__1798\,
            I => \N__1791\
        );

    \I__196\ : InMux
    port map (
            O => \N__1797\,
            I => \N__1788\
        );

    \I__195\ : Span4Mux_v
    port map (
            O => \N__1794\,
            I => \N__1781\
        );

    \I__194\ : LocalMux
    port map (
            O => \N__1791\,
            I => \N__1781\
        );

    \I__193\ : LocalMux
    port map (
            O => \N__1788\,
            I => \N__1781\
        );

    \I__192\ : Span4Mux_v
    port map (
            O => \N__1781\,
            I => \N__1778\
        );

    \I__191\ : Span4Mux_h
    port map (
            O => \N__1778\,
            I => \N__1775\
        );

    \I__190\ : Span4Mux_v
    port map (
            O => \N__1775\,
            I => \N__1772\
        );

    \I__189\ : Odrv4
    port map (
            O => \N__1772\,
            I => \DIVIDE_4_\
        );

    \I__188\ : InMux
    port map (
            O => \N__1769\,
            I => n421
        );

    \I__187\ : CascadeMux
    port map (
            O => \N__1766\,
            I => \N__1763\
        );

    \I__186\ : InMux
    port map (
            O => \N__1763\,
            I => \N__1759\
        );

    \I__185\ : InMux
    port map (
            O => \N__1762\,
            I => \N__1756\
        );

    \I__184\ : LocalMux
    port map (
            O => \N__1759\,
            I => \N__1751\
        );

    \I__183\ : LocalMux
    port map (
            O => \N__1756\,
            I => \N__1751\
        );

    \I__182\ : Span4Mux_v
    port map (
            O => \N__1751\,
            I => \N__1747\
        );

    \I__181\ : InMux
    port map (
            O => \N__1750\,
            I => \N__1744\
        );

    \I__180\ : Sp12to4
    port map (
            O => \N__1747\,
            I => \N__1739\
        );

    \I__179\ : LocalMux
    port map (
            O => \N__1744\,
            I => \N__1739\
        );

    \I__178\ : Odrv12
    port map (
            O => \N__1739\,
            I => \DIVIDE_5_\
        );

    \I__177\ : InMux
    port map (
            O => \N__1736\,
            I => n422
        );

    \I__176\ : CascadeMux
    port map (
            O => \N__1733\,
            I => \N__1730\
        );

    \I__175\ : InMux
    port map (
            O => \N__1730\,
            I => \N__1727\
        );

    \I__174\ : LocalMux
    port map (
            O => \N__1727\,
            I => \N__1724\
        );

    \I__173\ : Odrv4
    port map (
            O => \N__1724\,
            I => n11
        );

    \I__172\ : InMux
    port map (
            O => \N__1721\,
            I => n423
        );

    \I__171\ : InMux
    port map (
            O => \N__1718\,
            I => n424
        );

    \I__170\ : CascadeMux
    port map (
            O => \N__1715\,
            I => \N__1712\
        );

    \I__169\ : InMux
    port map (
            O => \N__1712\,
            I => \N__1709\
        );

    \I__168\ : LocalMux
    port map (
            O => \N__1709\,
            I => \N__1706\
        );

    \I__167\ : Odrv4
    port map (
            O => \N__1706\,
            I => n9
        );

    \I__166\ : InMux
    port map (
            O => \N__1703\,
            I => \bfn_1_10_0_\
        );

    \I__165\ : InMux
    port map (
            O => \N__1700\,
            I => \N__1695\
        );

    \I__164\ : InMux
    port map (
            O => \N__1699\,
            I => \N__1692\
        );

    \I__163\ : InMux
    port map (
            O => \N__1698\,
            I => \N__1689\
        );

    \I__162\ : LocalMux
    port map (
            O => \N__1695\,
            I => \N__1686\
        );

    \I__161\ : LocalMux
    port map (
            O => \N__1692\,
            I => \N__1681\
        );

    \I__160\ : LocalMux
    port map (
            O => \N__1689\,
            I => \N__1681\
        );

    \I__159\ : Sp12to4
    port map (
            O => \N__1686\,
            I => \N__1678\
        );

    \I__158\ : Span4Mux_v
    port map (
            O => \N__1681\,
            I => \N__1675\
        );

    \I__157\ : Span12Mux_s5_h
    port map (
            O => \N__1678\,
            I => \N__1670\
        );

    \I__156\ : Sp12to4
    port map (
            O => \N__1675\,
            I => \N__1670\
        );

    \I__155\ : Span12Mux_v
    port map (
            O => \N__1670\,
            I => \N__1667\
        );

    \I__154\ : Odrv12
    port map (
            O => \N__1667\,
            I => \DIVIDE_9_\
        );

    \I__153\ : InMux
    port map (
            O => \N__1664\,
            I => n426
        );

    \I__152\ : InMux
    port map (
            O => \N__1661\,
            I => n427
        );

    \I__151\ : InMux
    port map (
            O => \N__1658\,
            I => n428
        );

    \I__150\ : CascadeMux
    port map (
            O => \N__1655\,
            I => \N__1652\
        );

    \I__149\ : InMux
    port map (
            O => \N__1652\,
            I => \N__1649\
        );

    \I__148\ : LocalMux
    port map (
            O => \N__1649\,
            I => \N__1646\
        );

    \I__147\ : Sp12to4
    port map (
            O => \N__1646\,
            I => \N__1643\
        );

    \I__146\ : Span12Mux_v
    port map (
            O => \N__1643\,
            I => \N__1640\
        );

    \I__145\ : Odrv12
    port map (
            O => \N__1640\,
            I => \DIVIDE_0_\
        );

    \I__144\ : InMux
    port map (
            O => \N__1637\,
            I => \bfn_1_9_0_\
        );

    \I__143\ : InMux
    port map (
            O => \N__1634\,
            I => \N__1631\
        );

    \I__142\ : LocalMux
    port map (
            O => \N__1631\,
            I => n16
        );

    \I__141\ : InMux
    port map (
            O => \N__1628\,
            I => n418
        );

    \I__140\ : InMux
    port map (
            O => \N__1625\,
            I => \N__1622\
        );

    \I__139\ : LocalMux
    port map (
            O => \N__1622\,
            I => n15
        );

    \I__138\ : InMux
    port map (
            O => \N__1619\,
            I => n419
        );

    \IN_MUX_bfv_1_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_9_0_\
        );

    \IN_MUX_bfv_1_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n425,
            carryinitout => \bfn_1_10_0_\
        );

    \IN_MUX_bfv_2_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_9_0_\
        );

    \IN_MUX_bfv_2_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n395,
            carryinitout => \bfn_2_10_0_\
        );

    \IN_MUX_bfv_2_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_7_0_\
        );

    \IN_MUX_bfv_2_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n410,
            carryinitout => \bfn_2_8_0_\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \i200_4_lut_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__2203\,
            in1 => \N__2005\,
            in2 => \N__2255\,
            in3 => \N__2026\,
            lcout => n447,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \t0on_i4_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__1750\,
            in1 => \N__3344\,
            in2 => \_gnd_net_\,
            in3 => \N__2240\,
            lcout => t0on_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3678\,
            ce => \N__3406\,
            sr => \_gnd_net_\
        );

    \sub_34_inv_0_i7_1_lut_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2082\,
            lcout => n11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \t0on_i0_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__2144\,
            in1 => \N__3337\,
            in2 => \_gnd_net_\,
            in3 => \N__2015\,
            lcout => t0on_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3680\,
            ce => \N__3412\,
            sr => \_gnd_net_\
        );

    \t0on_i8_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__3341\,
            in1 => \N__1698\,
            in2 => \_gnd_net_\,
            in3 => \N__2168\,
            lcout => t0on_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3680\,
            ce => \N__3412\,
            sr => \_gnd_net_\
        );

    \t0on_i13_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__3338\,
            in1 => \N__1926\,
            in2 => \_gnd_net_\,
            in3 => \N__2285\,
            lcout => t0on_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3680\,
            ce => \N__3412\,
            sr => \_gnd_net_\
        );

    \t0on_i5_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__1859\,
            in1 => \N__3340\,
            in2 => \_gnd_net_\,
            in3 => \N__2213\,
            lcout => t0on_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3680\,
            ce => \N__3412\,
            sr => \_gnd_net_\
        );

    \t0on_i3_LC_1_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__3339\,
            in1 => \N__1797\,
            in2 => \_gnd_net_\,
            in3 => \N__1970\,
            lcout => t0on_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3680\,
            ce => \N__3412\,
            sr => \_gnd_net_\
        );

    \sub_34_inv_0_i2_1_lut_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__2056\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sub_34_inv_0_i5_1_lut_LC_1_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__1762\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sub_34_inv_0_i13_1_lut_LC_1_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2491\,
            lcout => n5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sub_34_inv_0_i14_1_lut_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__1927\,
            lcout => n4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sub_34_inv_0_i4_1_lut_LC_1_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__1798\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10_4_lut_adj_1_LC_1_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__2296\,
            in1 => \N__1981\,
            in2 => \N__2230\,
            in3 => \N__2179\,
            lcout => n26_adj_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sub_34_inv_0_i9_1_lut_LC_1_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__1699\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sub_34_inv_0_i3_1_lut_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2544\,
            lcout => n15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sub_34_add_2_2_lut_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2105\,
            in2 => \N__1655\,
            in3 => \N__1637\,
            lcout => \t0off_15_N_67_0\,
            ltout => OPEN,
            carryin => \bfn_1_9_0_\,
            carryout => n418,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sub_34_add_2_3_lut_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1634\,
            in2 => \N__2143\,
            in3 => \N__1628\,
            lcout => \t0off_15_N_67_1\,
            ltout => OPEN,
            carryin => n418,
            carryout => n419,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sub_34_add_2_4_lut_LC_1_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1625\,
            in2 => \N__2060\,
            in3 => \N__1619\,
            lcout => \t0off_15_N_67_2\,
            ltout => OPEN,
            carryin => n419,
            carryout => n420,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sub_34_add_2_5_lut_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1820\,
            in2 => \N__2549\,
            in3 => \N__1814\,
            lcout => \t0off_15_N_67_3\,
            ltout => OPEN,
            carryin => n420,
            carryout => n421,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sub_34_add_2_6_lut_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1811\,
            in2 => \N__1805\,
            in3 => \N__1769\,
            lcout => \t0off_15_N_67_4\,
            ltout => OPEN,
            carryin => n421,
            carryout => n422,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sub_34_add_2_7_lut_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1829\,
            in2 => \N__1766\,
            in3 => \N__1736\,
            lcout => \t0off_15_N_67_5\,
            ltout => OPEN,
            carryin => n422,
            carryout => n423,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sub_34_add_2_8_lut_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1858\,
            in2 => \N__1733\,
            in3 => \N__1721\,
            lcout => \t0off_15_N_67_6\,
            ltout => OPEN,
            carryin => n423,
            carryout => n424,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sub_34_add_2_9_lut_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1868\,
            in2 => \N__2096\,
            in3 => \N__1718\,
            lcout => \t0off_15_N_67_7\,
            ltout => OPEN,
            carryin => n424,
            carryout => n425,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sub_34_add_2_10_lut_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2434\,
            in2 => \N__1715\,
            in3 => \N__1703\,
            lcout => \t0off_15_N_67_8\,
            ltout => OPEN,
            carryin => \bfn_1_10_0_\,
            carryout => n426,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sub_34_add_2_11_lut_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1700\,
            in2 => \N__2894\,
            in3 => \N__1664\,
            lcout => \t0off_15_N_67_9\,
            ltout => OPEN,
            carryin => n426,
            carryout => n427,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sub_34_add_2_12_lut_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2908\,
            in2 => \N__1889\,
            in3 => \N__1661\,
            lcout => \t0off_15_N_67_10\,
            ltout => OPEN,
            carryin => n427,
            carryout => n428,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sub_34_add_2_13_lut_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2930\,
            in2 => \N__2609\,
            in3 => \N__1658\,
            lcout => \t0off_15_N_67_11\,
            ltout => OPEN,
            carryin => n428,
            carryout => n429,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sub_34_add_2_14_lut_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2944\,
            in2 => \N__1961\,
            in3 => \N__1949\,
            lcout => \t0off_15_N_67_12\,
            ltout => OPEN,
            carryin => n429,
            carryout => n430,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sub_34_add_2_15_lut_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2495\,
            in2 => \N__1946\,
            in3 => \N__1934\,
            lcout => \t0off_15_N_67_13\,
            ltout => OPEN,
            carryin => n430,
            carryout => n431,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sub_34_add_2_16_lut_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2150\,
            in2 => \N__1931\,
            in3 => \N__1895\,
            lcout => \t0off_15_N_67_14\,
            ltout => OPEN,
            carryin => n431,
            carryout => n432,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \t0off_i15_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100001110100"
        )
    port map (
            in0 => \N__3007\,
            in1 => \N__3402\,
            in2 => \N__2618\,
            in3 => \N__1892\,
            lcout => t0off_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3648\,
            ce => \N__3545\,
            sr => \_gnd_net_\
        );

    \sub_34_inv_0_i11_1_lut_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2607\,
            lcout => n7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \t_clk_24_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3811\,
            lcout => \OCLK\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3614\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sub_34_inv_0_i8_1_lut_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__2433\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sub_34_inv_0_i6_1_lut_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__1851\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => n12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sub_34_inv_0_i15_1_lut_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2994\,
            lcout => n3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sub_34_inv_0_i1_1_lut_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2136\,
            lcout => n17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \t0on_i6_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__3343\,
            in1 => \N__2089\,
            in2 => \_gnd_net_\,
            in3 => \N__2192\,
            lcout => t0on_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3679\,
            ce => \N__3407\,
            sr => \_gnd_net_\
        );

    \t0on_i1_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__2049\,
            in1 => \N__1994\,
            in2 => \_gnd_net_\,
            in3 => \N__3342\,
            lcout => t0on_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3679\,
            ce => \N__3407\,
            sr => \_gnd_net_\
        );

    \add_32_2_lut_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2027\,
            in2 => \_gnd_net_\,
            in3 => \N__2009\,
            lcout => \t0on_15_N_35_0\,
            ltout => OPEN,
            carryin => \bfn_2_7_0_\,
            carryout => n403,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_32_3_lut_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2006\,
            in2 => \N__2768\,
            in3 => \N__1988\,
            lcout => \t0on_15_N_35_1\,
            ltout => OPEN,
            carryin => n403,
            carryout => n404,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_32_4_lut_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2507\,
            in2 => \N__2771\,
            in3 => \N__1985\,
            lcout => \t0on_15_N_35_2\,
            ltout => OPEN,
            carryin => n404,
            carryout => n405,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_32_5_lut_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__1982\,
            in2 => \N__2769\,
            in3 => \N__1964\,
            lcout => \t0on_15_N_35_3\,
            ltout => OPEN,
            carryin => n405,
            carryout => n406,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_32_6_lut_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2254\,
            in2 => \N__2772\,
            in3 => \N__2234\,
            lcout => \t0on_15_N_35_4\,
            ltout => OPEN,
            carryin => n406,
            carryout => n407,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_32_7_lut_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2709\,
            in2 => \N__2231\,
            in3 => \N__2207\,
            lcout => \t0on_15_N_35_5\,
            ltout => OPEN,
            carryin => n407,
            carryout => n408,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_32_8_lut_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2204\,
            in2 => \N__2773\,
            in3 => \N__2186\,
            lcout => \t0on_15_N_35_6\,
            ltout => OPEN,
            carryin => n408,
            carryout => n409,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_32_9_lut_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2386\,
            in2 => \N__2770\,
            in3 => \N__2183\,
            lcout => \t0on_15_N_35_7\,
            ltout => OPEN,
            carryin => n409,
            carryout => n410,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_32_10_lut_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2180\,
            in2 => \N__2774\,
            in3 => \N__2162\,
            lcout => \t0on_15_N_35_8\,
            ltout => OPEN,
            carryin => \bfn_2_8_0_\,
            carryout => n411,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_32_11_lut_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2716\,
            in2 => \N__3023\,
            in3 => \N__2159\,
            lcout => \t0on_15_N_35_9\,
            ltout => OPEN,
            carryin => n411,
            carryout => n412,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_32_12_lut_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2561\,
            in2 => \N__2775\,
            in3 => \N__2156\,
            lcout => \t0on_15_N_35_10\,
            ltout => OPEN,
            carryin => n412,
            carryout => n413,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_32_13_lut_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2720\,
            in2 => \N__2351\,
            in3 => \N__2153\,
            lcout => \t0on_15_N_35_11\,
            ltout => OPEN,
            carryin => n413,
            carryout => n414,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_32_14_lut_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2447\,
            in2 => \N__2776\,
            in3 => \N__2303\,
            lcout => \t0on_15_N_35_12\,
            ltout => OPEN,
            carryin => n414,
            carryout => n415,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_32_15_lut_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2724\,
            in2 => \N__2300\,
            in3 => \N__2279\,
            lcout => \t0on_15_N_35_13\,
            ltout => OPEN,
            carryin => n415,
            carryout => n416,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_32_16_lut_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2969\,
            in2 => \N__2777\,
            in3 => \N__2276\,
            lcout => \t0on_15_N_35_14\,
            ltout => OPEN,
            carryin => n416,
            carryout => n417,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \t0on_i15_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__2371\,
            in1 => \N__2728\,
            in2 => \_gnd_net_\,
            in3 => \N__2273\,
            lcout => t0on_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3681\,
            ce => \N__3413\,
            sr => \N__3425\
        );

    \add_33_2_lut_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3931\,
            in2 => \_gnd_net_\,
            in3 => \N__2270\,
            lcout => \t0off_15_N_51_0\,
            ltout => OPEN,
            carryin => \bfn_2_9_0_\,
            carryout => n388,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_33_3_lut_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3964\,
            in2 => \N__2778\,
            in3 => \N__2267\,
            lcout => \t0off_15_N_51_1\,
            ltout => OPEN,
            carryin => n388,
            carryout => n389,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_33_4_lut_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3220\,
            in2 => \N__2782\,
            in3 => \N__2264\,
            lcout => \t0off_15_N_51_2\,
            ltout => OPEN,
            carryin => n389,
            carryout => n390,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_33_5_lut_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4055\,
            in2 => \N__2779\,
            in3 => \N__2261\,
            lcout => \t0off_15_N_51_3\,
            ltout => OPEN,
            carryin => n390,
            carryout => n391,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_33_6_lut_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3946\,
            in2 => \N__2783\,
            in3 => \N__2258\,
            lcout => \t0off_15_N_51_4\,
            ltout => OPEN,
            carryin => n391,
            carryout => n392,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_33_7_lut_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3890\,
            in2 => \N__2780\,
            in3 => \N__2333\,
            lcout => \t0off_15_N_51_5\,
            ltout => OPEN,
            carryin => n392,
            carryout => n393,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_33_8_lut_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3851\,
            in2 => \N__2784\,
            in3 => \N__2330\,
            lcout => \t0off_15_N_51_6\,
            ltout => OPEN,
            carryin => n393,
            carryout => n394,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_33_9_lut_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3202\,
            in2 => \N__2781\,
            in3 => \N__2327\,
            lcout => \t0off_15_N_51_7\,
            ltout => OPEN,
            carryin => n394,
            carryout => n395,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_33_10_lut_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4039\,
            in2 => \N__2805\,
            in3 => \N__2324\,
            lcout => \t0off_15_N_51_8\,
            ltout => OPEN,
            carryin => \bfn_2_10_0_\,
            carryout => n396,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_33_11_lut_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3986\,
            in2 => \N__2809\,
            in3 => \N__2321\,
            lcout => \t0off_15_N_51_9\,
            ltout => OPEN,
            carryin => n396,
            carryout => n397,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_33_12_lut_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3187\,
            in2 => \N__2806\,
            in3 => \N__2318\,
            lcout => \t0off_15_N_51_10\,
            ltout => OPEN,
            carryin => n397,
            carryout => n398,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_33_13_lut_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3707\,
            in2 => \N__2810\,
            in3 => \N__2315\,
            lcout => \t0off_15_N_51_11\,
            ltout => OPEN,
            carryin => n398,
            carryout => n399,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_33_14_lut_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3235\,
            in2 => \N__2807\,
            in3 => \N__2312\,
            lcout => \t0off_15_N_51_12\,
            ltout => OPEN,
            carryin => n399,
            carryout => n400,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_33_15_lut_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2794\,
            in2 => \N__4073\,
            in3 => \N__2309\,
            lcout => \t0off_15_N_51_13\,
            ltout => OPEN,
            carryin => n400,
            carryout => n401,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_33_16_lut_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4018\,
            in2 => \N__2808\,
            in3 => \N__2306\,
            lcout => \t0off_15_N_51_14\,
            ltout => OPEN,
            carryin => n401,
            carryout => n402,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \add_33_17_lut_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__2804\,
            in1 => \N__4000\,
            in2 => \_gnd_net_\,
            in3 => \N__2621\,
            lcout => \t0off_15_N_51_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i11_4_lut_adj_2_LC_3_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__2446\,
            in1 => \N__2506\,
            in2 => \N__2387\,
            in3 => \N__2560\,
            lcout => n27_adj_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \t0on_i10_LC_3_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__2608\,
            in1 => \N__3333\,
            in2 => \_gnd_net_\,
            in3 => \N__2567\,
            lcout => t0on_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3691\,
            ce => \N__3411\,
            sr => \_gnd_net_\
        );

    \t0on_i2_LC_3_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__3335\,
            in1 => \N__2548\,
            in2 => \_gnd_net_\,
            in3 => \N__2513\,
            lcout => t0on_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3691\,
            ce => \N__3411\,
            sr => \_gnd_net_\
        );

    \t0on_i12_LC_3_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__2490\,
            in1 => \N__3334\,
            in2 => \_gnd_net_\,
            in3 => \N__2453\,
            lcout => t0on_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3691\,
            ce => \N__3411\,
            sr => \_gnd_net_\
        );

    \t0on_i7_LC_3_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__3336\,
            in1 => \N__2435\,
            in2 => \_gnd_net_\,
            in3 => \N__2393\,
            lcout => t0on_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3691\,
            ce => \N__3411\,
            sr => \_gnd_net_\
        );

    \i12_4_lut_LC_3_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__2968\,
            in1 => \N__3019\,
            in2 => \N__2372\,
            in3 => \N__2344\,
            lcout => n28_adj_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \t0on_i11_LC_3_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__2357\,
            in1 => \_gnd_net_\,
            in2 => \N__3324\,
            in3 => \N__2957\,
            lcout => t0on_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3676\,
            ce => \N__3398\,
            sr => \_gnd_net_\
        );

    \t0on_i9_LC_3_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__2918\,
            in1 => \N__3029\,
            in2 => \_gnd_net_\,
            in3 => \N__3298\,
            lcout => t0on_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3676\,
            ce => \N__3398\,
            sr => \_gnd_net_\
        );

    \t0on_i14_LC_3_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__3297\,
            in1 => \N__3008\,
            in2 => \_gnd_net_\,
            in3 => \N__2975\,
            lcout => t0on_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3676\,
            ce => \N__3398\,
            sr => \_gnd_net_\
        );

    \sub_34_inv_0_i12_1_lut_LC_3_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2956\,
            lcout => n6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sub_34_inv_0_i10_1_lut_LC_3_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2917\,
            lcout => n8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \t0off_i3_LC_3_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__2879\,
            in1 => \N__3815\,
            in2 => \_gnd_net_\,
            in3 => \N__2870\,
            lcout => t0off_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3677\,
            ce => \N__3540\,
            sr => \_gnd_net_\
        );

    \t0off_i8_LC_3_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__3817\,
            in1 => \N__2864\,
            in2 => \_gnd_net_\,
            in3 => \N__2852\,
            lcout => t0off_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3677\,
            ce => \N__3540\,
            sr => \_gnd_net_\
        );

    \t0off_i2_LC_3_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__2846\,
            in1 => \N__3814\,
            in2 => \_gnd_net_\,
            in3 => \N__2837\,
            lcout => t0off_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3677\,
            ce => \N__3540\,
            sr => \_gnd_net_\
        );

    \t0off_i10_LC_3_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__3812\,
            in1 => \_gnd_net_\,
            in2 => \N__2831\,
            in3 => \N__2816\,
            lcout => t0off_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3677\,
            ce => \N__3540\,
            sr => \_gnd_net_\
        );

    \t0off_i13_LC_3_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__3161\,
            in1 => \N__3813\,
            in2 => \_gnd_net_\,
            in3 => \N__3149\,
            lcout => t0off_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3677\,
            ce => \N__3540\,
            sr => \_gnd_net_\
        );

    \t0off_i7_LC_3_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__3816\,
            in1 => \N__3143\,
            in2 => \_gnd_net_\,
            in3 => \N__3134\,
            lcout => t0off_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3677\,
            ce => \N__3540\,
            sr => \_gnd_net_\
        );

    \t0off_i12_LC_3_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__3128\,
            in1 => \N__3820\,
            in2 => \_gnd_net_\,
            in3 => \N__3119\,
            lcout => t0off_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3675\,
            ce => \N__3541\,
            sr => \_gnd_net_\
        );

    \t0off_i9_LC_3_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__3824\,
            in1 => \N__3113\,
            in2 => \_gnd_net_\,
            in3 => \N__3107\,
            lcout => t0off_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3675\,
            ce => \N__3541\,
            sr => \_gnd_net_\
        );

    \t0off_i14_LC_3_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__3098\,
            in1 => \N__3821\,
            in2 => \_gnd_net_\,
            in3 => \N__3089\,
            lcout => t0off_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3675\,
            ce => \N__3541\,
            sr => \_gnd_net_\
        );

    \t0off_i4_LC_3_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__3823\,
            in1 => \N__3083\,
            in2 => \_gnd_net_\,
            in3 => \N__3071\,
            lcout => t0off_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3675\,
            ce => \N__3541\,
            sr => \_gnd_net_\
        );

    \t0off_i1_LC_3_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__3065\,
            in1 => \N__3822\,
            in2 => \_gnd_net_\,
            in3 => \N__3053\,
            lcout => t0off_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3675\,
            ce => \N__3541\,
            sr => \_gnd_net_\
        );

    \t0off_i0_LC_3_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__3047\,
            in1 => \N__3035\,
            in2 => \_gnd_net_\,
            in3 => \N__3819\,
            lcout => t0off_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3675\,
            ce => \N__3541\,
            sr => \_gnd_net_\
        );

    \div_state_i1_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3277\,
            in2 => \_gnd_net_\,
            in3 => \N__3762\,
            lcout => div_state_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3692\,
            ce => \N__3443\,
            sr => \_gnd_net_\
        );

    \i206_4_lut_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3494\,
            in1 => \N__3482\,
            in2 => \N__3470\,
            in3 => \N__3458\,
            lcout => n441,
            ltout => \n441_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i214_2_lut_4_lut_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011110111111"
        )
    port map (
            in0 => \N__3757\,
            in1 => \N__3276\,
            in2 => \N__3446\,
            in3 => \N__3169\,
            lcout => n6_adj_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \div_state_i0_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101001111"
        )
    port map (
            in0 => \N__3758\,
            in1 => \N__3431\,
            in2 => \N__3293\,
            in3 => \N__3170\,
            lcout => div_state_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3689\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i217_2_lut_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3271\,
            in2 => \_gnd_net_\,
            in3 => \N__3755\,
            lcout => n386,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i218_1_lut_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__3754\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \div_state_1__N_88\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i208_2_lut_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3272\,
            in2 => \_gnd_net_\,
            in3 => \N__3756\,
            lcout => n307,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i11_4_lut_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3239\,
            in1 => \N__3221\,
            in2 => \N__3206\,
            in3 => \N__3188\,
            lcout => OPEN,
            ltout => \n27_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i205_4_lut_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3971\,
            in1 => \N__4025\,
            in2 => \N__3173\,
            in3 => \N__3917\,
            lcout => n442,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i10_4_lut_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__4072\,
            in1 => \N__4054\,
            in2 => \N__3889\,
            in3 => \N__4040\,
            lcout => n26,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12_4_lut_adj_3_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3703\,
            in1 => \N__4019\,
            in2 => \N__4004\,
            in3 => \N__3985\,
            lcout => n28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i202_4_lut_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__3847\,
            in1 => \N__3965\,
            in2 => \N__3950\,
            in3 => \N__3932\,
            lcout => n444,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \t0off_i5_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__3911\,
            in1 => \N__3780\,
            in2 => \_gnd_net_\,
            in3 => \N__3902\,
            lcout => t0off_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3690\,
            ce => \N__3529\,
            sr => \_gnd_net_\
        );

    \t0off_i6_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__3781\,
            in1 => \N__3869\,
            in2 => \_gnd_net_\,
            in3 => \N__3860\,
            lcout => t0off_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3690\,
            ce => \N__3529\,
            sr => \_gnd_net_\
        );

    \t0off_i11_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__3836\,
            in1 => \N__3818\,
            in2 => \_gnd_net_\,
            in3 => \N__3716\,
            lcout => t0off_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3688\,
            ce => \N__3533\,
            sr => \_gnd_net_\
        );
end \INTERFACE\;
