// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Dec 7 2021 19:29:43

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "zim" view "INTERFACE"

module zim (
    VAC_DRDY,
    IAC_FLT1,
    DDS_SCK,
    ICE_IOR_166,
    ICE_IOR_119,
    DDS_MOSI,
    VAC_MISO,
    DDS_MOSI1,
    ICE_IOR_146,
    VDC_CLK,
    ICE_IOT_222,
    IAC_CS,
    ICE_IOL_18B,
    ICE_IOL_13A,
    ICE_IOB_81,
    VAC_OSR1,
    IAC_MOSI,
    DDS_CS1,
    ICE_IOL_4B,
    ICE_IOB_94,
    VAC_CS,
    VAC_CLK,
    ICE_SPI_CE0,
    ICE_IOR_167,
    ICE_IOR_118,
    RTD_SDO,
    IAC_OSR0,
    VDC_SCLK,
    VAC_FLT1,
    ICE_SPI_MOSI,
    ICE_IOR_165,
    ICE_IOR_147,
    ICE_IOL_14A,
    ICE_IOL_13B,
    ICE_IOB_91,
    ICE_GPMO_0,
    DDS_RNG_0,
    VDC_RNG0,
    ICE_SPI_SCLK,
    ICE_IOR_152,
    ICE_IOL_12A,
    RTD_DRDY,
    ICE_SPI_MISO,
    ICE_IOT_177,
    ICE_IOR_141,
    ICE_IOB_80,
    ICE_IOB_102,
    ICE_GPMO_2,
    ICE_GPMI_0,
    IAC_MISO,
    VAC_OSR0,
    VAC_MOSI,
    TEST_LED,
    ICE_IOR_148,
    STAT_COMM,
    ICE_SYSCLK,
    ICE_IOR_161,
    ICE_IOB_95,
    ICE_IOB_82,
    ICE_IOB_104,
    IAC_CLK,
    DDS_CS,
    SELIRNG0,
    RTD_SDI,
    ICE_IOT_221,
    ICE_IOT_197,
    DDS_MCLK,
    RTD_SCLK,
    RTD_CS,
    ICE_IOR_137,
    IAC_OSR1,
    VAC_FLT0,
    ICE_IOR_144,
    ICE_IOR_128,
    ICE_GPMO_1,
    IAC_SCLK,
    EIS_SYNCCLK,
    ICE_IOR_139,
    ICE_IOL_4A,
    VAC_SCLK,
    THERMOSTAT,
    ICE_IOR_164,
    ICE_IOB_103,
    AMPV_POW,
    VDC_SDO,
    ICE_IOT_174,
    ICE_IOR_140,
    ICE_IOB_96,
    CONT_SD,
    AC_ADC_SYNC,
    SELIRNG1,
    ICE_IOL_12B,
    ICE_IOR_160,
    ICE_IOR_136,
    DDS_MCLK1,
    ICE_IOT_198,
    ICE_IOT_173,
    IAC_DRDY,
    ICE_IOT_178,
    ICE_IOR_138,
    ICE_IOR_120,
    IAC_FLT0,
    DDS_SCK1);

    input VAC_DRDY;
    output IAC_FLT1;
    output DDS_SCK;
    input ICE_IOR_166;
    input ICE_IOR_119;
    output DDS_MOSI;
    input VAC_MISO;
    output DDS_MOSI1;
    input ICE_IOR_146;
    output VDC_CLK;
    input ICE_IOT_222;
    output IAC_CS;
    input ICE_IOL_18B;
    input ICE_IOL_13A;
    input ICE_IOB_81;
    output VAC_OSR1;
    output IAC_MOSI;
    output DDS_CS1;
    input ICE_IOL_4B;
    input ICE_IOB_94;
    output VAC_CS;
    output VAC_CLK;
    input ICE_SPI_CE0;
    input ICE_IOR_167;
    input ICE_IOR_118;
    input RTD_SDO;
    output IAC_OSR0;
    output VDC_SCLK;
    output VAC_FLT1;
    input ICE_SPI_MOSI;
    input ICE_IOR_165;
    input ICE_IOR_147;
    input ICE_IOL_14A;
    input ICE_IOL_13B;
    input ICE_IOB_91;
    input ICE_GPMO_0;
    output DDS_RNG_0;
    output VDC_RNG0;
    input ICE_SPI_SCLK;
    input ICE_IOR_152;
    input ICE_IOL_12A;
    input RTD_DRDY;
    output ICE_SPI_MISO;
    input ICE_IOT_177;
    input ICE_IOR_141;
    input ICE_IOB_80;
    input ICE_IOB_102;
    input ICE_GPMO_2;
    output ICE_GPMI_0;
    input IAC_MISO;
    output VAC_OSR0;
    output VAC_MOSI;
    output TEST_LED;
    input ICE_IOR_148;
    output STAT_COMM;
    input ICE_SYSCLK;
    input ICE_IOR_161;
    input ICE_IOB_95;
    input ICE_IOB_82;
    input ICE_IOB_104;
    output IAC_CLK;
    output DDS_CS;
    output SELIRNG0;
    output RTD_SDI;
    input ICE_IOT_221;
    input ICE_IOT_197;
    output DDS_MCLK;
    output RTD_SCLK;
    output RTD_CS;
    input ICE_IOR_137;
    output IAC_OSR1;
    output VAC_FLT0;
    input ICE_IOR_144;
    input ICE_IOR_128;
    input ICE_GPMO_1;
    output IAC_SCLK;
    input EIS_SYNCCLK;
    input ICE_IOR_139;
    input ICE_IOL_4A;
    output VAC_SCLK;
    input THERMOSTAT;
    input ICE_IOR_164;
    input ICE_IOB_103;
    output AMPV_POW;
    input VDC_SDO;
    input ICE_IOT_174;
    input ICE_IOR_140;
    input ICE_IOB_96;
    output CONT_SD;
    output AC_ADC_SYNC;
    output SELIRNG1;
    input ICE_IOL_12B;
    input ICE_IOR_160;
    input ICE_IOR_136;
    output DDS_MCLK1;
    input ICE_IOT_198;
    input ICE_IOT_173;
    input IAC_DRDY;
    input ICE_IOT_178;
    input ICE_IOR_138;
    input ICE_IOR_120;
    output IAC_FLT0;
    output DDS_SCK1;

    wire N__59914;
    wire N__59913;
    wire N__59912;
    wire N__59905;
    wire N__59904;
    wire N__59903;
    wire N__59896;
    wire N__59895;
    wire N__59894;
    wire N__59887;
    wire N__59886;
    wire N__59885;
    wire N__59878;
    wire N__59877;
    wire N__59876;
    wire N__59869;
    wire N__59868;
    wire N__59867;
    wire N__59860;
    wire N__59859;
    wire N__59858;
    wire N__59851;
    wire N__59850;
    wire N__59849;
    wire N__59842;
    wire N__59841;
    wire N__59840;
    wire N__59833;
    wire N__59832;
    wire N__59831;
    wire N__59824;
    wire N__59823;
    wire N__59822;
    wire N__59815;
    wire N__59814;
    wire N__59813;
    wire N__59806;
    wire N__59805;
    wire N__59804;
    wire N__59797;
    wire N__59796;
    wire N__59795;
    wire N__59788;
    wire N__59787;
    wire N__59786;
    wire N__59779;
    wire N__59778;
    wire N__59777;
    wire N__59770;
    wire N__59769;
    wire N__59768;
    wire N__59761;
    wire N__59760;
    wire N__59759;
    wire N__59752;
    wire N__59751;
    wire N__59750;
    wire N__59743;
    wire N__59742;
    wire N__59741;
    wire N__59734;
    wire N__59733;
    wire N__59732;
    wire N__59725;
    wire N__59724;
    wire N__59723;
    wire N__59716;
    wire N__59715;
    wire N__59714;
    wire N__59707;
    wire N__59706;
    wire N__59705;
    wire N__59698;
    wire N__59697;
    wire N__59696;
    wire N__59689;
    wire N__59688;
    wire N__59687;
    wire N__59680;
    wire N__59679;
    wire N__59678;
    wire N__59671;
    wire N__59670;
    wire N__59669;
    wire N__59662;
    wire N__59661;
    wire N__59660;
    wire N__59653;
    wire N__59652;
    wire N__59651;
    wire N__59644;
    wire N__59643;
    wire N__59642;
    wire N__59635;
    wire N__59634;
    wire N__59633;
    wire N__59626;
    wire N__59625;
    wire N__59624;
    wire N__59617;
    wire N__59616;
    wire N__59615;
    wire N__59608;
    wire N__59607;
    wire N__59606;
    wire N__59599;
    wire N__59598;
    wire N__59597;
    wire N__59590;
    wire N__59589;
    wire N__59588;
    wire N__59581;
    wire N__59580;
    wire N__59579;
    wire N__59572;
    wire N__59571;
    wire N__59570;
    wire N__59563;
    wire N__59562;
    wire N__59561;
    wire N__59554;
    wire N__59553;
    wire N__59552;
    wire N__59545;
    wire N__59544;
    wire N__59543;
    wire N__59536;
    wire N__59535;
    wire N__59534;
    wire N__59527;
    wire N__59526;
    wire N__59525;
    wire N__59518;
    wire N__59517;
    wire N__59516;
    wire N__59509;
    wire N__59508;
    wire N__59507;
    wire N__59500;
    wire N__59499;
    wire N__59498;
    wire N__59491;
    wire N__59490;
    wire N__59489;
    wire N__59482;
    wire N__59481;
    wire N__59480;
    wire N__59473;
    wire N__59472;
    wire N__59471;
    wire N__59464;
    wire N__59463;
    wire N__59462;
    wire N__59455;
    wire N__59454;
    wire N__59453;
    wire N__59446;
    wire N__59445;
    wire N__59444;
    wire N__59437;
    wire N__59436;
    wire N__59435;
    wire N__59428;
    wire N__59427;
    wire N__59426;
    wire N__59419;
    wire N__59418;
    wire N__59417;
    wire N__59410;
    wire N__59409;
    wire N__59408;
    wire N__59401;
    wire N__59400;
    wire N__59399;
    wire N__59392;
    wire N__59391;
    wire N__59390;
    wire N__59383;
    wire N__59382;
    wire N__59381;
    wire N__59374;
    wire N__59373;
    wire N__59372;
    wire N__59365;
    wire N__59364;
    wire N__59363;
    wire N__59356;
    wire N__59355;
    wire N__59354;
    wire N__59347;
    wire N__59346;
    wire N__59345;
    wire N__59338;
    wire N__59337;
    wire N__59336;
    wire N__59329;
    wire N__59328;
    wire N__59327;
    wire N__59320;
    wire N__59319;
    wire N__59318;
    wire N__59311;
    wire N__59310;
    wire N__59309;
    wire N__59302;
    wire N__59301;
    wire N__59300;
    wire N__59293;
    wire N__59292;
    wire N__59291;
    wire N__59284;
    wire N__59283;
    wire N__59282;
    wire N__59275;
    wire N__59274;
    wire N__59273;
    wire N__59266;
    wire N__59265;
    wire N__59264;
    wire N__59257;
    wire N__59256;
    wire N__59255;
    wire N__59248;
    wire N__59247;
    wire N__59246;
    wire N__59239;
    wire N__59238;
    wire N__59237;
    wire N__59230;
    wire N__59229;
    wire N__59228;
    wire N__59221;
    wire N__59220;
    wire N__59219;
    wire N__59212;
    wire N__59211;
    wire N__59210;
    wire N__59203;
    wire N__59202;
    wire N__59201;
    wire N__59194;
    wire N__59193;
    wire N__59192;
    wire N__59185;
    wire N__59184;
    wire N__59183;
    wire N__59176;
    wire N__59175;
    wire N__59174;
    wire N__59167;
    wire N__59166;
    wire N__59165;
    wire N__59158;
    wire N__59157;
    wire N__59156;
    wire N__59149;
    wire N__59148;
    wire N__59147;
    wire N__59140;
    wire N__59139;
    wire N__59138;
    wire N__59131;
    wire N__59130;
    wire N__59129;
    wire N__59122;
    wire N__59121;
    wire N__59120;
    wire N__59113;
    wire N__59112;
    wire N__59111;
    wire N__59104;
    wire N__59103;
    wire N__59102;
    wire N__59095;
    wire N__59094;
    wire N__59093;
    wire N__59086;
    wire N__59085;
    wire N__59084;
    wire N__59077;
    wire N__59076;
    wire N__59075;
    wire N__59068;
    wire N__59067;
    wire N__59066;
    wire N__59059;
    wire N__59058;
    wire N__59057;
    wire N__59050;
    wire N__59049;
    wire N__59048;
    wire N__59041;
    wire N__59040;
    wire N__59039;
    wire N__59032;
    wire N__59031;
    wire N__59030;
    wire N__59023;
    wire N__59022;
    wire N__59021;
    wire N__59014;
    wire N__59013;
    wire N__59012;
    wire N__59005;
    wire N__59004;
    wire N__59003;
    wire N__58996;
    wire N__58995;
    wire N__58994;
    wire N__58977;
    wire N__58974;
    wire N__58973;
    wire N__58972;
    wire N__58969;
    wire N__58968;
    wire N__58965;
    wire N__58962;
    wire N__58959;
    wire N__58956;
    wire N__58953;
    wire N__58950;
    wire N__58945;
    wire N__58942;
    wire N__58939;
    wire N__58934;
    wire N__58931;
    wire N__58926;
    wire N__58923;
    wire N__58920;
    wire N__58917;
    wire N__58914;
    wire N__58911;
    wire N__58910;
    wire N__58907;
    wire N__58904;
    wire N__58899;
    wire N__58896;
    wire N__58893;
    wire N__58892;
    wire N__58891;
    wire N__58888;
    wire N__58885;
    wire N__58882;
    wire N__58875;
    wire N__58874;
    wire N__58871;
    wire N__58868;
    wire N__58863;
    wire N__58860;
    wire N__58857;
    wire N__58856;
    wire N__58853;
    wire N__58850;
    wire N__58847;
    wire N__58844;
    wire N__58839;
    wire N__58836;
    wire N__58833;
    wire N__58830;
    wire N__58827;
    wire N__58824;
    wire N__58821;
    wire N__58818;
    wire N__58817;
    wire N__58816;
    wire N__58809;
    wire N__58806;
    wire N__58803;
    wire N__58800;
    wire N__58797;
    wire N__58796;
    wire N__58793;
    wire N__58790;
    wire N__58789;
    wire N__58784;
    wire N__58781;
    wire N__58776;
    wire N__58775;
    wire N__58774;
    wire N__58773;
    wire N__58770;
    wire N__58767;
    wire N__58766;
    wire N__58765;
    wire N__58764;
    wire N__58763;
    wire N__58762;
    wire N__58759;
    wire N__58758;
    wire N__58755;
    wire N__58754;
    wire N__58753;
    wire N__58752;
    wire N__58751;
    wire N__58750;
    wire N__58749;
    wire N__58748;
    wire N__58747;
    wire N__58746;
    wire N__58745;
    wire N__58744;
    wire N__58743;
    wire N__58738;
    wire N__58735;
    wire N__58732;
    wire N__58729;
    wire N__58728;
    wire N__58725;
    wire N__58722;
    wire N__58721;
    wire N__58720;
    wire N__58719;
    wire N__58718;
    wire N__58717;
    wire N__58716;
    wire N__58715;
    wire N__58712;
    wire N__58709;
    wire N__58708;
    wire N__58707;
    wire N__58706;
    wire N__58705;
    wire N__58704;
    wire N__58703;
    wire N__58702;
    wire N__58699;
    wire N__58696;
    wire N__58695;
    wire N__58692;
    wire N__58691;
    wire N__58688;
    wire N__58687;
    wire N__58684;
    wire N__58683;
    wire N__58680;
    wire N__58679;
    wire N__58676;
    wire N__58675;
    wire N__58672;
    wire N__58671;
    wire N__58668;
    wire N__58665;
    wire N__58664;
    wire N__58661;
    wire N__58660;
    wire N__58657;
    wire N__58656;
    wire N__58653;
    wire N__58644;
    wire N__58641;
    wire N__58636;
    wire N__58633;
    wire N__58630;
    wire N__58627;
    wire N__58626;
    wire N__58623;
    wire N__58622;
    wire N__58619;
    wire N__58618;
    wire N__58615;
    wire N__58614;
    wire N__58611;
    wire N__58608;
    wire N__58605;
    wire N__58598;
    wire N__58589;
    wire N__58586;
    wire N__58571;
    wire N__58554;
    wire N__58539;
    wire N__58534;
    wire N__58525;
    wire N__58508;
    wire N__58503;
    wire N__58498;
    wire N__58495;
    wire N__58490;
    wire N__58487;
    wire N__58486;
    wire N__58481;
    wire N__58478;
    wire N__58475;
    wire N__58472;
    wire N__58469;
    wire N__58466;
    wire N__58463;
    wire N__58460;
    wire N__58455;
    wire N__58450;
    wire N__58441;
    wire N__58438;
    wire N__58431;
    wire N__58430;
    wire N__58427;
    wire N__58424;
    wire N__58421;
    wire N__58418;
    wire N__58413;
    wire N__58412;
    wire N__58409;
    wire N__58408;
    wire N__58407;
    wire N__58406;
    wire N__58403;
    wire N__58402;
    wire N__58401;
    wire N__58400;
    wire N__58399;
    wire N__58396;
    wire N__58393;
    wire N__58392;
    wire N__58391;
    wire N__58388;
    wire N__58385;
    wire N__58384;
    wire N__58381;
    wire N__58378;
    wire N__58375;
    wire N__58372;
    wire N__58371;
    wire N__58368;
    wire N__58367;
    wire N__58362;
    wire N__58359;
    wire N__58358;
    wire N__58357;
    wire N__58356;
    wire N__58353;
    wire N__58352;
    wire N__58347;
    wire N__58344;
    wire N__58341;
    wire N__58338;
    wire N__58337;
    wire N__58332;
    wire N__58329;
    wire N__58328;
    wire N__58325;
    wire N__58322;
    wire N__58317;
    wire N__58314;
    wire N__58311;
    wire N__58308;
    wire N__58307;
    wire N__58304;
    wire N__58301;
    wire N__58298;
    wire N__58295;
    wire N__58290;
    wire N__58287;
    wire N__58284;
    wire N__58281;
    wire N__58278;
    wire N__58273;
    wire N__58270;
    wire N__58267;
    wire N__58264;
    wire N__58261;
    wire N__58258;
    wire N__58257;
    wire N__58252;
    wire N__58243;
    wire N__58236;
    wire N__58231;
    wire N__58222;
    wire N__58219;
    wire N__58216;
    wire N__58211;
    wire N__58206;
    wire N__58203;
    wire N__58194;
    wire N__58193;
    wire N__58192;
    wire N__58187;
    wire N__58184;
    wire N__58181;
    wire N__58178;
    wire N__58173;
    wire N__58170;
    wire N__58167;
    wire N__58166;
    wire N__58165;
    wire N__58164;
    wire N__58163;
    wire N__58162;
    wire N__58161;
    wire N__58160;
    wire N__58159;
    wire N__58158;
    wire N__58157;
    wire N__58156;
    wire N__58153;
    wire N__58150;
    wire N__58149;
    wire N__58146;
    wire N__58145;
    wire N__58140;
    wire N__58139;
    wire N__58136;
    wire N__58133;
    wire N__58132;
    wire N__58131;
    wire N__58128;
    wire N__58127;
    wire N__58126;
    wire N__58123;
    wire N__58122;
    wire N__58121;
    wire N__58120;
    wire N__58117;
    wire N__58114;
    wire N__58113;
    wire N__58110;
    wire N__58109;
    wire N__58108;
    wire N__58101;
    wire N__58098;
    wire N__58095;
    wire N__58092;
    wire N__58081;
    wire N__58074;
    wire N__58071;
    wire N__58068;
    wire N__58067;
    wire N__58066;
    wire N__58065;
    wire N__58060;
    wire N__58059;
    wire N__58058;
    wire N__58055;
    wire N__58054;
    wire N__58053;
    wire N__58052;
    wire N__58051;
    wire N__58048;
    wire N__58045;
    wire N__58038;
    wire N__58035;
    wire N__58030;
    wire N__58023;
    wire N__58018;
    wire N__58013;
    wire N__58010;
    wire N__58007;
    wire N__58002;
    wire N__57999;
    wire N__57994;
    wire N__57989;
    wire N__57988;
    wire N__57987;
    wire N__57982;
    wire N__57979;
    wire N__57976;
    wire N__57973;
    wire N__57970;
    wire N__57967;
    wire N__57960;
    wire N__57957;
    wire N__57950;
    wire N__57945;
    wire N__57940;
    wire N__57935;
    wire N__57932;
    wire N__57929;
    wire N__57926;
    wire N__57919;
    wire N__57916;
    wire N__57903;
    wire N__57900;
    wire N__57897;
    wire N__57896;
    wire N__57893;
    wire N__57890;
    wire N__57887;
    wire N__57882;
    wire N__57879;
    wire N__57878;
    wire N__57875;
    wire N__57872;
    wire N__57869;
    wire N__57866;
    wire N__57861;
    wire N__57858;
    wire N__57855;
    wire N__57854;
    wire N__57851;
    wire N__57848;
    wire N__57845;
    wire N__57840;
    wire N__57837;
    wire N__57836;
    wire N__57833;
    wire N__57830;
    wire N__57827;
    wire N__57824;
    wire N__57819;
    wire N__57816;
    wire N__57813;
    wire N__57812;
    wire N__57809;
    wire N__57806;
    wire N__57803;
    wire N__57798;
    wire N__57795;
    wire N__57794;
    wire N__57791;
    wire N__57788;
    wire N__57785;
    wire N__57782;
    wire N__57777;
    wire N__57774;
    wire N__57773;
    wire N__57770;
    wire N__57767;
    wire N__57764;
    wire N__57759;
    wire N__57756;
    wire N__57753;
    wire N__57750;
    wire N__57749;
    wire N__57746;
    wire N__57743;
    wire N__57740;
    wire N__57735;
    wire N__57734;
    wire N__57731;
    wire N__57728;
    wire N__57725;
    wire N__57722;
    wire N__57719;
    wire N__57714;
    wire N__57713;
    wire N__57710;
    wire N__57707;
    wire N__57704;
    wire N__57699;
    wire N__57696;
    wire N__57695;
    wire N__57692;
    wire N__57689;
    wire N__57686;
    wire N__57681;
    wire N__57678;
    wire N__57677;
    wire N__57674;
    wire N__57671;
    wire N__57668;
    wire N__57665;
    wire N__57660;
    wire N__57657;
    wire N__57654;
    wire N__57653;
    wire N__57650;
    wire N__57647;
    wire N__57644;
    wire N__57639;
    wire N__57636;
    wire N__57635;
    wire N__57632;
    wire N__57629;
    wire N__57626;
    wire N__57623;
    wire N__57620;
    wire N__57615;
    wire N__57612;
    wire N__57609;
    wire N__57606;
    wire N__57605;
    wire N__57602;
    wire N__57599;
    wire N__57596;
    wire N__57591;
    wire N__57588;
    wire N__57587;
    wire N__57584;
    wire N__57581;
    wire N__57578;
    wire N__57575;
    wire N__57570;
    wire N__57567;
    wire N__57564;
    wire N__57563;
    wire N__57560;
    wire N__57557;
    wire N__57554;
    wire N__57549;
    wire N__57546;
    wire N__57543;
    wire N__57540;
    wire N__57537;
    wire N__57536;
    wire N__57535;
    wire N__57532;
    wire N__57529;
    wire N__57526;
    wire N__57519;
    wire N__57516;
    wire N__57515;
    wire N__57512;
    wire N__57509;
    wire N__57506;
    wire N__57503;
    wire N__57500;
    wire N__57497;
    wire N__57492;
    wire N__57491;
    wire N__57488;
    wire N__57485;
    wire N__57482;
    wire N__57479;
    wire N__57474;
    wire N__57471;
    wire N__57470;
    wire N__57467;
    wire N__57464;
    wire N__57459;
    wire N__57456;
    wire N__57453;
    wire N__57450;
    wire N__57447;
    wire N__57444;
    wire N__57441;
    wire N__57438;
    wire N__57437;
    wire N__57434;
    wire N__57431;
    wire N__57430;
    wire N__57425;
    wire N__57422;
    wire N__57417;
    wire N__57414;
    wire N__57413;
    wire N__57410;
    wire N__57407;
    wire N__57402;
    wire N__57399;
    wire N__57396;
    wire N__57395;
    wire N__57392;
    wire N__57389;
    wire N__57386;
    wire N__57383;
    wire N__57378;
    wire N__57375;
    wire N__57372;
    wire N__57371;
    wire N__57368;
    wire N__57365;
    wire N__57362;
    wire N__57359;
    wire N__57354;
    wire N__57351;
    wire N__57348;
    wire N__57345;
    wire N__57342;
    wire N__57339;
    wire N__57336;
    wire N__57333;
    wire N__57330;
    wire N__57327;
    wire N__57324;
    wire N__57321;
    wire N__57318;
    wire N__57315;
    wire N__57312;
    wire N__57309;
    wire N__57306;
    wire N__57303;
    wire N__57300;
    wire N__57297;
    wire N__57294;
    wire N__57291;
    wire N__57288;
    wire N__57285;
    wire N__57282;
    wire N__57279;
    wire N__57276;
    wire N__57273;
    wire N__57272;
    wire N__57271;
    wire N__57270;
    wire N__57269;
    wire N__57268;
    wire N__57267;
    wire N__57266;
    wire N__57265;
    wire N__57264;
    wire N__57263;
    wire N__57262;
    wire N__57261;
    wire N__57260;
    wire N__57259;
    wire N__57258;
    wire N__57257;
    wire N__57254;
    wire N__57253;
    wire N__57252;
    wire N__57251;
    wire N__57250;
    wire N__57249;
    wire N__57246;
    wire N__57243;
    wire N__57240;
    wire N__57239;
    wire N__57238;
    wire N__57233;
    wire N__57230;
    wire N__57227;
    wire N__57224;
    wire N__57221;
    wire N__57218;
    wire N__57217;
    wire N__57214;
    wire N__57213;
    wire N__57212;
    wire N__57211;
    wire N__57210;
    wire N__57209;
    wire N__57208;
    wire N__57207;
    wire N__57206;
    wire N__57205;
    wire N__57204;
    wire N__57203;
    wire N__57202;
    wire N__57199;
    wire N__57198;
    wire N__57197;
    wire N__57196;
    wire N__57195;
    wire N__57194;
    wire N__57191;
    wire N__57188;
    wire N__57187;
    wire N__57186;
    wire N__57185;
    wire N__57184;
    wire N__57181;
    wire N__57180;
    wire N__57179;
    wire N__57170;
    wire N__57167;
    wire N__57164;
    wire N__57163;
    wire N__57162;
    wire N__57159;
    wire N__57152;
    wire N__57151;
    wire N__57150;
    wire N__57149;
    wire N__57148;
    wire N__57147;
    wire N__57146;
    wire N__57143;
    wire N__57140;
    wire N__57137;
    wire N__57136;
    wire N__57135;
    wire N__57134;
    wire N__57133;
    wire N__57132;
    wire N__57131;
    wire N__57130;
    wire N__57129;
    wire N__57128;
    wire N__57127;
    wire N__57122;
    wire N__57115;
    wire N__57114;
    wire N__57113;
    wire N__57112;
    wire N__57111;
    wire N__57110;
    wire N__57109;
    wire N__57106;
    wire N__57105;
    wire N__57102;
    wire N__57101;
    wire N__57100;
    wire N__57099;
    wire N__57098;
    wire N__57097;
    wire N__57094;
    wire N__57093;
    wire N__57092;
    wire N__57091;
    wire N__57088;
    wire N__57083;
    wire N__57080;
    wire N__57077;
    wire N__57072;
    wire N__57067;
    wire N__57062;
    wire N__57059;
    wire N__57052;
    wire N__57049;
    wire N__57046;
    wire N__57043;
    wire N__57038;
    wire N__57035;
    wire N__57032;
    wire N__57029;
    wire N__57028;
    wire N__57027;
    wire N__57026;
    wire N__57025;
    wire N__57024;
    wire N__57023;
    wire N__57018;
    wire N__57015;
    wire N__57012;
    wire N__57007;
    wire N__57004;
    wire N__56999;
    wire N__56996;
    wire N__56993;
    wire N__56986;
    wire N__56983;
    wire N__56980;
    wire N__56975;
    wire N__56972;
    wire N__56961;
    wire N__56960;
    wire N__56959;
    wire N__56958;
    wire N__56957;
    wire N__56954;
    wire N__56949;
    wire N__56946;
    wire N__56943;
    wire N__56938;
    wire N__56937;
    wire N__56934;
    wire N__56931;
    wire N__56928;
    wire N__56925;
    wire N__56918;
    wire N__56915;
    wire N__56914;
    wire N__56913;
    wire N__56910;
    wire N__56901;
    wire N__56900;
    wire N__56899;
    wire N__56898;
    wire N__56895;
    wire N__56892;
    wire N__56889;
    wire N__56884;
    wire N__56881;
    wire N__56878;
    wire N__56875;
    wire N__56874;
    wire N__56873;
    wire N__56870;
    wire N__56869;
    wire N__56868;
    wire N__56867;
    wire N__56866;
    wire N__56865;
    wire N__56856;
    wire N__56853;
    wire N__56848;
    wire N__56843;
    wire N__56836;
    wire N__56827;
    wire N__56822;
    wire N__56807;
    wire N__56802;
    wire N__56791;
    wire N__56788;
    wire N__56787;
    wire N__56784;
    wire N__56783;
    wire N__56778;
    wire N__56767;
    wire N__56764;
    wire N__56753;
    wire N__56752;
    wire N__56751;
    wire N__56748;
    wire N__56743;
    wire N__56738;
    wire N__56731;
    wire N__56728;
    wire N__56723;
    wire N__56720;
    wire N__56713;
    wire N__56710;
    wire N__56707;
    wire N__56704;
    wire N__56697;
    wire N__56692;
    wire N__56687;
    wire N__56680;
    wire N__56669;
    wire N__56660;
    wire N__56655;
    wire N__56650;
    wire N__56645;
    wire N__56628;
    wire N__56601;
    wire N__56598;
    wire N__56595;
    wire N__56592;
    wire N__56589;
    wire N__56586;
    wire N__56583;
    wire N__56582;
    wire N__56579;
    wire N__56578;
    wire N__56575;
    wire N__56574;
    wire N__56573;
    wire N__56572;
    wire N__56571;
    wire N__56568;
    wire N__56565;
    wire N__56562;
    wire N__56557;
    wire N__56552;
    wire N__56541;
    wire N__56538;
    wire N__56537;
    wire N__56534;
    wire N__56531;
    wire N__56526;
    wire N__56523;
    wire N__56520;
    wire N__56517;
    wire N__56514;
    wire N__56511;
    wire N__56508;
    wire N__56505;
    wire N__56504;
    wire N__56503;
    wire N__56500;
    wire N__56497;
    wire N__56494;
    wire N__56487;
    wire N__56486;
    wire N__56483;
    wire N__56480;
    wire N__56477;
    wire N__56474;
    wire N__56469;
    wire N__56466;
    wire N__56463;
    wire N__56460;
    wire N__56457;
    wire N__56454;
    wire N__56451;
    wire N__56448;
    wire N__56447;
    wire N__56446;
    wire N__56443;
    wire N__56438;
    wire N__56435;
    wire N__56432;
    wire N__56429;
    wire N__56426;
    wire N__56421;
    wire N__56418;
    wire N__56415;
    wire N__56412;
    wire N__56409;
    wire N__56406;
    wire N__56403;
    wire N__56402;
    wire N__56401;
    wire N__56394;
    wire N__56391;
    wire N__56388;
    wire N__56385;
    wire N__56382;
    wire N__56381;
    wire N__56378;
    wire N__56375;
    wire N__56370;
    wire N__56369;
    wire N__56366;
    wire N__56363;
    wire N__56358;
    wire N__56357;
    wire N__56354;
    wire N__56351;
    wire N__56348;
    wire N__56345;
    wire N__56340;
    wire N__56339;
    wire N__56336;
    wire N__56333;
    wire N__56328;
    wire N__56325;
    wire N__56322;
    wire N__56319;
    wire N__56316;
    wire N__56313;
    wire N__56310;
    wire N__56307;
    wire N__56304;
    wire N__56301;
    wire N__56298;
    wire N__56297;
    wire N__56294;
    wire N__56291;
    wire N__56288;
    wire N__56285;
    wire N__56280;
    wire N__56279;
    wire N__56276;
    wire N__56273;
    wire N__56270;
    wire N__56265;
    wire N__56264;
    wire N__56261;
    wire N__56258;
    wire N__56255;
    wire N__56250;
    wire N__56249;
    wire N__56246;
    wire N__56243;
    wire N__56238;
    wire N__56235;
    wire N__56232;
    wire N__56231;
    wire N__56230;
    wire N__56229;
    wire N__56228;
    wire N__56225;
    wire N__56222;
    wire N__56217;
    wire N__56214;
    wire N__56205;
    wire N__56202;
    wire N__56199;
    wire N__56198;
    wire N__56195;
    wire N__56192;
    wire N__56187;
    wire N__56184;
    wire N__56181;
    wire N__56180;
    wire N__56177;
    wire N__56174;
    wire N__56169;
    wire N__56168;
    wire N__56165;
    wire N__56162;
    wire N__56159;
    wire N__56154;
    wire N__56151;
    wire N__56148;
    wire N__56147;
    wire N__56144;
    wire N__56141;
    wire N__56140;
    wire N__56135;
    wire N__56132;
    wire N__56129;
    wire N__56126;
    wire N__56121;
    wire N__56118;
    wire N__56115;
    wire N__56112;
    wire N__56109;
    wire N__56106;
    wire N__56103;
    wire N__56102;
    wire N__56101;
    wire N__56100;
    wire N__56099;
    wire N__56098;
    wire N__56097;
    wire N__56096;
    wire N__56095;
    wire N__56094;
    wire N__56093;
    wire N__56092;
    wire N__56091;
    wire N__56090;
    wire N__56089;
    wire N__56088;
    wire N__56087;
    wire N__56086;
    wire N__56085;
    wire N__56084;
    wire N__56083;
    wire N__56082;
    wire N__56081;
    wire N__56080;
    wire N__56079;
    wire N__56078;
    wire N__56077;
    wire N__56076;
    wire N__56075;
    wire N__56074;
    wire N__56073;
    wire N__56072;
    wire N__56071;
    wire N__56070;
    wire N__56069;
    wire N__56068;
    wire N__56067;
    wire N__56066;
    wire N__56065;
    wire N__56064;
    wire N__56063;
    wire N__56062;
    wire N__56061;
    wire N__56060;
    wire N__56059;
    wire N__56058;
    wire N__56057;
    wire N__56056;
    wire N__56055;
    wire N__56054;
    wire N__56053;
    wire N__56052;
    wire N__56051;
    wire N__56050;
    wire N__56049;
    wire N__56048;
    wire N__56047;
    wire N__56046;
    wire N__56045;
    wire N__56044;
    wire N__56043;
    wire N__56042;
    wire N__56041;
    wire N__56040;
    wire N__56039;
    wire N__56038;
    wire N__56037;
    wire N__56036;
    wire N__56035;
    wire N__56034;
    wire N__56033;
    wire N__56032;
    wire N__56031;
    wire N__56030;
    wire N__56029;
    wire N__56028;
    wire N__56027;
    wire N__56026;
    wire N__56025;
    wire N__56024;
    wire N__56023;
    wire N__56022;
    wire N__56021;
    wire N__56020;
    wire N__56019;
    wire N__56018;
    wire N__56017;
    wire N__56016;
    wire N__56015;
    wire N__56014;
    wire N__56013;
    wire N__56012;
    wire N__56011;
    wire N__56010;
    wire N__56009;
    wire N__56008;
    wire N__56007;
    wire N__56006;
    wire N__56005;
    wire N__56004;
    wire N__56003;
    wire N__56002;
    wire N__56001;
    wire N__56000;
    wire N__55999;
    wire N__55998;
    wire N__55997;
    wire N__55996;
    wire N__55995;
    wire N__55994;
    wire N__55993;
    wire N__55992;
    wire N__55991;
    wire N__55990;
    wire N__55989;
    wire N__55988;
    wire N__55987;
    wire N__55986;
    wire N__55985;
    wire N__55984;
    wire N__55983;
    wire N__55982;
    wire N__55981;
    wire N__55980;
    wire N__55979;
    wire N__55978;
    wire N__55977;
    wire N__55976;
    wire N__55975;
    wire N__55974;
    wire N__55973;
    wire N__55972;
    wire N__55971;
    wire N__55970;
    wire N__55969;
    wire N__55968;
    wire N__55967;
    wire N__55966;
    wire N__55965;
    wire N__55964;
    wire N__55963;
    wire N__55962;
    wire N__55961;
    wire N__55960;
    wire N__55959;
    wire N__55958;
    wire N__55957;
    wire N__55956;
    wire N__55955;
    wire N__55954;
    wire N__55953;
    wire N__55952;
    wire N__55951;
    wire N__55950;
    wire N__55949;
    wire N__55948;
    wire N__55947;
    wire N__55946;
    wire N__55945;
    wire N__55944;
    wire N__55943;
    wire N__55942;
    wire N__55941;
    wire N__55940;
    wire N__55939;
    wire N__55938;
    wire N__55937;
    wire N__55602;
    wire N__55599;
    wire N__55596;
    wire N__55593;
    wire N__55590;
    wire N__55587;
    wire N__55584;
    wire N__55581;
    wire N__55578;
    wire N__55575;
    wire N__55574;
    wire N__55573;
    wire N__55572;
    wire N__55571;
    wire N__55568;
    wire N__55565;
    wire N__55564;
    wire N__55563;
    wire N__55562;
    wire N__55559;
    wire N__55554;
    wire N__55553;
    wire N__55548;
    wire N__55545;
    wire N__55544;
    wire N__55541;
    wire N__55538;
    wire N__55537;
    wire N__55536;
    wire N__55533;
    wire N__55530;
    wire N__55527;
    wire N__55524;
    wire N__55521;
    wire N__55518;
    wire N__55513;
    wire N__55508;
    wire N__55503;
    wire N__55496;
    wire N__55489;
    wire N__55482;
    wire N__55479;
    wire N__55478;
    wire N__55475;
    wire N__55474;
    wire N__55473;
    wire N__55472;
    wire N__55471;
    wire N__55470;
    wire N__55469;
    wire N__55468;
    wire N__55467;
    wire N__55466;
    wire N__55465;
    wire N__55464;
    wire N__55463;
    wire N__55462;
    wire N__55461;
    wire N__55460;
    wire N__55459;
    wire N__55456;
    wire N__55455;
    wire N__55452;
    wire N__55441;
    wire N__55440;
    wire N__55439;
    wire N__55438;
    wire N__55437;
    wire N__55436;
    wire N__55435;
    wire N__55434;
    wire N__55433;
    wire N__55432;
    wire N__55431;
    wire N__55430;
    wire N__55429;
    wire N__55428;
    wire N__55427;
    wire N__55424;
    wire N__55423;
    wire N__55422;
    wire N__55421;
    wire N__55420;
    wire N__55419;
    wire N__55418;
    wire N__55415;
    wire N__55414;
    wire N__55411;
    wire N__55410;
    wire N__55407;
    wire N__55406;
    wire N__55403;
    wire N__55402;
    wire N__55399;
    wire N__55396;
    wire N__55389;
    wire N__55388;
    wire N__55387;
    wire N__55384;
    wire N__55381;
    wire N__55378;
    wire N__55373;
    wire N__55368;
    wire N__55359;
    wire N__55358;
    wire N__55355;
    wire N__55352;
    wire N__55347;
    wire N__55346;
    wire N__55343;
    wire N__55336;
    wire N__55325;
    wire N__55322;
    wire N__55319;
    wire N__55302;
    wire N__55299;
    wire N__55298;
    wire N__55297;
    wire N__55296;
    wire N__55295;
    wire N__55294;
    wire N__55293;
    wire N__55292;
    wire N__55289;
    wire N__55288;
    wire N__55287;
    wire N__55286;
    wire N__55285;
    wire N__55282;
    wire N__55281;
    wire N__55280;
    wire N__55279;
    wire N__55276;
    wire N__55273;
    wire N__55272;
    wire N__55271;
    wire N__55270;
    wire N__55269;
    wire N__55268;
    wire N__55255;
    wire N__55252;
    wire N__55251;
    wire N__55250;
    wire N__55249;
    wire N__55248;
    wire N__55247;
    wire N__55244;
    wire N__55239;
    wire N__55238;
    wire N__55237;
    wire N__55236;
    wire N__55235;
    wire N__55234;
    wire N__55233;
    wire N__55230;
    wire N__55227;
    wire N__55216;
    wire N__55213;
    wire N__55208;
    wire N__55207;
    wire N__55204;
    wire N__55195;
    wire N__55192;
    wire N__55187;
    wire N__55184;
    wire N__55183;
    wire N__55182;
    wire N__55181;
    wire N__55180;
    wire N__55177;
    wire N__55174;
    wire N__55171;
    wire N__55166;
    wire N__55165;
    wire N__55164;
    wire N__55163;
    wire N__55160;
    wire N__55157;
    wire N__55154;
    wire N__55149;
    wire N__55144;
    wire N__55141;
    wire N__55136;
    wire N__55131;
    wire N__55126;
    wire N__55121;
    wire N__55120;
    wire N__55109;
    wire N__55108;
    wire N__55105;
    wire N__55104;
    wire N__55101;
    wire N__55096;
    wire N__55091;
    wire N__55088;
    wire N__55085;
    wire N__55076;
    wire N__55069;
    wire N__55068;
    wire N__55067;
    wire N__55066;
    wire N__55065;
    wire N__55062;
    wire N__55059;
    wire N__55056;
    wire N__55051;
    wire N__55044;
    wire N__55033;
    wire N__55030;
    wire N__55029;
    wire N__55028;
    wire N__55027;
    wire N__55024;
    wire N__55017;
    wire N__55014;
    wire N__55011;
    wire N__55008;
    wire N__55005;
    wire N__55002;
    wire N__54995;
    wire N__54990;
    wire N__54985;
    wire N__54980;
    wire N__54977;
    wire N__54974;
    wire N__54965;
    wire N__54958;
    wire N__54951;
    wire N__54946;
    wire N__54941;
    wire N__54934;
    wire N__54931;
    wire N__54924;
    wire N__54903;
    wire N__54900;
    wire N__54897;
    wire N__54894;
    wire N__54893;
    wire N__54892;
    wire N__54891;
    wire N__54888;
    wire N__54887;
    wire N__54886;
    wire N__54885;
    wire N__54884;
    wire N__54881;
    wire N__54876;
    wire N__54875;
    wire N__54874;
    wire N__54871;
    wire N__54864;
    wire N__54863;
    wire N__54862;
    wire N__54861;
    wire N__54860;
    wire N__54859;
    wire N__54858;
    wire N__54857;
    wire N__54854;
    wire N__54853;
    wire N__54852;
    wire N__54851;
    wire N__54848;
    wire N__54847;
    wire N__54844;
    wire N__54843;
    wire N__54842;
    wire N__54841;
    wire N__54840;
    wire N__54839;
    wire N__54836;
    wire N__54833;
    wire N__54828;
    wire N__54827;
    wire N__54826;
    wire N__54825;
    wire N__54822;
    wire N__54811;
    wire N__54810;
    wire N__54807;
    wire N__54804;
    wire N__54803;
    wire N__54800;
    wire N__54797;
    wire N__54796;
    wire N__54795;
    wire N__54792;
    wire N__54789;
    wire N__54788;
    wire N__54787;
    wire N__54784;
    wire N__54781;
    wire N__54778;
    wire N__54777;
    wire N__54774;
    wire N__54771;
    wire N__54766;
    wire N__54761;
    wire N__54758;
    wire N__54755;
    wire N__54754;
    wire N__54753;
    wire N__54750;
    wire N__54747;
    wire N__54744;
    wire N__54741;
    wire N__54740;
    wire N__54739;
    wire N__54738;
    wire N__54737;
    wire N__54734;
    wire N__54731;
    wire N__54728;
    wire N__54725;
    wire N__54716;
    wire N__54711;
    wire N__54710;
    wire N__54707;
    wire N__54706;
    wire N__54703;
    wire N__54696;
    wire N__54691;
    wire N__54686;
    wire N__54685;
    wire N__54684;
    wire N__54683;
    wire N__54680;
    wire N__54675;
    wire N__54670;
    wire N__54667;
    wire N__54662;
    wire N__54659;
    wire N__54652;
    wire N__54649;
    wire N__54646;
    wire N__54643;
    wire N__54640;
    wire N__54633;
    wire N__54626;
    wire N__54617;
    wire N__54610;
    wire N__54603;
    wire N__54594;
    wire N__54573;
    wire N__54572;
    wire N__54571;
    wire N__54568;
    wire N__54567;
    wire N__54566;
    wire N__54563;
    wire N__54560;
    wire N__54557;
    wire N__54556;
    wire N__54555;
    wire N__54554;
    wire N__54553;
    wire N__54552;
    wire N__54551;
    wire N__54550;
    wire N__54549;
    wire N__54548;
    wire N__54547;
    wire N__54546;
    wire N__54545;
    wire N__54544;
    wire N__54543;
    wire N__54542;
    wire N__54541;
    wire N__54538;
    wire N__54535;
    wire N__54534;
    wire N__54531;
    wire N__54526;
    wire N__54525;
    wire N__54522;
    wire N__54519;
    wire N__54518;
    wire N__54517;
    wire N__54516;
    wire N__54515;
    wire N__54514;
    wire N__54511;
    wire N__54510;
    wire N__54509;
    wire N__54508;
    wire N__54507;
    wire N__54506;
    wire N__54505;
    wire N__54504;
    wire N__54503;
    wire N__54502;
    wire N__54501;
    wire N__54500;
    wire N__54499;
    wire N__54498;
    wire N__54495;
    wire N__54494;
    wire N__54491;
    wire N__54490;
    wire N__54489;
    wire N__54488;
    wire N__54487;
    wire N__54486;
    wire N__54485;
    wire N__54484;
    wire N__54467;
    wire N__54464;
    wire N__54461;
    wire N__54458;
    wire N__54455;
    wire N__54452;
    wire N__54449;
    wire N__54444;
    wire N__54441;
    wire N__54440;
    wire N__54439;
    wire N__54438;
    wire N__54437;
    wire N__54436;
    wire N__54435;
    wire N__54434;
    wire N__54433;
    wire N__54432;
    wire N__54431;
    wire N__54430;
    wire N__54429;
    wire N__54426;
    wire N__54423;
    wire N__54418;
    wire N__54417;
    wire N__54414;
    wire N__54411;
    wire N__54410;
    wire N__54409;
    wire N__54406;
    wire N__54403;
    wire N__54402;
    wire N__54401;
    wire N__54400;
    wire N__54397;
    wire N__54390;
    wire N__54381;
    wire N__54380;
    wire N__54379;
    wire N__54376;
    wire N__54375;
    wire N__54374;
    wire N__54371;
    wire N__54368;
    wire N__54367;
    wire N__54366;
    wire N__54363;
    wire N__54360;
    wire N__54357;
    wire N__54350;
    wire N__54343;
    wire N__54342;
    wire N__54341;
    wire N__54340;
    wire N__54339;
    wire N__54338;
    wire N__54337;
    wire N__54336;
    wire N__54335;
    wire N__54334;
    wire N__54333;
    wire N__54332;
    wire N__54331;
    wire N__54326;
    wire N__54323;
    wire N__54308;
    wire N__54303;
    wire N__54300;
    wire N__54293;
    wire N__54276;
    wire N__54269;
    wire N__54266;
    wire N__54263;
    wire N__54256;
    wire N__54251;
    wire N__54248;
    wire N__54245;
    wire N__54242;
    wire N__54235;
    wire N__54232;
    wire N__54225;
    wire N__54222;
    wire N__54217;
    wire N__54212;
    wire N__54201;
    wire N__54200;
    wire N__54199;
    wire N__54198;
    wire N__54197;
    wire N__54196;
    wire N__54195;
    wire N__54194;
    wire N__54193;
    wire N__54192;
    wire N__54191;
    wire N__54188;
    wire N__54185;
    wire N__54184;
    wire N__54183;
    wire N__54180;
    wire N__54179;
    wire N__54178;
    wire N__54177;
    wire N__54174;
    wire N__54173;
    wire N__54172;
    wire N__54155;
    wire N__54152;
    wire N__54141;
    wire N__54136;
    wire N__54129;
    wire N__54126;
    wire N__54115;
    wire N__54112;
    wire N__54103;
    wire N__54086;
    wire N__54081;
    wire N__54078;
    wire N__54075;
    wire N__54068;
    wire N__54063;
    wire N__54054;
    wire N__54047;
    wire N__54042;
    wire N__54037;
    wire N__54032;
    wire N__54009;
    wire N__54008;
    wire N__54007;
    wire N__54006;
    wire N__54005;
    wire N__54004;
    wire N__54003;
    wire N__54002;
    wire N__54001;
    wire N__53998;
    wire N__53997;
    wire N__53994;
    wire N__53989;
    wire N__53988;
    wire N__53987;
    wire N__53986;
    wire N__53983;
    wire N__53982;
    wire N__53981;
    wire N__53980;
    wire N__53979;
    wire N__53978;
    wire N__53977;
    wire N__53970;
    wire N__53969;
    wire N__53966;
    wire N__53965;
    wire N__53964;
    wire N__53963;
    wire N__53962;
    wire N__53959;
    wire N__53956;
    wire N__53951;
    wire N__53948;
    wire N__53947;
    wire N__53946;
    wire N__53943;
    wire N__53940;
    wire N__53931;
    wire N__53924;
    wire N__53923;
    wire N__53922;
    wire N__53921;
    wire N__53920;
    wire N__53919;
    wire N__53916;
    wire N__53913;
    wire N__53910;
    wire N__53905;
    wire N__53900;
    wire N__53897;
    wire N__53894;
    wire N__53889;
    wire N__53886;
    wire N__53883;
    wire N__53880;
    wire N__53877;
    wire N__53874;
    wire N__53873;
    wire N__53872;
    wire N__53871;
    wire N__53870;
    wire N__53869;
    wire N__53868;
    wire N__53865;
    wire N__53860;
    wire N__53853;
    wire N__53850;
    wire N__53845;
    wire N__53838;
    wire N__53833;
    wire N__53830;
    wire N__53823;
    wire N__53820;
    wire N__53811;
    wire N__53806;
    wire N__53793;
    wire N__53790;
    wire N__53775;
    wire N__53772;
    wire N__53769;
    wire N__53766;
    wire N__53763;
    wire N__53760;
    wire N__53757;
    wire N__53756;
    wire N__53753;
    wire N__53750;
    wire N__53747;
    wire N__53742;
    wire N__53741;
    wire N__53738;
    wire N__53735;
    wire N__53732;
    wire N__53727;
    wire N__53726;
    wire N__53723;
    wire N__53720;
    wire N__53717;
    wire N__53712;
    wire N__53711;
    wire N__53708;
    wire N__53705;
    wire N__53702;
    wire N__53697;
    wire N__53694;
    wire N__53691;
    wire N__53688;
    wire N__53685;
    wire N__53682;
    wire N__53679;
    wire N__53676;
    wire N__53675;
    wire N__53674;
    wire N__53671;
    wire N__53666;
    wire N__53663;
    wire N__53660;
    wire N__53655;
    wire N__53652;
    wire N__53649;
    wire N__53646;
    wire N__53645;
    wire N__53644;
    wire N__53641;
    wire N__53640;
    wire N__53637;
    wire N__53636;
    wire N__53633;
    wire N__53630;
    wire N__53627;
    wire N__53624;
    wire N__53621;
    wire N__53620;
    wire N__53619;
    wire N__53612;
    wire N__53607;
    wire N__53604;
    wire N__53601;
    wire N__53600;
    wire N__53597;
    wire N__53594;
    wire N__53591;
    wire N__53588;
    wire N__53585;
    wire N__53584;
    wire N__53581;
    wire N__53578;
    wire N__53573;
    wire N__53570;
    wire N__53567;
    wire N__53556;
    wire N__53553;
    wire N__53552;
    wire N__53549;
    wire N__53546;
    wire N__53543;
    wire N__53538;
    wire N__53535;
    wire N__53532;
    wire N__53529;
    wire N__53526;
    wire N__53523;
    wire N__53520;
    wire N__53517;
    wire N__53514;
    wire N__53511;
    wire N__53510;
    wire N__53507;
    wire N__53504;
    wire N__53503;
    wire N__53500;
    wire N__53499;
    wire N__53496;
    wire N__53493;
    wire N__53490;
    wire N__53487;
    wire N__53482;
    wire N__53477;
    wire N__53474;
    wire N__53471;
    wire N__53466;
    wire N__53463;
    wire N__53462;
    wire N__53459;
    wire N__53458;
    wire N__53455;
    wire N__53452;
    wire N__53449;
    wire N__53448;
    wire N__53445;
    wire N__53442;
    wire N__53439;
    wire N__53438;
    wire N__53437;
    wire N__53436;
    wire N__53435;
    wire N__53432;
    wire N__53425;
    wire N__53424;
    wire N__53423;
    wire N__53418;
    wire N__53415;
    wire N__53412;
    wire N__53407;
    wire N__53404;
    wire N__53401;
    wire N__53398;
    wire N__53393;
    wire N__53390;
    wire N__53387;
    wire N__53384;
    wire N__53381;
    wire N__53378;
    wire N__53375;
    wire N__53370;
    wire N__53367;
    wire N__53358;
    wire N__53355;
    wire N__53352;
    wire N__53349;
    wire N__53346;
    wire N__53345;
    wire N__53344;
    wire N__53343;
    wire N__53342;
    wire N__53339;
    wire N__53336;
    wire N__53333;
    wire N__53332;
    wire N__53331;
    wire N__53328;
    wire N__53325;
    wire N__53322;
    wire N__53319;
    wire N__53316;
    wire N__53313;
    wire N__53310;
    wire N__53305;
    wire N__53298;
    wire N__53293;
    wire N__53292;
    wire N__53291;
    wire N__53288;
    wire N__53283;
    wire N__53280;
    wire N__53277;
    wire N__53268;
    wire N__53267;
    wire N__53264;
    wire N__53261;
    wire N__53256;
    wire N__53253;
    wire N__53250;
    wire N__53247;
    wire N__53244;
    wire N__53241;
    wire N__53238;
    wire N__53235;
    wire N__53234;
    wire N__53231;
    wire N__53228;
    wire N__53227;
    wire N__53226;
    wire N__53225;
    wire N__53222;
    wire N__53219;
    wire N__53218;
    wire N__53217;
    wire N__53214;
    wire N__53211;
    wire N__53208;
    wire N__53205;
    wire N__53202;
    wire N__53199;
    wire N__53196;
    wire N__53195;
    wire N__53192;
    wire N__53189;
    wire N__53184;
    wire N__53177;
    wire N__53174;
    wire N__53171;
    wire N__53166;
    wire N__53161;
    wire N__53160;
    wire N__53157;
    wire N__53152;
    wire N__53149;
    wire N__53142;
    wire N__53141;
    wire N__53138;
    wire N__53135;
    wire N__53132;
    wire N__53131;
    wire N__53130;
    wire N__53129;
    wire N__53128;
    wire N__53127;
    wire N__53126;
    wire N__53123;
    wire N__53120;
    wire N__53117;
    wire N__53114;
    wire N__53109;
    wire N__53106;
    wire N__53103;
    wire N__53088;
    wire N__53087;
    wire N__53084;
    wire N__53081;
    wire N__53078;
    wire N__53073;
    wire N__53072;
    wire N__53071;
    wire N__53070;
    wire N__53069;
    wire N__53068;
    wire N__53067;
    wire N__53066;
    wire N__53065;
    wire N__53064;
    wire N__53063;
    wire N__53062;
    wire N__53061;
    wire N__53058;
    wire N__53053;
    wire N__53052;
    wire N__53051;
    wire N__53050;
    wire N__53049;
    wire N__53048;
    wire N__53047;
    wire N__53046;
    wire N__53043;
    wire N__53042;
    wire N__53037;
    wire N__53034;
    wire N__53033;
    wire N__53032;
    wire N__53031;
    wire N__53030;
    wire N__53029;
    wire N__53028;
    wire N__53025;
    wire N__53014;
    wire N__53009;
    wire N__53002;
    wire N__52993;
    wire N__52992;
    wire N__52991;
    wire N__52990;
    wire N__52989;
    wire N__52988;
    wire N__52987;
    wire N__52986;
    wire N__52983;
    wire N__52980;
    wire N__52975;
    wire N__52966;
    wire N__52963;
    wire N__52960;
    wire N__52951;
    wire N__52948;
    wire N__52939;
    wire N__52938;
    wire N__52933;
    wire N__52930;
    wire N__52927;
    wire N__52920;
    wire N__52915;
    wire N__52908;
    wire N__52905;
    wire N__52890;
    wire N__52887;
    wire N__52884;
    wire N__52883;
    wire N__52882;
    wire N__52881;
    wire N__52880;
    wire N__52879;
    wire N__52872;
    wire N__52869;
    wire N__52864;
    wire N__52863;
    wire N__52862;
    wire N__52861;
    wire N__52860;
    wire N__52859;
    wire N__52858;
    wire N__52857;
    wire N__52856;
    wire N__52855;
    wire N__52852;
    wire N__52849;
    wire N__52846;
    wire N__52839;
    wire N__52828;
    wire N__52825;
    wire N__52820;
    wire N__52813;
    wire N__52810;
    wire N__52803;
    wire N__52800;
    wire N__52799;
    wire N__52798;
    wire N__52797;
    wire N__52796;
    wire N__52795;
    wire N__52794;
    wire N__52793;
    wire N__52784;
    wire N__52783;
    wire N__52782;
    wire N__52781;
    wire N__52778;
    wire N__52775;
    wire N__52772;
    wire N__52771;
    wire N__52770;
    wire N__52769;
    wire N__52768;
    wire N__52767;
    wire N__52764;
    wire N__52763;
    wire N__52762;
    wire N__52759;
    wire N__52756;
    wire N__52753;
    wire N__52750;
    wire N__52745;
    wire N__52740;
    wire N__52727;
    wire N__52724;
    wire N__52719;
    wire N__52712;
    wire N__52707;
    wire N__52704;
    wire N__52701;
    wire N__52698;
    wire N__52695;
    wire N__52692;
    wire N__52691;
    wire N__52690;
    wire N__52685;
    wire N__52682;
    wire N__52679;
    wire N__52674;
    wire N__52669;
    wire N__52664;
    wire N__52661;
    wire N__52658;
    wire N__52653;
    wire N__52650;
    wire N__52647;
    wire N__52644;
    wire N__52641;
    wire N__52638;
    wire N__52635;
    wire N__52632;
    wire N__52631;
    wire N__52628;
    wire N__52625;
    wire N__52622;
    wire N__52619;
    wire N__52616;
    wire N__52613;
    wire N__52610;
    wire N__52607;
    wire N__52602;
    wire N__52599;
    wire N__52596;
    wire N__52593;
    wire N__52590;
    wire N__52587;
    wire N__52584;
    wire N__52581;
    wire N__52578;
    wire N__52575;
    wire N__52572;
    wire N__52569;
    wire N__52566;
    wire N__52565;
    wire N__52564;
    wire N__52563;
    wire N__52562;
    wire N__52561;
    wire N__52560;
    wire N__52559;
    wire N__52558;
    wire N__52557;
    wire N__52556;
    wire N__52555;
    wire N__52554;
    wire N__52553;
    wire N__52546;
    wire N__52539;
    wire N__52532;
    wire N__52527;
    wire N__52524;
    wire N__52523;
    wire N__52522;
    wire N__52521;
    wire N__52520;
    wire N__52517;
    wire N__52514;
    wire N__52513;
    wire N__52512;
    wire N__52503;
    wire N__52500;
    wire N__52495;
    wire N__52490;
    wire N__52487;
    wire N__52484;
    wire N__52481;
    wire N__52478;
    wire N__52475;
    wire N__52468;
    wire N__52463;
    wire N__52460;
    wire N__52449;
    wire N__52448;
    wire N__52447;
    wire N__52446;
    wire N__52445;
    wire N__52444;
    wire N__52443;
    wire N__52440;
    wire N__52439;
    wire N__52438;
    wire N__52437;
    wire N__52436;
    wire N__52435;
    wire N__52434;
    wire N__52433;
    wire N__52432;
    wire N__52429;
    wire N__52426;
    wire N__52423;
    wire N__52420;
    wire N__52415;
    wire N__52412;
    wire N__52411;
    wire N__52410;
    wire N__52409;
    wire N__52406;
    wire N__52401;
    wire N__52396;
    wire N__52395;
    wire N__52394;
    wire N__52393;
    wire N__52392;
    wire N__52383;
    wire N__52382;
    wire N__52381;
    wire N__52380;
    wire N__52379;
    wire N__52378;
    wire N__52377;
    wire N__52376;
    wire N__52371;
    wire N__52364;
    wire N__52355;
    wire N__52350;
    wire N__52345;
    wire N__52340;
    wire N__52337;
    wire N__52334;
    wire N__52325;
    wire N__52320;
    wire N__52313;
    wire N__52304;
    wire N__52299;
    wire N__52290;
    wire N__52287;
    wire N__52286;
    wire N__52285;
    wire N__52282;
    wire N__52279;
    wire N__52278;
    wire N__52277;
    wire N__52276;
    wire N__52275;
    wire N__52272;
    wire N__52269;
    wire N__52266;
    wire N__52263;
    wire N__52260;
    wire N__52257;
    wire N__52254;
    wire N__52251;
    wire N__52246;
    wire N__52243;
    wire N__52240;
    wire N__52237;
    wire N__52234;
    wire N__52231;
    wire N__52228;
    wire N__52225;
    wire N__52220;
    wire N__52217;
    wire N__52214;
    wire N__52209;
    wire N__52200;
    wire N__52197;
    wire N__52194;
    wire N__52191;
    wire N__52188;
    wire N__52185;
    wire N__52182;
    wire N__52179;
    wire N__52176;
    wire N__52173;
    wire N__52170;
    wire N__52169;
    wire N__52166;
    wire N__52163;
    wire N__52160;
    wire N__52157;
    wire N__52152;
    wire N__52151;
    wire N__52150;
    wire N__52147;
    wire N__52144;
    wire N__52141;
    wire N__52138;
    wire N__52135;
    wire N__52132;
    wire N__52129;
    wire N__52122;
    wire N__52119;
    wire N__52116;
    wire N__52113;
    wire N__52110;
    wire N__52107;
    wire N__52104;
    wire N__52101;
    wire N__52098;
    wire N__52095;
    wire N__52094;
    wire N__52091;
    wire N__52090;
    wire N__52087;
    wire N__52084;
    wire N__52081;
    wire N__52078;
    wire N__52075;
    wire N__52072;
    wire N__52069;
    wire N__52064;
    wire N__52059;
    wire N__52056;
    wire N__52055;
    wire N__52052;
    wire N__52049;
    wire N__52044;
    wire N__52041;
    wire N__52038;
    wire N__52035;
    wire N__52032;
    wire N__52029;
    wire N__52026;
    wire N__52023;
    wire N__52020;
    wire N__52017;
    wire N__52014;
    wire N__52011;
    wire N__52008;
    wire N__52005;
    wire N__52004;
    wire N__52001;
    wire N__52000;
    wire N__51997;
    wire N__51994;
    wire N__51993;
    wire N__51990;
    wire N__51987;
    wire N__51986;
    wire N__51985;
    wire N__51982;
    wire N__51979;
    wire N__51976;
    wire N__51975;
    wire N__51974;
    wire N__51971;
    wire N__51966;
    wire N__51959;
    wire N__51954;
    wire N__51951;
    wire N__51948;
    wire N__51943;
    wire N__51942;
    wire N__51939;
    wire N__51934;
    wire N__51931;
    wire N__51928;
    wire N__51923;
    wire N__51918;
    wire N__51915;
    wire N__51912;
    wire N__51911;
    wire N__51910;
    wire N__51909;
    wire N__51908;
    wire N__51905;
    wire N__51904;
    wire N__51903;
    wire N__51900;
    wire N__51897;
    wire N__51896;
    wire N__51895;
    wire N__51894;
    wire N__51893;
    wire N__51892;
    wire N__51889;
    wire N__51886;
    wire N__51883;
    wire N__51882;
    wire N__51881;
    wire N__51880;
    wire N__51877;
    wire N__51874;
    wire N__51871;
    wire N__51868;
    wire N__51867;
    wire N__51864;
    wire N__51861;
    wire N__51860;
    wire N__51859;
    wire N__51858;
    wire N__51857;
    wire N__51856;
    wire N__51853;
    wire N__51846;
    wire N__51843;
    wire N__51840;
    wire N__51833;
    wire N__51828;
    wire N__51823;
    wire N__51820;
    wire N__51817;
    wire N__51814;
    wire N__51811;
    wire N__51806;
    wire N__51803;
    wire N__51800;
    wire N__51789;
    wire N__51786;
    wire N__51783;
    wire N__51762;
    wire N__51761;
    wire N__51760;
    wire N__51759;
    wire N__51758;
    wire N__51755;
    wire N__51754;
    wire N__51753;
    wire N__51750;
    wire N__51747;
    wire N__51746;
    wire N__51745;
    wire N__51744;
    wire N__51741;
    wire N__51738;
    wire N__51735;
    wire N__51732;
    wire N__51729;
    wire N__51726;
    wire N__51723;
    wire N__51722;
    wire N__51721;
    wire N__51720;
    wire N__51717;
    wire N__51714;
    wire N__51713;
    wire N__51712;
    wire N__51711;
    wire N__51710;
    wire N__51709;
    wire N__51708;
    wire N__51707;
    wire N__51706;
    wire N__51705;
    wire N__51704;
    wire N__51703;
    wire N__51702;
    wire N__51701;
    wire N__51700;
    wire N__51699;
    wire N__51698;
    wire N__51697;
    wire N__51696;
    wire N__51691;
    wire N__51690;
    wire N__51687;
    wire N__51684;
    wire N__51681;
    wire N__51674;
    wire N__51669;
    wire N__51666;
    wire N__51661;
    wire N__51652;
    wire N__51649;
    wire N__51648;
    wire N__51645;
    wire N__51642;
    wire N__51641;
    wire N__51640;
    wire N__51639;
    wire N__51638;
    wire N__51637;
    wire N__51636;
    wire N__51635;
    wire N__51634;
    wire N__51625;
    wire N__51616;
    wire N__51609;
    wire N__51606;
    wire N__51603;
    wire N__51602;
    wire N__51601;
    wire N__51600;
    wire N__51599;
    wire N__51596;
    wire N__51593;
    wire N__51590;
    wire N__51587;
    wire N__51578;
    wire N__51575;
    wire N__51560;
    wire N__51557;
    wire N__51550;
    wire N__51539;
    wire N__51530;
    wire N__51521;
    wire N__51518;
    wire N__51501;
    wire N__51500;
    wire N__51499;
    wire N__51498;
    wire N__51497;
    wire N__51496;
    wire N__51495;
    wire N__51494;
    wire N__51493;
    wire N__51492;
    wire N__51491;
    wire N__51490;
    wire N__51489;
    wire N__51488;
    wire N__51485;
    wire N__51484;
    wire N__51483;
    wire N__51482;
    wire N__51481;
    wire N__51480;
    wire N__51479;
    wire N__51478;
    wire N__51477;
    wire N__51476;
    wire N__51475;
    wire N__51474;
    wire N__51473;
    wire N__51470;
    wire N__51457;
    wire N__51456;
    wire N__51455;
    wire N__51452;
    wire N__51449;
    wire N__51446;
    wire N__51443;
    wire N__51442;
    wire N__51437;
    wire N__51424;
    wire N__51421;
    wire N__51416;
    wire N__51415;
    wire N__51414;
    wire N__51413;
    wire N__51412;
    wire N__51409;
    wire N__51402;
    wire N__51399;
    wire N__51396;
    wire N__51391;
    wire N__51386;
    wire N__51385;
    wire N__51380;
    wire N__51377;
    wire N__51374;
    wire N__51371;
    wire N__51368;
    wire N__51365;
    wire N__51364;
    wire N__51363;
    wire N__51362;
    wire N__51361;
    wire N__51358;
    wire N__51357;
    wire N__51356;
    wire N__51355;
    wire N__51352;
    wire N__51349;
    wire N__51346;
    wire N__51345;
    wire N__51344;
    wire N__51339;
    wire N__51332;
    wire N__51331;
    wire N__51330;
    wire N__51329;
    wire N__51328;
    wire N__51327;
    wire N__51324;
    wire N__51321;
    wire N__51312;
    wire N__51309;
    wire N__51306;
    wire N__51295;
    wire N__51286;
    wire N__51281;
    wire N__51278;
    wire N__51275;
    wire N__51272;
    wire N__51269;
    wire N__51264;
    wire N__51257;
    wire N__51254;
    wire N__51251;
    wire N__51246;
    wire N__51237;
    wire N__51216;
    wire N__51213;
    wire N__51212;
    wire N__51211;
    wire N__51210;
    wire N__51209;
    wire N__51208;
    wire N__51205;
    wire N__51204;
    wire N__51203;
    wire N__51198;
    wire N__51197;
    wire N__51194;
    wire N__51191;
    wire N__51188;
    wire N__51185;
    wire N__51184;
    wire N__51181;
    wire N__51180;
    wire N__51179;
    wire N__51176;
    wire N__51175;
    wire N__51174;
    wire N__51171;
    wire N__51168;
    wire N__51163;
    wire N__51158;
    wire N__51155;
    wire N__51154;
    wire N__51153;
    wire N__51152;
    wire N__51151;
    wire N__51150;
    wire N__51149;
    wire N__51146;
    wire N__51145;
    wire N__51142;
    wire N__51139;
    wire N__51136;
    wire N__51133;
    wire N__51130;
    wire N__51125;
    wire N__51118;
    wire N__51111;
    wire N__51104;
    wire N__51101;
    wire N__51098;
    wire N__51075;
    wire N__51072;
    wire N__51069;
    wire N__51066;
    wire N__51063;
    wire N__51060;
    wire N__51057;
    wire N__51054;
    wire N__51051;
    wire N__51048;
    wire N__51045;
    wire N__51044;
    wire N__51041;
    wire N__51038;
    wire N__51033;
    wire N__51030;
    wire N__51027;
    wire N__51024;
    wire N__51021;
    wire N__51020;
    wire N__51015;
    wire N__51012;
    wire N__51009;
    wire N__51006;
    wire N__51005;
    wire N__51002;
    wire N__50999;
    wire N__50994;
    wire N__50991;
    wire N__50990;
    wire N__50987;
    wire N__50984;
    wire N__50983;
    wire N__50982;
    wire N__50981;
    wire N__50980;
    wire N__50977;
    wire N__50972;
    wire N__50969;
    wire N__50966;
    wire N__50963;
    wire N__50960;
    wire N__50957;
    wire N__50954;
    wire N__50953;
    wire N__50952;
    wire N__50949;
    wire N__50946;
    wire N__50941;
    wire N__50938;
    wire N__50933;
    wire N__50928;
    wire N__50925;
    wire N__50922;
    wire N__50919;
    wire N__50916;
    wire N__50913;
    wire N__50908;
    wire N__50905;
    wire N__50902;
    wire N__50899;
    wire N__50892;
    wire N__50891;
    wire N__50888;
    wire N__50885;
    wire N__50884;
    wire N__50879;
    wire N__50876;
    wire N__50875;
    wire N__50870;
    wire N__50869;
    wire N__50866;
    wire N__50863;
    wire N__50860;
    wire N__50857;
    wire N__50852;
    wire N__50849;
    wire N__50846;
    wire N__50843;
    wire N__50840;
    wire N__50837;
    wire N__50832;
    wire N__50829;
    wire N__50826;
    wire N__50823;
    wire N__50820;
    wire N__50817;
    wire N__50814;
    wire N__50811;
    wire N__50810;
    wire N__50807;
    wire N__50804;
    wire N__50803;
    wire N__50800;
    wire N__50799;
    wire N__50798;
    wire N__50797;
    wire N__50796;
    wire N__50795;
    wire N__50794;
    wire N__50793;
    wire N__50792;
    wire N__50791;
    wire N__50790;
    wire N__50789;
    wire N__50788;
    wire N__50787;
    wire N__50786;
    wire N__50785;
    wire N__50784;
    wire N__50783;
    wire N__50782;
    wire N__50781;
    wire N__50778;
    wire N__50733;
    wire N__50730;
    wire N__50729;
    wire N__50724;
    wire N__50721;
    wire N__50720;
    wire N__50717;
    wire N__50714;
    wire N__50711;
    wire N__50710;
    wire N__50707;
    wire N__50704;
    wire N__50701;
    wire N__50698;
    wire N__50691;
    wire N__50688;
    wire N__50685;
    wire N__50682;
    wire N__50679;
    wire N__50676;
    wire N__50673;
    wire N__50670;
    wire N__50667;
    wire N__50664;
    wire N__50663;
    wire N__50660;
    wire N__50657;
    wire N__50654;
    wire N__50649;
    wire N__50648;
    wire N__50645;
    wire N__50644;
    wire N__50641;
    wire N__50638;
    wire N__50635;
    wire N__50628;
    wire N__50625;
    wire N__50622;
    wire N__50621;
    wire N__50618;
    wire N__50615;
    wire N__50612;
    wire N__50607;
    wire N__50606;
    wire N__50605;
    wire N__50600;
    wire N__50597;
    wire N__50592;
    wire N__50589;
    wire N__50586;
    wire N__50583;
    wire N__50580;
    wire N__50577;
    wire N__50574;
    wire N__50571;
    wire N__50568;
    wire N__50567;
    wire N__50564;
    wire N__50561;
    wire N__50556;
    wire N__50553;
    wire N__50552;
    wire N__50549;
    wire N__50546;
    wire N__50543;
    wire N__50538;
    wire N__50535;
    wire N__50534;
    wire N__50531;
    wire N__50528;
    wire N__50525;
    wire N__50520;
    wire N__50517;
    wire N__50516;
    wire N__50513;
    wire N__50510;
    wire N__50505;
    wire N__50502;
    wire N__50501;
    wire N__50498;
    wire N__50495;
    wire N__50490;
    wire N__50487;
    wire N__50484;
    wire N__50481;
    wire N__50478;
    wire N__50475;
    wire N__50472;
    wire N__50469;
    wire N__50466;
    wire N__50463;
    wire N__50462;
    wire N__50459;
    wire N__50456;
    wire N__50455;
    wire N__50450;
    wire N__50447;
    wire N__50442;
    wire N__50439;
    wire N__50436;
    wire N__50433;
    wire N__50430;
    wire N__50427;
    wire N__50424;
    wire N__50423;
    wire N__50422;
    wire N__50419;
    wire N__50418;
    wire N__50415;
    wire N__50414;
    wire N__50411;
    wire N__50406;
    wire N__50403;
    wire N__50400;
    wire N__50397;
    wire N__50394;
    wire N__50391;
    wire N__50388;
    wire N__50385;
    wire N__50382;
    wire N__50375;
    wire N__50370;
    wire N__50367;
    wire N__50364;
    wire N__50361;
    wire N__50358;
    wire N__50355;
    wire N__50354;
    wire N__50351;
    wire N__50348;
    wire N__50343;
    wire N__50342;
    wire N__50341;
    wire N__50338;
    wire N__50335;
    wire N__50334;
    wire N__50333;
    wire N__50330;
    wire N__50325;
    wire N__50322;
    wire N__50321;
    wire N__50318;
    wire N__50315;
    wire N__50312;
    wire N__50309;
    wire N__50306;
    wire N__50305;
    wire N__50302;
    wire N__50299;
    wire N__50296;
    wire N__50291;
    wire N__50288;
    wire N__50285;
    wire N__50282;
    wire N__50279;
    wire N__50276;
    wire N__50265;
    wire N__50262;
    wire N__50261;
    wire N__50258;
    wire N__50255;
    wire N__50254;
    wire N__50251;
    wire N__50250;
    wire N__50247;
    wire N__50244;
    wire N__50243;
    wire N__50240;
    wire N__50237;
    wire N__50232;
    wire N__50231;
    wire N__50228;
    wire N__50227;
    wire N__50224;
    wire N__50219;
    wire N__50216;
    wire N__50213;
    wire N__50210;
    wire N__50207;
    wire N__50204;
    wire N__50201;
    wire N__50198;
    wire N__50191;
    wire N__50184;
    wire N__50181;
    wire N__50178;
    wire N__50175;
    wire N__50172;
    wire N__50169;
    wire N__50166;
    wire N__50165;
    wire N__50162;
    wire N__50159;
    wire N__50158;
    wire N__50157;
    wire N__50156;
    wire N__50153;
    wire N__50150;
    wire N__50147;
    wire N__50146;
    wire N__50145;
    wire N__50142;
    wire N__50139;
    wire N__50136;
    wire N__50131;
    wire N__50128;
    wire N__50125;
    wire N__50122;
    wire N__50119;
    wire N__50114;
    wire N__50109;
    wire N__50108;
    wire N__50105;
    wire N__50098;
    wire N__50095;
    wire N__50094;
    wire N__50091;
    wire N__50088;
    wire N__50085;
    wire N__50082;
    wire N__50073;
    wire N__50072;
    wire N__50069;
    wire N__50066;
    wire N__50061;
    wire N__50058;
    wire N__50055;
    wire N__50052;
    wire N__50049;
    wire N__50046;
    wire N__50043;
    wire N__50040;
    wire N__50037;
    wire N__50034;
    wire N__50031;
    wire N__50028;
    wire N__50025;
    wire N__50022;
    wire N__50019;
    wire N__50016;
    wire N__50013;
    wire N__50010;
    wire N__50007;
    wire N__50004;
    wire N__50003;
    wire N__50002;
    wire N__49999;
    wire N__49994;
    wire N__49993;
    wire N__49988;
    wire N__49985;
    wire N__49982;
    wire N__49977;
    wire N__49974;
    wire N__49973;
    wire N__49970;
    wire N__49967;
    wire N__49964;
    wire N__49959;
    wire N__49956;
    wire N__49953;
    wire N__49950;
    wire N__49947;
    wire N__49944;
    wire N__49943;
    wire N__49942;
    wire N__49939;
    wire N__49936;
    wire N__49933;
    wire N__49932;
    wire N__49931;
    wire N__49928;
    wire N__49923;
    wire N__49920;
    wire N__49917;
    wire N__49908;
    wire N__49905;
    wire N__49902;
    wire N__49899;
    wire N__49896;
    wire N__49893;
    wire N__49890;
    wire N__49887;
    wire N__49884;
    wire N__49881;
    wire N__49878;
    wire N__49877;
    wire N__49876;
    wire N__49875;
    wire N__49872;
    wire N__49869;
    wire N__49868;
    wire N__49867;
    wire N__49864;
    wire N__49861;
    wire N__49860;
    wire N__49857;
    wire N__49856;
    wire N__49853;
    wire N__49850;
    wire N__49847;
    wire N__49844;
    wire N__49841;
    wire N__49838;
    wire N__49835;
    wire N__49832;
    wire N__49827;
    wire N__49824;
    wire N__49821;
    wire N__49816;
    wire N__49811;
    wire N__49810;
    wire N__49805;
    wire N__49798;
    wire N__49795;
    wire N__49788;
    wire N__49785;
    wire N__49782;
    wire N__49779;
    wire N__49776;
    wire N__49773;
    wire N__49770;
    wire N__49767;
    wire N__49764;
    wire N__49761;
    wire N__49758;
    wire N__49755;
    wire N__49752;
    wire N__49749;
    wire N__49746;
    wire N__49745;
    wire N__49742;
    wire N__49739;
    wire N__49736;
    wire N__49733;
    wire N__49730;
    wire N__49727;
    wire N__49724;
    wire N__49723;
    wire N__49722;
    wire N__49721;
    wire N__49718;
    wire N__49717;
    wire N__49714;
    wire N__49711;
    wire N__49708;
    wire N__49705;
    wire N__49704;
    wire N__49701;
    wire N__49698;
    wire N__49693;
    wire N__49690;
    wire N__49687;
    wire N__49684;
    wire N__49679;
    wire N__49678;
    wire N__49675;
    wire N__49672;
    wire N__49669;
    wire N__49666;
    wire N__49663;
    wire N__49660;
    wire N__49659;
    wire N__49656;
    wire N__49649;
    wire N__49644;
    wire N__49641;
    wire N__49632;
    wire N__49629;
    wire N__49626;
    wire N__49623;
    wire N__49620;
    wire N__49617;
    wire N__49614;
    wire N__49611;
    wire N__49608;
    wire N__49605;
    wire N__49602;
    wire N__49599;
    wire N__49596;
    wire N__49593;
    wire N__49590;
    wire N__49587;
    wire N__49586;
    wire N__49585;
    wire N__49582;
    wire N__49579;
    wire N__49576;
    wire N__49573;
    wire N__49570;
    wire N__49569;
    wire N__49568;
    wire N__49567;
    wire N__49564;
    wire N__49561;
    wire N__49558;
    wire N__49557;
    wire N__49554;
    wire N__49549;
    wire N__49546;
    wire N__49541;
    wire N__49538;
    wire N__49537;
    wire N__49534;
    wire N__49531;
    wire N__49524;
    wire N__49521;
    wire N__49518;
    wire N__49515;
    wire N__49512;
    wire N__49505;
    wire N__49500;
    wire N__49497;
    wire N__49496;
    wire N__49495;
    wire N__49494;
    wire N__49491;
    wire N__49488;
    wire N__49487;
    wire N__49486;
    wire N__49483;
    wire N__49480;
    wire N__49477;
    wire N__49474;
    wire N__49471;
    wire N__49468;
    wire N__49465;
    wire N__49462;
    wire N__49459;
    wire N__49456;
    wire N__49453;
    wire N__49450;
    wire N__49445;
    wire N__49440;
    wire N__49433;
    wire N__49428;
    wire N__49425;
    wire N__49424;
    wire N__49421;
    wire N__49418;
    wire N__49413;
    wire N__49410;
    wire N__49407;
    wire N__49404;
    wire N__49401;
    wire N__49398;
    wire N__49395;
    wire N__49392;
    wire N__49391;
    wire N__49390;
    wire N__49389;
    wire N__49388;
    wire N__49387;
    wire N__49386;
    wire N__49385;
    wire N__49384;
    wire N__49383;
    wire N__49382;
    wire N__49379;
    wire N__49378;
    wire N__49377;
    wire N__49376;
    wire N__49375;
    wire N__49374;
    wire N__49371;
    wire N__49370;
    wire N__49369;
    wire N__49366;
    wire N__49365;
    wire N__49362;
    wire N__49361;
    wire N__49356;
    wire N__49355;
    wire N__49352;
    wire N__49351;
    wire N__49350;
    wire N__49347;
    wire N__49342;
    wire N__49341;
    wire N__49338;
    wire N__49337;
    wire N__49336;
    wire N__49335;
    wire N__49332;
    wire N__49331;
    wire N__49326;
    wire N__49325;
    wire N__49324;
    wire N__49323;
    wire N__49322;
    wire N__49319;
    wire N__49318;
    wire N__49317;
    wire N__49316;
    wire N__49313;
    wire N__49312;
    wire N__49311;
    wire N__49310;
    wire N__49309;
    wire N__49306;
    wire N__49305;
    wire N__49304;
    wire N__49303;
    wire N__49302;
    wire N__49301;
    wire N__49298;
    wire N__49297;
    wire N__49294;
    wire N__49291;
    wire N__49284;
    wire N__49281;
    wire N__49280;
    wire N__49279;
    wire N__49276;
    wire N__49273;
    wire N__49272;
    wire N__49269;
    wire N__49264;
    wire N__49259;
    wire N__49258;
    wire N__49255;
    wire N__49252;
    wire N__49249;
    wire N__49244;
    wire N__49243;
    wire N__49242;
    wire N__49239;
    wire N__49236;
    wire N__49235;
    wire N__49234;
    wire N__49231;
    wire N__49224;
    wire N__49221;
    wire N__49216;
    wire N__49215;
    wire N__49214;
    wire N__49211;
    wire N__49210;
    wire N__49209;
    wire N__49208;
    wire N__49207;
    wire N__49204;
    wire N__49203;
    wire N__49200;
    wire N__49197;
    wire N__49194;
    wire N__49191;
    wire N__49188;
    wire N__49185;
    wire N__49180;
    wire N__49173;
    wire N__49170;
    wire N__49167;
    wire N__49164;
    wire N__49159;
    wire N__49156;
    wire N__49151;
    wire N__49148;
    wire N__49143;
    wire N__49140;
    wire N__49135;
    wire N__49134;
    wire N__49133;
    wire N__49132;
    wire N__49131;
    wire N__49128;
    wire N__49127;
    wire N__49126;
    wire N__49125;
    wire N__49124;
    wire N__49123;
    wire N__49120;
    wire N__49113;
    wire N__49112;
    wire N__49109;
    wire N__49108;
    wire N__49105;
    wire N__49104;
    wire N__49103;
    wire N__49100;
    wire N__49093;
    wire N__49088;
    wire N__49083;
    wire N__49070;
    wire N__49063;
    wire N__49062;
    wire N__49061;
    wire N__49060;
    wire N__49059;
    wire N__49056;
    wire N__49053;
    wire N__49050;
    wire N__49043;
    wire N__49030;
    wire N__49021;
    wire N__49016;
    wire N__49013;
    wire N__49008;
    wire N__48999;
    wire N__48992;
    wire N__48987;
    wire N__48984;
    wire N__48973;
    wire N__48966;
    wire N__48959;
    wire N__48956;
    wire N__48949;
    wire N__48946;
    wire N__48943;
    wire N__48936;
    wire N__48931;
    wire N__48926;
    wire N__48913;
    wire N__48910;
    wire N__48891;
    wire N__48888;
    wire N__48885;
    wire N__48882;
    wire N__48879;
    wire N__48876;
    wire N__48873;
    wire N__48870;
    wire N__48867;
    wire N__48864;
    wire N__48861;
    wire N__48858;
    wire N__48855;
    wire N__48852;
    wire N__48851;
    wire N__48848;
    wire N__48847;
    wire N__48844;
    wire N__48841;
    wire N__48838;
    wire N__48831;
    wire N__48828;
    wire N__48825;
    wire N__48822;
    wire N__48821;
    wire N__48820;
    wire N__48817;
    wire N__48812;
    wire N__48807;
    wire N__48804;
    wire N__48801;
    wire N__48798;
    wire N__48795;
    wire N__48792;
    wire N__48791;
    wire N__48788;
    wire N__48785;
    wire N__48782;
    wire N__48779;
    wire N__48776;
    wire N__48773;
    wire N__48768;
    wire N__48765;
    wire N__48764;
    wire N__48763;
    wire N__48758;
    wire N__48755;
    wire N__48750;
    wire N__48749;
    wire N__48746;
    wire N__48743;
    wire N__48742;
    wire N__48741;
    wire N__48738;
    wire N__48735;
    wire N__48732;
    wire N__48729;
    wire N__48720;
    wire N__48717;
    wire N__48714;
    wire N__48711;
    wire N__48708;
    wire N__48707;
    wire N__48704;
    wire N__48703;
    wire N__48700;
    wire N__48699;
    wire N__48698;
    wire N__48697;
    wire N__48696;
    wire N__48693;
    wire N__48690;
    wire N__48687;
    wire N__48684;
    wire N__48681;
    wire N__48678;
    wire N__48677;
    wire N__48676;
    wire N__48673;
    wire N__48668;
    wire N__48659;
    wire N__48656;
    wire N__48653;
    wire N__48650;
    wire N__48645;
    wire N__48640;
    wire N__48635;
    wire N__48632;
    wire N__48629;
    wire N__48624;
    wire N__48621;
    wire N__48618;
    wire N__48615;
    wire N__48612;
    wire N__48609;
    wire N__48606;
    wire N__48603;
    wire N__48600;
    wire N__48599;
    wire N__48598;
    wire N__48597;
    wire N__48596;
    wire N__48595;
    wire N__48592;
    wire N__48589;
    wire N__48588;
    wire N__48585;
    wire N__48582;
    wire N__48579;
    wire N__48576;
    wire N__48573;
    wire N__48572;
    wire N__48569;
    wire N__48566;
    wire N__48563;
    wire N__48560;
    wire N__48557;
    wire N__48554;
    wire N__48551;
    wire N__48548;
    wire N__48543;
    wire N__48540;
    wire N__48535;
    wire N__48528;
    wire N__48525;
    wire N__48520;
    wire N__48517;
    wire N__48510;
    wire N__48507;
    wire N__48504;
    wire N__48501;
    wire N__48498;
    wire N__48495;
    wire N__48492;
    wire N__48489;
    wire N__48486;
    wire N__48483;
    wire N__48480;
    wire N__48477;
    wire N__48474;
    wire N__48471;
    wire N__48468;
    wire N__48465;
    wire N__48462;
    wire N__48459;
    wire N__48456;
    wire N__48453;
    wire N__48450;
    wire N__48447;
    wire N__48444;
    wire N__48441;
    wire N__48438;
    wire N__48435;
    wire N__48432;
    wire N__48429;
    wire N__48426;
    wire N__48423;
    wire N__48420;
    wire N__48417;
    wire N__48414;
    wire N__48411;
    wire N__48410;
    wire N__48409;
    wire N__48408;
    wire N__48407;
    wire N__48404;
    wire N__48401;
    wire N__48398;
    wire N__48395;
    wire N__48392;
    wire N__48389;
    wire N__48384;
    wire N__48381;
    wire N__48378;
    wire N__48375;
    wire N__48370;
    wire N__48363;
    wire N__48360;
    wire N__48359;
    wire N__48358;
    wire N__48355;
    wire N__48350;
    wire N__48345;
    wire N__48342;
    wire N__48341;
    wire N__48338;
    wire N__48335;
    wire N__48330;
    wire N__48327;
    wire N__48324;
    wire N__48321;
    wire N__48318;
    wire N__48315;
    wire N__48312;
    wire N__48309;
    wire N__48306;
    wire N__48303;
    wire N__48300;
    wire N__48297;
    wire N__48294;
    wire N__48293;
    wire N__48290;
    wire N__48287;
    wire N__48284;
    wire N__48281;
    wire N__48276;
    wire N__48273;
    wire N__48270;
    wire N__48267;
    wire N__48266;
    wire N__48263;
    wire N__48260;
    wire N__48259;
    wire N__48258;
    wire N__48257;
    wire N__48254;
    wire N__48251;
    wire N__48248;
    wire N__48245;
    wire N__48242;
    wire N__48241;
    wire N__48238;
    wire N__48237;
    wire N__48232;
    wire N__48229;
    wire N__48226;
    wire N__48223;
    wire N__48220;
    wire N__48217;
    wire N__48208;
    wire N__48201;
    wire N__48198;
    wire N__48195;
    wire N__48192;
    wire N__48189;
    wire N__48188;
    wire N__48185;
    wire N__48182;
    wire N__48177;
    wire N__48174;
    wire N__48171;
    wire N__48168;
    wire N__48165;
    wire N__48162;
    wire N__48161;
    wire N__48156;
    wire N__48153;
    wire N__48150;
    wire N__48147;
    wire N__48144;
    wire N__48141;
    wire N__48140;
    wire N__48139;
    wire N__48138;
    wire N__48137;
    wire N__48134;
    wire N__48131;
    wire N__48128;
    wire N__48125;
    wire N__48122;
    wire N__48117;
    wire N__48110;
    wire N__48107;
    wire N__48104;
    wire N__48099;
    wire N__48096;
    wire N__48093;
    wire N__48090;
    wire N__48087;
    wire N__48084;
    wire N__48081;
    wire N__48078;
    wire N__48075;
    wire N__48072;
    wire N__48069;
    wire N__48066;
    wire N__48063;
    wire N__48060;
    wire N__48057;
    wire N__48054;
    wire N__48051;
    wire N__48048;
    wire N__48045;
    wire N__48042;
    wire N__48039;
    wire N__48036;
    wire N__48033;
    wire N__48030;
    wire N__48027;
    wire N__48024;
    wire N__48021;
    wire N__48018;
    wire N__48015;
    wire N__48012;
    wire N__48009;
    wire N__48006;
    wire N__48003;
    wire N__48000;
    wire N__47997;
    wire N__47994;
    wire N__47991;
    wire N__47988;
    wire N__47985;
    wire N__47982;
    wire N__47979;
    wire N__47976;
    wire N__47973;
    wire N__47970;
    wire N__47967;
    wire N__47964;
    wire N__47961;
    wire N__47958;
    wire N__47955;
    wire N__47952;
    wire N__47949;
    wire N__47946;
    wire N__47943;
    wire N__47940;
    wire N__47937;
    wire N__47934;
    wire N__47931;
    wire N__47928;
    wire N__47925;
    wire N__47924;
    wire N__47923;
    wire N__47922;
    wire N__47921;
    wire N__47920;
    wire N__47917;
    wire N__47916;
    wire N__47911;
    wire N__47910;
    wire N__47909;
    wire N__47908;
    wire N__47907;
    wire N__47906;
    wire N__47905;
    wire N__47902;
    wire N__47899;
    wire N__47896;
    wire N__47893;
    wire N__47890;
    wire N__47887;
    wire N__47882;
    wire N__47873;
    wire N__47868;
    wire N__47865;
    wire N__47864;
    wire N__47863;
    wire N__47862;
    wire N__47859;
    wire N__47856;
    wire N__47847;
    wire N__47844;
    wire N__47841;
    wire N__47836;
    wire N__47829;
    wire N__47820;
    wire N__47819;
    wire N__47816;
    wire N__47815;
    wire N__47812;
    wire N__47809;
    wire N__47806;
    wire N__47803;
    wire N__47800;
    wire N__47799;
    wire N__47796;
    wire N__47791;
    wire N__47788;
    wire N__47787;
    wire N__47786;
    wire N__47783;
    wire N__47778;
    wire N__47775;
    wire N__47774;
    wire N__47771;
    wire N__47768;
    wire N__47763;
    wire N__47760;
    wire N__47759;
    wire N__47756;
    wire N__47751;
    wire N__47748;
    wire N__47745;
    wire N__47742;
    wire N__47733;
    wire N__47730;
    wire N__47729;
    wire N__47728;
    wire N__47725;
    wire N__47724;
    wire N__47723;
    wire N__47722;
    wire N__47721;
    wire N__47718;
    wire N__47717;
    wire N__47716;
    wire N__47713;
    wire N__47712;
    wire N__47711;
    wire N__47710;
    wire N__47709;
    wire N__47708;
    wire N__47707;
    wire N__47706;
    wire N__47705;
    wire N__47704;
    wire N__47703;
    wire N__47702;
    wire N__47701;
    wire N__47700;
    wire N__47699;
    wire N__47698;
    wire N__47697;
    wire N__47696;
    wire N__47695;
    wire N__47694;
    wire N__47693;
    wire N__47692;
    wire N__47691;
    wire N__47688;
    wire N__47679;
    wire N__47678;
    wire N__47677;
    wire N__47676;
    wire N__47675;
    wire N__47674;
    wire N__47673;
    wire N__47672;
    wire N__47671;
    wire N__47668;
    wire N__47667;
    wire N__47666;
    wire N__47665;
    wire N__47664;
    wire N__47663;
    wire N__47662;
    wire N__47661;
    wire N__47658;
    wire N__47649;
    wire N__47644;
    wire N__47643;
    wire N__47642;
    wire N__47639;
    wire N__47638;
    wire N__47637;
    wire N__47628;
    wire N__47625;
    wire N__47622;
    wire N__47613;
    wire N__47608;
    wire N__47605;
    wire N__47602;
    wire N__47601;
    wire N__47594;
    wire N__47589;
    wire N__47578;
    wire N__47571;
    wire N__47568;
    wire N__47565;
    wire N__47564;
    wire N__47563;
    wire N__47560;
    wire N__47557;
    wire N__47548;
    wire N__47541;
    wire N__47538;
    wire N__47537;
    wire N__47536;
    wire N__47533;
    wire N__47532;
    wire N__47531;
    wire N__47530;
    wire N__47529;
    wire N__47524;
    wire N__47521;
    wire N__47520;
    wire N__47519;
    wire N__47518;
    wire N__47517;
    wire N__47516;
    wire N__47515;
    wire N__47510;
    wire N__47507;
    wire N__47502;
    wire N__47501;
    wire N__47500;
    wire N__47495;
    wire N__47492;
    wire N__47485;
    wire N__47478;
    wire N__47473;
    wire N__47468;
    wire N__47461;
    wire N__47458;
    wire N__47457;
    wire N__47454;
    wire N__47453;
    wire N__47452;
    wire N__47451;
    wire N__47450;
    wire N__47449;
    wire N__47446;
    wire N__47443;
    wire N__47436;
    wire N__47431;
    wire N__47424;
    wire N__47419;
    wire N__47416;
    wire N__47409;
    wire N__47404;
    wire N__47397;
    wire N__47394;
    wire N__47387;
    wire N__47384;
    wire N__47381;
    wire N__47378;
    wire N__47375;
    wire N__47370;
    wire N__47365;
    wire N__47360;
    wire N__47347;
    wire N__47342;
    wire N__47337;
    wire N__47316;
    wire N__47313;
    wire N__47310;
    wire N__47307;
    wire N__47304;
    wire N__47301;
    wire N__47298;
    wire N__47295;
    wire N__47292;
    wire N__47289;
    wire N__47286;
    wire N__47283;
    wire N__47280;
    wire N__47277;
    wire N__47274;
    wire N__47271;
    wire N__47270;
    wire N__47269;
    wire N__47268;
    wire N__47267;
    wire N__47264;
    wire N__47263;
    wire N__47262;
    wire N__47259;
    wire N__47258;
    wire N__47257;
    wire N__47256;
    wire N__47255;
    wire N__47254;
    wire N__47253;
    wire N__47252;
    wire N__47251;
    wire N__47250;
    wire N__47249;
    wire N__47246;
    wire N__47245;
    wire N__47244;
    wire N__47243;
    wire N__47240;
    wire N__47237;
    wire N__47234;
    wire N__47233;
    wire N__47232;
    wire N__47227;
    wire N__47224;
    wire N__47221;
    wire N__47218;
    wire N__47215;
    wire N__47212;
    wire N__47209;
    wire N__47204;
    wire N__47197;
    wire N__47196;
    wire N__47195;
    wire N__47194;
    wire N__47193;
    wire N__47192;
    wire N__47191;
    wire N__47190;
    wire N__47187;
    wire N__47182;
    wire N__47179;
    wire N__47176;
    wire N__47171;
    wire N__47166;
    wire N__47165;
    wire N__47164;
    wire N__47163;
    wire N__47160;
    wire N__47159;
    wire N__47158;
    wire N__47155;
    wire N__47154;
    wire N__47153;
    wire N__47150;
    wire N__47137;
    wire N__47136;
    wire N__47135;
    wire N__47134;
    wire N__47133;
    wire N__47132;
    wire N__47131;
    wire N__47128;
    wire N__47123;
    wire N__47120;
    wire N__47117;
    wire N__47112;
    wire N__47107;
    wire N__47098;
    wire N__47095;
    wire N__47092;
    wire N__47091;
    wire N__47088;
    wire N__47085;
    wire N__47080;
    wire N__47077;
    wire N__47072;
    wire N__47067;
    wire N__47058;
    wire N__47055;
    wire N__47052;
    wire N__47049;
    wire N__47048;
    wire N__47041;
    wire N__47034;
    wire N__47029;
    wire N__47026;
    wire N__47009;
    wire N__47006;
    wire N__47003;
    wire N__47000;
    wire N__46997;
    wire N__46994;
    wire N__46991;
    wire N__46986;
    wire N__46971;
    wire N__46968;
    wire N__46965;
    wire N__46962;
    wire N__46959;
    wire N__46958;
    wire N__46957;
    wire N__46954;
    wire N__46951;
    wire N__46948;
    wire N__46943;
    wire N__46938;
    wire N__46935;
    wire N__46934;
    wire N__46931;
    wire N__46928;
    wire N__46925;
    wire N__46922;
    wire N__46917;
    wire N__46916;
    wire N__46915;
    wire N__46914;
    wire N__46911;
    wire N__46910;
    wire N__46909;
    wire N__46906;
    wire N__46903;
    wire N__46900;
    wire N__46899;
    wire N__46898;
    wire N__46895;
    wire N__46894;
    wire N__46891;
    wire N__46890;
    wire N__46889;
    wire N__46886;
    wire N__46885;
    wire N__46878;
    wire N__46875;
    wire N__46874;
    wire N__46873;
    wire N__46872;
    wire N__46869;
    wire N__46866;
    wire N__46859;
    wire N__46856;
    wire N__46853;
    wire N__46850;
    wire N__46847;
    wire N__46842;
    wire N__46839;
    wire N__46836;
    wire N__46833;
    wire N__46828;
    wire N__46823;
    wire N__46818;
    wire N__46811;
    wire N__46810;
    wire N__46807;
    wire N__46804;
    wire N__46801;
    wire N__46796;
    wire N__46793;
    wire N__46790;
    wire N__46787;
    wire N__46784;
    wire N__46781;
    wire N__46770;
    wire N__46767;
    wire N__46766;
    wire N__46765;
    wire N__46764;
    wire N__46763;
    wire N__46760;
    wire N__46757;
    wire N__46756;
    wire N__46755;
    wire N__46754;
    wire N__46747;
    wire N__46746;
    wire N__46745;
    wire N__46742;
    wire N__46739;
    wire N__46734;
    wire N__46733;
    wire N__46732;
    wire N__46729;
    wire N__46726;
    wire N__46723;
    wire N__46720;
    wire N__46717;
    wire N__46712;
    wire N__46709;
    wire N__46706;
    wire N__46703;
    wire N__46700;
    wire N__46697;
    wire N__46696;
    wire N__46689;
    wire N__46686;
    wire N__46681;
    wire N__46676;
    wire N__46673;
    wire N__46670;
    wire N__46665;
    wire N__46662;
    wire N__46653;
    wire N__46650;
    wire N__46647;
    wire N__46644;
    wire N__46641;
    wire N__46640;
    wire N__46637;
    wire N__46634;
    wire N__46631;
    wire N__46628;
    wire N__46625;
    wire N__46620;
    wire N__46617;
    wire N__46616;
    wire N__46613;
    wire N__46610;
    wire N__46607;
    wire N__46602;
    wire N__46599;
    wire N__46598;
    wire N__46595;
    wire N__46594;
    wire N__46591;
    wire N__46588;
    wire N__46585;
    wire N__46578;
    wire N__46575;
    wire N__46572;
    wire N__46571;
    wire N__46568;
    wire N__46567;
    wire N__46564;
    wire N__46561;
    wire N__46558;
    wire N__46551;
    wire N__46548;
    wire N__46545;
    wire N__46544;
    wire N__46541;
    wire N__46538;
    wire N__46535;
    wire N__46530;
    wire N__46527;
    wire N__46526;
    wire N__46523;
    wire N__46520;
    wire N__46519;
    wire N__46516;
    wire N__46513;
    wire N__46510;
    wire N__46505;
    wire N__46500;
    wire N__46497;
    wire N__46494;
    wire N__46491;
    wire N__46488;
    wire N__46485;
    wire N__46484;
    wire N__46483;
    wire N__46482;
    wire N__46481;
    wire N__46480;
    wire N__46479;
    wire N__46478;
    wire N__46477;
    wire N__46476;
    wire N__46475;
    wire N__46474;
    wire N__46473;
    wire N__46472;
    wire N__46471;
    wire N__46470;
    wire N__46469;
    wire N__46468;
    wire N__46467;
    wire N__46466;
    wire N__46465;
    wire N__46464;
    wire N__46463;
    wire N__46462;
    wire N__46461;
    wire N__46460;
    wire N__46459;
    wire N__46458;
    wire N__46457;
    wire N__46456;
    wire N__46455;
    wire N__46454;
    wire N__46453;
    wire N__46450;
    wire N__46445;
    wire N__46438;
    wire N__46433;
    wire N__46430;
    wire N__46425;
    wire N__46418;
    wire N__46415;
    wire N__46412;
    wire N__46411;
    wire N__46410;
    wire N__46409;
    wire N__46408;
    wire N__46407;
    wire N__46406;
    wire N__46403;
    wire N__46402;
    wire N__46397;
    wire N__46392;
    wire N__46387;
    wire N__46384;
    wire N__46381;
    wire N__46378;
    wire N__46377;
    wire N__46376;
    wire N__46375;
    wire N__46374;
    wire N__46373;
    wire N__46372;
    wire N__46371;
    wire N__46370;
    wire N__46369;
    wire N__46360;
    wire N__46357;
    wire N__46354;
    wire N__46351;
    wire N__46346;
    wire N__46339;
    wire N__46336;
    wire N__46329;
    wire N__46324;
    wire N__46319;
    wire N__46318;
    wire N__46317;
    wire N__46312;
    wire N__46311;
    wire N__46310;
    wire N__46309;
    wire N__46308;
    wire N__46307;
    wire N__46306;
    wire N__46303;
    wire N__46302;
    wire N__46301;
    wire N__46300;
    wire N__46299;
    wire N__46298;
    wire N__46297;
    wire N__46296;
    wire N__46295;
    wire N__46292;
    wire N__46291;
    wire N__46290;
    wire N__46287;
    wire N__46278;
    wire N__46275;
    wire N__46272;
    wire N__46269;
    wire N__46262;
    wire N__46259;
    wire N__46258;
    wire N__46257;
    wire N__46256;
    wire N__46249;
    wire N__46244;
    wire N__46241;
    wire N__46238;
    wire N__46225;
    wire N__46224;
    wire N__46221;
    wire N__46218;
    wire N__46215;
    wire N__46210;
    wire N__46203;
    wire N__46200;
    wire N__46197;
    wire N__46186;
    wire N__46183;
    wire N__46178;
    wire N__46175;
    wire N__46172;
    wire N__46169;
    wire N__46160;
    wire N__46159;
    wire N__46152;
    wire N__46149;
    wire N__46146;
    wire N__46143;
    wire N__46132;
    wire N__46129;
    wire N__46122;
    wire N__46111;
    wire N__46098;
    wire N__46095;
    wire N__46092;
    wire N__46089;
    wire N__46084;
    wire N__46081;
    wire N__46072;
    wire N__46059;
    wire N__46056;
    wire N__46053;
    wire N__46050;
    wire N__46047;
    wire N__46044;
    wire N__46041;
    wire N__46038;
    wire N__46037;
    wire N__46036;
    wire N__46033;
    wire N__46030;
    wire N__46027;
    wire N__46024;
    wire N__46021;
    wire N__46018;
    wire N__46015;
    wire N__46010;
    wire N__46005;
    wire N__46002;
    wire N__45999;
    wire N__45996;
    wire N__45993;
    wire N__45990;
    wire N__45987;
    wire N__45984;
    wire N__45981;
    wire N__45978;
    wire N__45975;
    wire N__45972;
    wire N__45969;
    wire N__45966;
    wire N__45963;
    wire N__45960;
    wire N__45957;
    wire N__45954;
    wire N__45951;
    wire N__45948;
    wire N__45945;
    wire N__45942;
    wire N__45939;
    wire N__45936;
    wire N__45933;
    wire N__45930;
    wire N__45927;
    wire N__45924;
    wire N__45921;
    wire N__45918;
    wire N__45915;
    wire N__45912;
    wire N__45909;
    wire N__45906;
    wire N__45903;
    wire N__45902;
    wire N__45899;
    wire N__45896;
    wire N__45891;
    wire N__45888;
    wire N__45885;
    wire N__45882;
    wire N__45879;
    wire N__45878;
    wire N__45875;
    wire N__45874;
    wire N__45871;
    wire N__45870;
    wire N__45869;
    wire N__45868;
    wire N__45865;
    wire N__45864;
    wire N__45861;
    wire N__45858;
    wire N__45855;
    wire N__45852;
    wire N__45849;
    wire N__45848;
    wire N__45845;
    wire N__45842;
    wire N__45839;
    wire N__45836;
    wire N__45833;
    wire N__45830;
    wire N__45829;
    wire N__45824;
    wire N__45821;
    wire N__45818;
    wire N__45809;
    wire N__45806;
    wire N__45803;
    wire N__45800;
    wire N__45797;
    wire N__45794;
    wire N__45791;
    wire N__45788;
    wire N__45785;
    wire N__45782;
    wire N__45775;
    wire N__45768;
    wire N__45765;
    wire N__45762;
    wire N__45759;
    wire N__45756;
    wire N__45753;
    wire N__45750;
    wire N__45747;
    wire N__45744;
    wire N__45741;
    wire N__45738;
    wire N__45735;
    wire N__45732;
    wire N__45729;
    wire N__45728;
    wire N__45725;
    wire N__45722;
    wire N__45719;
    wire N__45718;
    wire N__45715;
    wire N__45712;
    wire N__45709;
    wire N__45706;
    wire N__45699;
    wire N__45696;
    wire N__45693;
    wire N__45690;
    wire N__45687;
    wire N__45684;
    wire N__45681;
    wire N__45678;
    wire N__45677;
    wire N__45674;
    wire N__45671;
    wire N__45670;
    wire N__45669;
    wire N__45666;
    wire N__45663;
    wire N__45658;
    wire N__45651;
    wire N__45648;
    wire N__45647;
    wire N__45646;
    wire N__45645;
    wire N__45642;
    wire N__45639;
    wire N__45636;
    wire N__45635;
    wire N__45634;
    wire N__45631;
    wire N__45628;
    wire N__45625;
    wire N__45622;
    wire N__45621;
    wire N__45620;
    wire N__45617;
    wire N__45616;
    wire N__45613;
    wire N__45610;
    wire N__45605;
    wire N__45602;
    wire N__45599;
    wire N__45596;
    wire N__45593;
    wire N__45590;
    wire N__45585;
    wire N__45582;
    wire N__45579;
    wire N__45576;
    wire N__45573;
    wire N__45568;
    wire N__45563;
    wire N__45554;
    wire N__45549;
    wire N__45546;
    wire N__45543;
    wire N__45540;
    wire N__45537;
    wire N__45534;
    wire N__45531;
    wire N__45528;
    wire N__45525;
    wire N__45522;
    wire N__45519;
    wire N__45516;
    wire N__45513;
    wire N__45510;
    wire N__45507;
    wire N__45504;
    wire N__45501;
    wire N__45498;
    wire N__45495;
    wire N__45492;
    wire N__45489;
    wire N__45486;
    wire N__45483;
    wire N__45480;
    wire N__45479;
    wire N__45476;
    wire N__45475;
    wire N__45472;
    wire N__45469;
    wire N__45466;
    wire N__45465;
    wire N__45462;
    wire N__45459;
    wire N__45456;
    wire N__45453;
    wire N__45450;
    wire N__45445;
    wire N__45442;
    wire N__45439;
    wire N__45434;
    wire N__45431;
    wire N__45428;
    wire N__45423;
    wire N__45420;
    wire N__45417;
    wire N__45414;
    wire N__45411;
    wire N__45408;
    wire N__45405;
    wire N__45402;
    wire N__45399;
    wire N__45396;
    wire N__45393;
    wire N__45390;
    wire N__45389;
    wire N__45388;
    wire N__45385;
    wire N__45382;
    wire N__45377;
    wire N__45374;
    wire N__45371;
    wire N__45366;
    wire N__45363;
    wire N__45360;
    wire N__45357;
    wire N__45356;
    wire N__45353;
    wire N__45352;
    wire N__45349;
    wire N__45348;
    wire N__45345;
    wire N__45342;
    wire N__45339;
    wire N__45336;
    wire N__45335;
    wire N__45334;
    wire N__45327;
    wire N__45326;
    wire N__45323;
    wire N__45320;
    wire N__45317;
    wire N__45314;
    wire N__45311;
    wire N__45306;
    wire N__45303;
    wire N__45302;
    wire N__45293;
    wire N__45290;
    wire N__45285;
    wire N__45282;
    wire N__45281;
    wire N__45280;
    wire N__45275;
    wire N__45272;
    wire N__45269;
    wire N__45266;
    wire N__45263;
    wire N__45260;
    wire N__45257;
    wire N__45252;
    wire N__45249;
    wire N__45246;
    wire N__45243;
    wire N__45240;
    wire N__45237;
    wire N__45234;
    wire N__45231;
    wire N__45228;
    wire N__45225;
    wire N__45222;
    wire N__45219;
    wire N__45216;
    wire N__45213;
    wire N__45212;
    wire N__45211;
    wire N__45210;
    wire N__45209;
    wire N__45206;
    wire N__45203;
    wire N__45200;
    wire N__45199;
    wire N__45196;
    wire N__45195;
    wire N__45194;
    wire N__45191;
    wire N__45186;
    wire N__45183;
    wire N__45180;
    wire N__45177;
    wire N__45174;
    wire N__45171;
    wire N__45170;
    wire N__45167;
    wire N__45164;
    wire N__45157;
    wire N__45154;
    wire N__45151;
    wire N__45148;
    wire N__45145;
    wire N__45140;
    wire N__45133;
    wire N__45126;
    wire N__45123;
    wire N__45120;
    wire N__45117;
    wire N__45114;
    wire N__45111;
    wire N__45108;
    wire N__45105;
    wire N__45102;
    wire N__45099;
    wire N__45096;
    wire N__45093;
    wire N__45090;
    wire N__45087;
    wire N__45084;
    wire N__45081;
    wire N__45078;
    wire N__45075;
    wire N__45072;
    wire N__45069;
    wire N__45066;
    wire N__45063;
    wire N__45060;
    wire N__45059;
    wire N__45056;
    wire N__45053;
    wire N__45050;
    wire N__45047;
    wire N__45042;
    wire N__45039;
    wire N__45036;
    wire N__45033;
    wire N__45032;
    wire N__45029;
    wire N__45026;
    wire N__45025;
    wire N__45020;
    wire N__45017;
    wire N__45016;
    wire N__45011;
    wire N__45008;
    wire N__45005;
    wire N__45000;
    wire N__44997;
    wire N__44994;
    wire N__44993;
    wire N__44992;
    wire N__44989;
    wire N__44986;
    wire N__44983;
    wire N__44976;
    wire N__44973;
    wire N__44970;
    wire N__44969;
    wire N__44968;
    wire N__44967;
    wire N__44964;
    wire N__44959;
    wire N__44956;
    wire N__44949;
    wire N__44946;
    wire N__44943;
    wire N__44940;
    wire N__44937;
    wire N__44934;
    wire N__44931;
    wire N__44928;
    wire N__44925;
    wire N__44922;
    wire N__44919;
    wire N__44916;
    wire N__44913;
    wire N__44910;
    wire N__44907;
    wire N__44904;
    wire N__44901;
    wire N__44898;
    wire N__44895;
    wire N__44892;
    wire N__44889;
    wire N__44886;
    wire N__44883;
    wire N__44880;
    wire N__44877;
    wire N__44874;
    wire N__44871;
    wire N__44868;
    wire N__44865;
    wire N__44862;
    wire N__44859;
    wire N__44856;
    wire N__44853;
    wire N__44850;
    wire N__44847;
    wire N__44844;
    wire N__44841;
    wire N__44838;
    wire N__44835;
    wire N__44832;
    wire N__44829;
    wire N__44826;
    wire N__44823;
    wire N__44822;
    wire N__44819;
    wire N__44816;
    wire N__44815;
    wire N__44810;
    wire N__44807;
    wire N__44804;
    wire N__44799;
    wire N__44796;
    wire N__44793;
    wire N__44792;
    wire N__44791;
    wire N__44788;
    wire N__44785;
    wire N__44782;
    wire N__44775;
    wire N__44772;
    wire N__44769;
    wire N__44766;
    wire N__44763;
    wire N__44760;
    wire N__44757;
    wire N__44754;
    wire N__44753;
    wire N__44752;
    wire N__44749;
    wire N__44748;
    wire N__44745;
    wire N__44744;
    wire N__44741;
    wire N__44738;
    wire N__44735;
    wire N__44730;
    wire N__44727;
    wire N__44726;
    wire N__44719;
    wire N__44716;
    wire N__44713;
    wire N__44710;
    wire N__44709;
    wire N__44708;
    wire N__44703;
    wire N__44702;
    wire N__44699;
    wire N__44696;
    wire N__44693;
    wire N__44690;
    wire N__44687;
    wire N__44684;
    wire N__44679;
    wire N__44670;
    wire N__44669;
    wire N__44668;
    wire N__44667;
    wire N__44664;
    wire N__44661;
    wire N__44658;
    wire N__44657;
    wire N__44654;
    wire N__44653;
    wire N__44652;
    wire N__44651;
    wire N__44650;
    wire N__44649;
    wire N__44648;
    wire N__44647;
    wire N__44646;
    wire N__44645;
    wire N__44644;
    wire N__44643;
    wire N__44642;
    wire N__44641;
    wire N__44640;
    wire N__44639;
    wire N__44638;
    wire N__44633;
    wire N__44630;
    wire N__44629;
    wire N__44628;
    wire N__44627;
    wire N__44626;
    wire N__44623;
    wire N__44620;
    wire N__44617;
    wire N__44602;
    wire N__44585;
    wire N__44582;
    wire N__44579;
    wire N__44570;
    wire N__44565;
    wire N__44550;
    wire N__44547;
    wire N__44544;
    wire N__44543;
    wire N__44540;
    wire N__44537;
    wire N__44534;
    wire N__44531;
    wire N__44528;
    wire N__44525;
    wire N__44520;
    wire N__44517;
    wire N__44516;
    wire N__44515;
    wire N__44512;
    wire N__44509;
    wire N__44508;
    wire N__44505;
    wire N__44504;
    wire N__44503;
    wire N__44500;
    wire N__44499;
    wire N__44498;
    wire N__44497;
    wire N__44496;
    wire N__44495;
    wire N__44494;
    wire N__44493;
    wire N__44492;
    wire N__44491;
    wire N__44488;
    wire N__44485;
    wire N__44482;
    wire N__44479;
    wire N__44476;
    wire N__44473;
    wire N__44456;
    wire N__44455;
    wire N__44454;
    wire N__44453;
    wire N__44452;
    wire N__44451;
    wire N__44450;
    wire N__44449;
    wire N__44446;
    wire N__44445;
    wire N__44444;
    wire N__44439;
    wire N__44436;
    wire N__44433;
    wire N__44430;
    wire N__44425;
    wire N__44410;
    wire N__44409;
    wire N__44408;
    wire N__44401;
    wire N__44394;
    wire N__44389;
    wire N__44388;
    wire N__44385;
    wire N__44380;
    wire N__44377;
    wire N__44376;
    wire N__44373;
    wire N__44370;
    wire N__44367;
    wire N__44360;
    wire N__44357;
    wire N__44354;
    wire N__44343;
    wire N__44340;
    wire N__44337;
    wire N__44334;
    wire N__44331;
    wire N__44330;
    wire N__44327;
    wire N__44324;
    wire N__44323;
    wire N__44320;
    wire N__44317;
    wire N__44314;
    wire N__44313;
    wire N__44312;
    wire N__44311;
    wire N__44304;
    wire N__44301;
    wire N__44298;
    wire N__44295;
    wire N__44288;
    wire N__44283;
    wire N__44280;
    wire N__44277;
    wire N__44274;
    wire N__44271;
    wire N__44268;
    wire N__44265;
    wire N__44262;
    wire N__44259;
    wire N__44256;
    wire N__44253;
    wire N__44250;
    wire N__44247;
    wire N__44244;
    wire N__44241;
    wire N__44238;
    wire N__44235;
    wire N__44232;
    wire N__44229;
    wire N__44226;
    wire N__44223;
    wire N__44220;
    wire N__44217;
    wire N__44214;
    wire N__44213;
    wire N__44210;
    wire N__44207;
    wire N__44204;
    wire N__44199;
    wire N__44196;
    wire N__44195;
    wire N__44194;
    wire N__44191;
    wire N__44188;
    wire N__44185;
    wire N__44182;
    wire N__44175;
    wire N__44172;
    wire N__44169;
    wire N__44166;
    wire N__44165;
    wire N__44164;
    wire N__44161;
    wire N__44156;
    wire N__44151;
    wire N__44148;
    wire N__44145;
    wire N__44142;
    wire N__44141;
    wire N__44140;
    wire N__44137;
    wire N__44132;
    wire N__44127;
    wire N__44124;
    wire N__44121;
    wire N__44118;
    wire N__44115;
    wire N__44114;
    wire N__44111;
    wire N__44108;
    wire N__44105;
    wire N__44102;
    wire N__44099;
    wire N__44096;
    wire N__44093;
    wire N__44090;
    wire N__44087;
    wire N__44082;
    wire N__44079;
    wire N__44078;
    wire N__44075;
    wire N__44072;
    wire N__44071;
    wire N__44068;
    wire N__44065;
    wire N__44062;
    wire N__44061;
    wire N__44060;
    wire N__44059;
    wire N__44054;
    wire N__44051;
    wire N__44048;
    wire N__44043;
    wire N__44040;
    wire N__44037;
    wire N__44032;
    wire N__44029;
    wire N__44026;
    wire N__44023;
    wire N__44016;
    wire N__44015;
    wire N__44014;
    wire N__44013;
    wire N__44010;
    wire N__44009;
    wire N__44006;
    wire N__44003;
    wire N__44002;
    wire N__44001;
    wire N__43998;
    wire N__43995;
    wire N__43992;
    wire N__43989;
    wire N__43986;
    wire N__43983;
    wire N__43980;
    wire N__43973;
    wire N__43966;
    wire N__43963;
    wire N__43962;
    wire N__43957;
    wire N__43954;
    wire N__43951;
    wire N__43944;
    wire N__43943;
    wire N__43940;
    wire N__43937;
    wire N__43936;
    wire N__43933;
    wire N__43930;
    wire N__43927;
    wire N__43926;
    wire N__43921;
    wire N__43916;
    wire N__43911;
    wire N__43910;
    wire N__43907;
    wire N__43904;
    wire N__43903;
    wire N__43900;
    wire N__43897;
    wire N__43894;
    wire N__43891;
    wire N__43888;
    wire N__43885;
    wire N__43882;
    wire N__43879;
    wire N__43876;
    wire N__43869;
    wire N__43866;
    wire N__43865;
    wire N__43862;
    wire N__43859;
    wire N__43856;
    wire N__43853;
    wire N__43850;
    wire N__43845;
    wire N__43844;
    wire N__43841;
    wire N__43840;
    wire N__43837;
    wire N__43834;
    wire N__43831;
    wire N__43828;
    wire N__43825;
    wire N__43818;
    wire N__43815;
    wire N__43812;
    wire N__43809;
    wire N__43806;
    wire N__43803;
    wire N__43800;
    wire N__43797;
    wire N__43794;
    wire N__43791;
    wire N__43788;
    wire N__43785;
    wire N__43782;
    wire N__43779;
    wire N__43776;
    wire N__43773;
    wire N__43770;
    wire N__43769;
    wire N__43766;
    wire N__43763;
    wire N__43758;
    wire N__43757;
    wire N__43754;
    wire N__43751;
    wire N__43748;
    wire N__43745;
    wire N__43742;
    wire N__43741;
    wire N__43738;
    wire N__43735;
    wire N__43732;
    wire N__43729;
    wire N__43726;
    wire N__43723;
    wire N__43720;
    wire N__43717;
    wire N__43710;
    wire N__43707;
    wire N__43704;
    wire N__43701;
    wire N__43698;
    wire N__43697;
    wire N__43694;
    wire N__43691;
    wire N__43686;
    wire N__43683;
    wire N__43680;
    wire N__43677;
    wire N__43676;
    wire N__43673;
    wire N__43672;
    wire N__43669;
    wire N__43666;
    wire N__43663;
    wire N__43656;
    wire N__43653;
    wire N__43650;
    wire N__43649;
    wire N__43648;
    wire N__43645;
    wire N__43642;
    wire N__43639;
    wire N__43636;
    wire N__43633;
    wire N__43626;
    wire N__43623;
    wire N__43620;
    wire N__43617;
    wire N__43614;
    wire N__43613;
    wire N__43610;
    wire N__43607;
    wire N__43602;
    wire N__43601;
    wire N__43598;
    wire N__43595;
    wire N__43592;
    wire N__43587;
    wire N__43584;
    wire N__43581;
    wire N__43578;
    wire N__43575;
    wire N__43572;
    wire N__43569;
    wire N__43566;
    wire N__43563;
    wire N__43560;
    wire N__43559;
    wire N__43556;
    wire N__43553;
    wire N__43550;
    wire N__43547;
    wire N__43542;
    wire N__43539;
    wire N__43538;
    wire N__43535;
    wire N__43534;
    wire N__43531;
    wire N__43528;
    wire N__43525;
    wire N__43518;
    wire N__43517;
    wire N__43514;
    wire N__43513;
    wire N__43510;
    wire N__43507;
    wire N__43504;
    wire N__43497;
    wire N__43494;
    wire N__43491;
    wire N__43488;
    wire N__43485;
    wire N__43482;
    wire N__43479;
    wire N__43476;
    wire N__43473;
    wire N__43472;
    wire N__43469;
    wire N__43466;
    wire N__43461;
    wire N__43458;
    wire N__43457;
    wire N__43454;
    wire N__43451;
    wire N__43448;
    wire N__43445;
    wire N__43442;
    wire N__43437;
    wire N__43436;
    wire N__43433;
    wire N__43432;
    wire N__43429;
    wire N__43426;
    wire N__43423;
    wire N__43416;
    wire N__43413;
    wire N__43410;
    wire N__43407;
    wire N__43404;
    wire N__43401;
    wire N__43398;
    wire N__43395;
    wire N__43392;
    wire N__43389;
    wire N__43388;
    wire N__43385;
    wire N__43382;
    wire N__43379;
    wire N__43378;
    wire N__43375;
    wire N__43372;
    wire N__43369;
    wire N__43364;
    wire N__43359;
    wire N__43356;
    wire N__43353;
    wire N__43350;
    wire N__43347;
    wire N__43344;
    wire N__43341;
    wire N__43338;
    wire N__43337;
    wire N__43336;
    wire N__43333;
    wire N__43330;
    wire N__43327;
    wire N__43326;
    wire N__43325;
    wire N__43324;
    wire N__43321;
    wire N__43318;
    wire N__43315;
    wire N__43312;
    wire N__43309;
    wire N__43306;
    wire N__43305;
    wire N__43302;
    wire N__43295;
    wire N__43292;
    wire N__43289;
    wire N__43286;
    wire N__43275;
    wire N__43274;
    wire N__43271;
    wire N__43268;
    wire N__43265;
    wire N__43264;
    wire N__43263;
    wire N__43260;
    wire N__43257;
    wire N__43254;
    wire N__43251;
    wire N__43250;
    wire N__43249;
    wire N__43242;
    wire N__43239;
    wire N__43236;
    wire N__43233;
    wire N__43230;
    wire N__43225;
    wire N__43222;
    wire N__43215;
    wire N__43212;
    wire N__43209;
    wire N__43206;
    wire N__43203;
    wire N__43200;
    wire N__43199;
    wire N__43198;
    wire N__43195;
    wire N__43194;
    wire N__43191;
    wire N__43188;
    wire N__43185;
    wire N__43182;
    wire N__43179;
    wire N__43176;
    wire N__43173;
    wire N__43170;
    wire N__43165;
    wire N__43162;
    wire N__43157;
    wire N__43152;
    wire N__43149;
    wire N__43146;
    wire N__43143;
    wire N__43140;
    wire N__43137;
    wire N__43134;
    wire N__43131;
    wire N__43128;
    wire N__43125;
    wire N__43122;
    wire N__43119;
    wire N__43116;
    wire N__43113;
    wire N__43110;
    wire N__43107;
    wire N__43106;
    wire N__43103;
    wire N__43100;
    wire N__43097;
    wire N__43094;
    wire N__43091;
    wire N__43086;
    wire N__43085;
    wire N__43082;
    wire N__43079;
    wire N__43078;
    wire N__43075;
    wire N__43072;
    wire N__43069;
    wire N__43064;
    wire N__43059;
    wire N__43056;
    wire N__43053;
    wire N__43050;
    wire N__43047;
    wire N__43044;
    wire N__43043;
    wire N__43042;
    wire N__43041;
    wire N__43038;
    wire N__43035;
    wire N__43032;
    wire N__43029;
    wire N__43028;
    wire N__43025;
    wire N__43018;
    wire N__43015;
    wire N__43012;
    wire N__43009;
    wire N__43002;
    wire N__42999;
    wire N__42996;
    wire N__42995;
    wire N__42994;
    wire N__42991;
    wire N__42986;
    wire N__42981;
    wire N__42978;
    wire N__42977;
    wire N__42974;
    wire N__42973;
    wire N__42970;
    wire N__42967;
    wire N__42964;
    wire N__42957;
    wire N__42954;
    wire N__42953;
    wire N__42950;
    wire N__42947;
    wire N__42944;
    wire N__42941;
    wire N__42938;
    wire N__42937;
    wire N__42934;
    wire N__42931;
    wire N__42928;
    wire N__42925;
    wire N__42918;
    wire N__42915;
    wire N__42912;
    wire N__42909;
    wire N__42906;
    wire N__42903;
    wire N__42900;
    wire N__42897;
    wire N__42894;
    wire N__42891;
    wire N__42888;
    wire N__42887;
    wire N__42884;
    wire N__42881;
    wire N__42880;
    wire N__42877;
    wire N__42874;
    wire N__42871;
    wire N__42866;
    wire N__42863;
    wire N__42860;
    wire N__42857;
    wire N__42852;
    wire N__42851;
    wire N__42848;
    wire N__42847;
    wire N__42840;
    wire N__42837;
    wire N__42836;
    wire N__42833;
    wire N__42830;
    wire N__42829;
    wire N__42826;
    wire N__42823;
    wire N__42820;
    wire N__42815;
    wire N__42812;
    wire N__42809;
    wire N__42806;
    wire N__42801;
    wire N__42798;
    wire N__42797;
    wire N__42796;
    wire N__42795;
    wire N__42792;
    wire N__42791;
    wire N__42788;
    wire N__42785;
    wire N__42782;
    wire N__42781;
    wire N__42780;
    wire N__42779;
    wire N__42778;
    wire N__42775;
    wire N__42772;
    wire N__42757;
    wire N__42750;
    wire N__42747;
    wire N__42746;
    wire N__42745;
    wire N__42744;
    wire N__42743;
    wire N__42742;
    wire N__42741;
    wire N__42740;
    wire N__42737;
    wire N__42722;
    wire N__42717;
    wire N__42714;
    wire N__42711;
    wire N__42710;
    wire N__42709;
    wire N__42708;
    wire N__42707;
    wire N__42704;
    wire N__42701;
    wire N__42698;
    wire N__42695;
    wire N__42692;
    wire N__42689;
    wire N__42686;
    wire N__42683;
    wire N__42680;
    wire N__42677;
    wire N__42672;
    wire N__42669;
    wire N__42666;
    wire N__42663;
    wire N__42660;
    wire N__42655;
    wire N__42648;
    wire N__42645;
    wire N__42642;
    wire N__42639;
    wire N__42636;
    wire N__42635;
    wire N__42632;
    wire N__42631;
    wire N__42630;
    wire N__42627;
    wire N__42624;
    wire N__42621;
    wire N__42618;
    wire N__42615;
    wire N__42612;
    wire N__42609;
    wire N__42606;
    wire N__42601;
    wire N__42598;
    wire N__42595;
    wire N__42588;
    wire N__42585;
    wire N__42582;
    wire N__42579;
    wire N__42576;
    wire N__42573;
    wire N__42570;
    wire N__42567;
    wire N__42564;
    wire N__42561;
    wire N__42558;
    wire N__42555;
    wire N__42554;
    wire N__42551;
    wire N__42550;
    wire N__42547;
    wire N__42544;
    wire N__42543;
    wire N__42542;
    wire N__42539;
    wire N__42536;
    wire N__42535;
    wire N__42532;
    wire N__42527;
    wire N__42524;
    wire N__42521;
    wire N__42518;
    wire N__42517;
    wire N__42512;
    wire N__42509;
    wire N__42504;
    wire N__42501;
    wire N__42498;
    wire N__42495;
    wire N__42490;
    wire N__42483;
    wire N__42480;
    wire N__42477;
    wire N__42474;
    wire N__42471;
    wire N__42468;
    wire N__42465;
    wire N__42462;
    wire N__42459;
    wire N__42456;
    wire N__42453;
    wire N__42450;
    wire N__42447;
    wire N__42446;
    wire N__42443;
    wire N__42440;
    wire N__42435;
    wire N__42434;
    wire N__42431;
    wire N__42430;
    wire N__42429;
    wire N__42426;
    wire N__42425;
    wire N__42424;
    wire N__42421;
    wire N__42418;
    wire N__42415;
    wire N__42414;
    wire N__42413;
    wire N__42412;
    wire N__42411;
    wire N__42410;
    wire N__42409;
    wire N__42406;
    wire N__42403;
    wire N__42400;
    wire N__42399;
    wire N__42398;
    wire N__42395;
    wire N__42394;
    wire N__42391;
    wire N__42388;
    wire N__42385;
    wire N__42384;
    wire N__42383;
    wire N__42380;
    wire N__42377;
    wire N__42374;
    wire N__42373;
    wire N__42372;
    wire N__42369;
    wire N__42366;
    wire N__42365;
    wire N__42364;
    wire N__42363;
    wire N__42362;
    wire N__42357;
    wire N__42354;
    wire N__42351;
    wire N__42348;
    wire N__42345;
    wire N__42342;
    wire N__42335;
    wire N__42334;
    wire N__42331;
    wire N__42328;
    wire N__42325;
    wire N__42320;
    wire N__42317;
    wire N__42314;
    wire N__42309;
    wire N__42306;
    wire N__42305;
    wire N__42302;
    wire N__42301;
    wire N__42298;
    wire N__42295;
    wire N__42286;
    wire N__42279;
    wire N__42276;
    wire N__42269;
    wire N__42264;
    wire N__42261;
    wire N__42256;
    wire N__42253;
    wire N__42250;
    wire N__42247;
    wire N__42244;
    wire N__42235;
    wire N__42230;
    wire N__42227;
    wire N__42222;
    wire N__42221;
    wire N__42218;
    wire N__42215;
    wire N__42212;
    wire N__42209;
    wire N__42204;
    wire N__42201;
    wire N__42198;
    wire N__42183;
    wire N__42180;
    wire N__42177;
    wire N__42174;
    wire N__42171;
    wire N__42168;
    wire N__42165;
    wire N__42162;
    wire N__42159;
    wire N__42156;
    wire N__42153;
    wire N__42152;
    wire N__42151;
    wire N__42148;
    wire N__42147;
    wire N__42144;
    wire N__42143;
    wire N__42140;
    wire N__42137;
    wire N__42134;
    wire N__42131;
    wire N__42128;
    wire N__42125;
    wire N__42120;
    wire N__42115;
    wire N__42112;
    wire N__42109;
    wire N__42102;
    wire N__42099;
    wire N__42096;
    wire N__42093;
    wire N__42090;
    wire N__42087;
    wire N__42084;
    wire N__42083;
    wire N__42080;
    wire N__42077;
    wire N__42072;
    wire N__42069;
    wire N__42066;
    wire N__42063;
    wire N__42060;
    wire N__42057;
    wire N__42054;
    wire N__42051;
    wire N__42050;
    wire N__42047;
    wire N__42046;
    wire N__42043;
    wire N__42040;
    wire N__42037;
    wire N__42032;
    wire N__42029;
    wire N__42026;
    wire N__42021;
    wire N__42018;
    wire N__42015;
    wire N__42012;
    wire N__42009;
    wire N__42008;
    wire N__42005;
    wire N__42002;
    wire N__42001;
    wire N__41998;
    wire N__41995;
    wire N__41992;
    wire N__41991;
    wire N__41990;
    wire N__41989;
    wire N__41988;
    wire N__41985;
    wire N__41982;
    wire N__41979;
    wire N__41974;
    wire N__41969;
    wire N__41966;
    wire N__41963;
    wire N__41960;
    wire N__41949;
    wire N__41946;
    wire N__41943;
    wire N__41940;
    wire N__41937;
    wire N__41934;
    wire N__41931;
    wire N__41928;
    wire N__41925;
    wire N__41922;
    wire N__41919;
    wire N__41916;
    wire N__41915;
    wire N__41912;
    wire N__41909;
    wire N__41904;
    wire N__41901;
    wire N__41900;
    wire N__41897;
    wire N__41894;
    wire N__41891;
    wire N__41886;
    wire N__41883;
    wire N__41880;
    wire N__41877;
    wire N__41874;
    wire N__41871;
    wire N__41868;
    wire N__41865;
    wire N__41862;
    wire N__41859;
    wire N__41856;
    wire N__41853;
    wire N__41850;
    wire N__41847;
    wire N__41844;
    wire N__41843;
    wire N__41840;
    wire N__41837;
    wire N__41834;
    wire N__41831;
    wire N__41828;
    wire N__41825;
    wire N__41822;
    wire N__41819;
    wire N__41816;
    wire N__41813;
    wire N__41810;
    wire N__41807;
    wire N__41804;
    wire N__41799;
    wire N__41798;
    wire N__41795;
    wire N__41792;
    wire N__41787;
    wire N__41784;
    wire N__41783;
    wire N__41780;
    wire N__41777;
    wire N__41772;
    wire N__41769;
    wire N__41766;
    wire N__41763;
    wire N__41760;
    wire N__41757;
    wire N__41754;
    wire N__41751;
    wire N__41748;
    wire N__41745;
    wire N__41742;
    wire N__41739;
    wire N__41736;
    wire N__41733;
    wire N__41730;
    wire N__41727;
    wire N__41724;
    wire N__41723;
    wire N__41722;
    wire N__41719;
    wire N__41714;
    wire N__41709;
    wire N__41706;
    wire N__41705;
    wire N__41702;
    wire N__41701;
    wire N__41698;
    wire N__41695;
    wire N__41692;
    wire N__41689;
    wire N__41686;
    wire N__41683;
    wire N__41680;
    wire N__41677;
    wire N__41670;
    wire N__41669;
    wire N__41668;
    wire N__41667;
    wire N__41666;
    wire N__41665;
    wire N__41664;
    wire N__41663;
    wire N__41662;
    wire N__41659;
    wire N__41658;
    wire N__41657;
    wire N__41654;
    wire N__41651;
    wire N__41648;
    wire N__41645;
    wire N__41644;
    wire N__41641;
    wire N__41638;
    wire N__41637;
    wire N__41634;
    wire N__41631;
    wire N__41628;
    wire N__41625;
    wire N__41622;
    wire N__41619;
    wire N__41616;
    wire N__41615;
    wire N__41614;
    wire N__41613;
    wire N__41610;
    wire N__41607;
    wire N__41604;
    wire N__41599;
    wire N__41596;
    wire N__41591;
    wire N__41584;
    wire N__41579;
    wire N__41574;
    wire N__41571;
    wire N__41568;
    wire N__41565;
    wire N__41560;
    wire N__41551;
    wire N__41538;
    wire N__41535;
    wire N__41532;
    wire N__41531;
    wire N__41530;
    wire N__41527;
    wire N__41522;
    wire N__41517;
    wire N__41514;
    wire N__41511;
    wire N__41508;
    wire N__41505;
    wire N__41502;
    wire N__41501;
    wire N__41498;
    wire N__41497;
    wire N__41494;
    wire N__41491;
    wire N__41488;
    wire N__41485;
    wire N__41478;
    wire N__41475;
    wire N__41472;
    wire N__41469;
    wire N__41466;
    wire N__41463;
    wire N__41460;
    wire N__41457;
    wire N__41456;
    wire N__41455;
    wire N__41452;
    wire N__41449;
    wire N__41446;
    wire N__41439;
    wire N__41438;
    wire N__41435;
    wire N__41432;
    wire N__41427;
    wire N__41424;
    wire N__41421;
    wire N__41418;
    wire N__41417;
    wire N__41414;
    wire N__41411;
    wire N__41406;
    wire N__41403;
    wire N__41400;
    wire N__41397;
    wire N__41394;
    wire N__41391;
    wire N__41388;
    wire N__41385;
    wire N__41382;
    wire N__41379;
    wire N__41376;
    wire N__41373;
    wire N__41370;
    wire N__41369;
    wire N__41366;
    wire N__41363;
    wire N__41360;
    wire N__41357;
    wire N__41354;
    wire N__41351;
    wire N__41348;
    wire N__41345;
    wire N__41342;
    wire N__41339;
    wire N__41336;
    wire N__41333;
    wire N__41330;
    wire N__41327;
    wire N__41324;
    wire N__41321;
    wire N__41318;
    wire N__41315;
    wire N__41312;
    wire N__41307;
    wire N__41304;
    wire N__41303;
    wire N__41300;
    wire N__41297;
    wire N__41296;
    wire N__41293;
    wire N__41290;
    wire N__41287;
    wire N__41284;
    wire N__41281;
    wire N__41278;
    wire N__41275;
    wire N__41272;
    wire N__41265;
    wire N__41262;
    wire N__41259;
    wire N__41256;
    wire N__41253;
    wire N__41250;
    wire N__41247;
    wire N__41244;
    wire N__41241;
    wire N__41238;
    wire N__41237;
    wire N__41234;
    wire N__41231;
    wire N__41228;
    wire N__41223;
    wire N__41220;
    wire N__41219;
    wire N__41216;
    wire N__41215;
    wire N__41212;
    wire N__41209;
    wire N__41206;
    wire N__41199;
    wire N__41196;
    wire N__41193;
    wire N__41192;
    wire N__41189;
    wire N__41188;
    wire N__41185;
    wire N__41182;
    wire N__41179;
    wire N__41172;
    wire N__41169;
    wire N__41166;
    wire N__41163;
    wire N__41162;
    wire N__41161;
    wire N__41158;
    wire N__41153;
    wire N__41148;
    wire N__41145;
    wire N__41142;
    wire N__41141;
    wire N__41140;
    wire N__41137;
    wire N__41134;
    wire N__41131;
    wire N__41124;
    wire N__41123;
    wire N__41122;
    wire N__41121;
    wire N__41120;
    wire N__41119;
    wire N__41116;
    wire N__41113;
    wire N__41108;
    wire N__41103;
    wire N__41102;
    wire N__41101;
    wire N__41100;
    wire N__41097;
    wire N__41096;
    wire N__41093;
    wire N__41088;
    wire N__41085;
    wire N__41080;
    wire N__41079;
    wire N__41076;
    wire N__41073;
    wire N__41064;
    wire N__41061;
    wire N__41052;
    wire N__41049;
    wire N__41046;
    wire N__41045;
    wire N__41040;
    wire N__41037;
    wire N__41034;
    wire N__41031;
    wire N__41028;
    wire N__41025;
    wire N__41022;
    wire N__41019;
    wire N__41016;
    wire N__41013;
    wire N__41010;
    wire N__41007;
    wire N__41004;
    wire N__41001;
    wire N__40998;
    wire N__40995;
    wire N__40994;
    wire N__40991;
    wire N__40988;
    wire N__40985;
    wire N__40982;
    wire N__40979;
    wire N__40976;
    wire N__40973;
    wire N__40970;
    wire N__40967;
    wire N__40964;
    wire N__40961;
    wire N__40958;
    wire N__40955;
    wire N__40952;
    wire N__40949;
    wire N__40946;
    wire N__40943;
    wire N__40940;
    wire N__40937;
    wire N__40932;
    wire N__40929;
    wire N__40926;
    wire N__40925;
    wire N__40922;
    wire N__40919;
    wire N__40916;
    wire N__40913;
    wire N__40910;
    wire N__40905;
    wire N__40902;
    wire N__40901;
    wire N__40898;
    wire N__40897;
    wire N__40894;
    wire N__40891;
    wire N__40888;
    wire N__40881;
    wire N__40878;
    wire N__40875;
    wire N__40872;
    wire N__40869;
    wire N__40866;
    wire N__40863;
    wire N__40860;
    wire N__40857;
    wire N__40854;
    wire N__40851;
    wire N__40848;
    wire N__40845;
    wire N__40842;
    wire N__40839;
    wire N__40836;
    wire N__40833;
    wire N__40830;
    wire N__40827;
    wire N__40824;
    wire N__40821;
    wire N__40818;
    wire N__40815;
    wire N__40812;
    wire N__40809;
    wire N__40806;
    wire N__40805;
    wire N__40802;
    wire N__40799;
    wire N__40794;
    wire N__40791;
    wire N__40788;
    wire N__40785;
    wire N__40782;
    wire N__40779;
    wire N__40776;
    wire N__40773;
    wire N__40770;
    wire N__40767;
    wire N__40764;
    wire N__40761;
    wire N__40758;
    wire N__40755;
    wire N__40752;
    wire N__40749;
    wire N__40746;
    wire N__40743;
    wire N__40740;
    wire N__40737;
    wire N__40734;
    wire N__40731;
    wire N__40728;
    wire N__40725;
    wire N__40722;
    wire N__40719;
    wire N__40716;
    wire N__40713;
    wire N__40710;
    wire N__40707;
    wire N__40704;
    wire N__40703;
    wire N__40700;
    wire N__40697;
    wire N__40694;
    wire N__40691;
    wire N__40688;
    wire N__40683;
    wire N__40682;
    wire N__40679;
    wire N__40678;
    wire N__40675;
    wire N__40672;
    wire N__40669;
    wire N__40666;
    wire N__40663;
    wire N__40656;
    wire N__40653;
    wire N__40650;
    wire N__40647;
    wire N__40644;
    wire N__40641;
    wire N__40638;
    wire N__40635;
    wire N__40632;
    wire N__40629;
    wire N__40626;
    wire N__40623;
    wire N__40622;
    wire N__40621;
    wire N__40618;
    wire N__40617;
    wire N__40616;
    wire N__40615;
    wire N__40614;
    wire N__40613;
    wire N__40612;
    wire N__40611;
    wire N__40610;
    wire N__40609;
    wire N__40608;
    wire N__40607;
    wire N__40604;
    wire N__40601;
    wire N__40598;
    wire N__40595;
    wire N__40592;
    wire N__40589;
    wire N__40586;
    wire N__40583;
    wire N__40582;
    wire N__40579;
    wire N__40576;
    wire N__40573;
    wire N__40570;
    wire N__40569;
    wire N__40566;
    wire N__40563;
    wire N__40558;
    wire N__40555;
    wire N__40550;
    wire N__40547;
    wire N__40542;
    wire N__40539;
    wire N__40538;
    wire N__40535;
    wire N__40530;
    wire N__40527;
    wire N__40524;
    wire N__40519;
    wire N__40516;
    wire N__40505;
    wire N__40502;
    wire N__40497;
    wire N__40492;
    wire N__40485;
    wire N__40482;
    wire N__40477;
    wire N__40474;
    wire N__40473;
    wire N__40470;
    wire N__40467;
    wire N__40464;
    wire N__40461;
    wire N__40452;
    wire N__40449;
    wire N__40448;
    wire N__40447;
    wire N__40444;
    wire N__40441;
    wire N__40438;
    wire N__40435;
    wire N__40430;
    wire N__40427;
    wire N__40422;
    wire N__40419;
    wire N__40416;
    wire N__40413;
    wire N__40410;
    wire N__40407;
    wire N__40404;
    wire N__40401;
    wire N__40398;
    wire N__40395;
    wire N__40392;
    wire N__40389;
    wire N__40386;
    wire N__40383;
    wire N__40380;
    wire N__40379;
    wire N__40376;
    wire N__40373;
    wire N__40370;
    wire N__40367;
    wire N__40364;
    wire N__40359;
    wire N__40358;
    wire N__40355;
    wire N__40352;
    wire N__40347;
    wire N__40344;
    wire N__40343;
    wire N__40340;
    wire N__40337;
    wire N__40332;
    wire N__40329;
    wire N__40328;
    wire N__40327;
    wire N__40326;
    wire N__40325;
    wire N__40324;
    wire N__40323;
    wire N__40322;
    wire N__40321;
    wire N__40320;
    wire N__40319;
    wire N__40318;
    wire N__40317;
    wire N__40316;
    wire N__40315;
    wire N__40314;
    wire N__40313;
    wire N__40312;
    wire N__40311;
    wire N__40310;
    wire N__40309;
    wire N__40308;
    wire N__40307;
    wire N__40306;
    wire N__40305;
    wire N__40296;
    wire N__40293;
    wire N__40284;
    wire N__40275;
    wire N__40266;
    wire N__40257;
    wire N__40248;
    wire N__40243;
    wire N__40230;
    wire N__40227;
    wire N__40226;
    wire N__40223;
    wire N__40220;
    wire N__40217;
    wire N__40212;
    wire N__40211;
    wire N__40208;
    wire N__40205;
    wire N__40200;
    wire N__40197;
    wire N__40194;
    wire N__40193;
    wire N__40190;
    wire N__40187;
    wire N__40182;
    wire N__40179;
    wire N__40178;
    wire N__40175;
    wire N__40172;
    wire N__40167;
    wire N__40164;
    wire N__40163;
    wire N__40160;
    wire N__40157;
    wire N__40152;
    wire N__40149;
    wire N__40148;
    wire N__40145;
    wire N__40142;
    wire N__40139;
    wire N__40134;
    wire N__40131;
    wire N__40130;
    wire N__40127;
    wire N__40124;
    wire N__40121;
    wire N__40116;
    wire N__40113;
    wire N__40112;
    wire N__40109;
    wire N__40106;
    wire N__40103;
    wire N__40098;
    wire N__40095;
    wire N__40094;
    wire N__40091;
    wire N__40088;
    wire N__40083;
    wire N__40080;
    wire N__40077;
    wire N__40074;
    wire N__40073;
    wire N__40070;
    wire N__40067;
    wire N__40064;
    wire N__40059;
    wire N__40056;
    wire N__40055;
    wire N__40052;
    wire N__40049;
    wire N__40046;
    wire N__40041;
    wire N__40038;
    wire N__40035;
    wire N__40034;
    wire N__40031;
    wire N__40028;
    wire N__40025;
    wire N__40020;
    wire N__40017;
    wire N__40016;
    wire N__40013;
    wire N__40010;
    wire N__40005;
    wire N__40002;
    wire N__39999;
    wire N__39998;
    wire N__39995;
    wire N__39992;
    wire N__39989;
    wire N__39984;
    wire N__39981;
    wire N__39980;
    wire N__39977;
    wire N__39974;
    wire N__39969;
    wire N__39966;
    wire N__39963;
    wire N__39962;
    wire N__39959;
    wire N__39956;
    wire N__39953;
    wire N__39948;
    wire N__39945;
    wire N__39944;
    wire N__39941;
    wire N__39938;
    wire N__39933;
    wire N__39930;
    wire N__39929;
    wire N__39926;
    wire N__39923;
    wire N__39918;
    wire N__39915;
    wire N__39914;
    wire N__39909;
    wire N__39906;
    wire N__39903;
    wire N__39900;
    wire N__39897;
    wire N__39894;
    wire N__39891;
    wire N__39888;
    wire N__39885;
    wire N__39882;
    wire N__39879;
    wire N__39876;
    wire N__39873;
    wire N__39870;
    wire N__39867;
    wire N__39864;
    wire N__39863;
    wire N__39860;
    wire N__39857;
    wire N__39854;
    wire N__39851;
    wire N__39848;
    wire N__39845;
    wire N__39842;
    wire N__39839;
    wire N__39836;
    wire N__39833;
    wire N__39830;
    wire N__39827;
    wire N__39824;
    wire N__39821;
    wire N__39818;
    wire N__39813;
    wire N__39812;
    wire N__39809;
    wire N__39806;
    wire N__39803;
    wire N__39798;
    wire N__39797;
    wire N__39794;
    wire N__39791;
    wire N__39786;
    wire N__39785;
    wire N__39782;
    wire N__39779;
    wire N__39774;
    wire N__39771;
    wire N__39768;
    wire N__39765;
    wire N__39762;
    wire N__39759;
    wire N__39758;
    wire N__39755;
    wire N__39752;
    wire N__39747;
    wire N__39744;
    wire N__39741;
    wire N__39740;
    wire N__39737;
    wire N__39734;
    wire N__39731;
    wire N__39726;
    wire N__39723;
    wire N__39722;
    wire N__39719;
    wire N__39716;
    wire N__39711;
    wire N__39708;
    wire N__39707;
    wire N__39704;
    wire N__39701;
    wire N__39696;
    wire N__39693;
    wire N__39692;
    wire N__39689;
    wire N__39686;
    wire N__39681;
    wire N__39678;
    wire N__39677;
    wire N__39674;
    wire N__39671;
    wire N__39666;
    wire N__39663;
    wire N__39662;
    wire N__39659;
    wire N__39656;
    wire N__39653;
    wire N__39650;
    wire N__39649;
    wire N__39646;
    wire N__39643;
    wire N__39642;
    wire N__39641;
    wire N__39640;
    wire N__39639;
    wire N__39636;
    wire N__39631;
    wire N__39628;
    wire N__39625;
    wire N__39622;
    wire N__39619;
    wire N__39616;
    wire N__39613;
    wire N__39600;
    wire N__39597;
    wire N__39596;
    wire N__39595;
    wire N__39592;
    wire N__39589;
    wire N__39586;
    wire N__39585;
    wire N__39582;
    wire N__39579;
    wire N__39574;
    wire N__39567;
    wire N__39564;
    wire N__39563;
    wire N__39560;
    wire N__39557;
    wire N__39554;
    wire N__39551;
    wire N__39548;
    wire N__39543;
    wire N__39540;
    wire N__39539;
    wire N__39538;
    wire N__39535;
    wire N__39532;
    wire N__39529;
    wire N__39528;
    wire N__39525;
    wire N__39520;
    wire N__39517;
    wire N__39516;
    wire N__39515;
    wire N__39514;
    wire N__39509;
    wire N__39506;
    wire N__39503;
    wire N__39498;
    wire N__39495;
    wire N__39490;
    wire N__39487;
    wire N__39484;
    wire N__39479;
    wire N__39474;
    wire N__39471;
    wire N__39468;
    wire N__39465;
    wire N__39462;
    wire N__39461;
    wire N__39460;
    wire N__39457;
    wire N__39454;
    wire N__39451;
    wire N__39444;
    wire N__39441;
    wire N__39438;
    wire N__39435;
    wire N__39432;
    wire N__39429;
    wire N__39426;
    wire N__39423;
    wire N__39420;
    wire N__39417;
    wire N__39414;
    wire N__39411;
    wire N__39408;
    wire N__39405;
    wire N__39402;
    wire N__39401;
    wire N__39398;
    wire N__39395;
    wire N__39392;
    wire N__39389;
    wire N__39386;
    wire N__39383;
    wire N__39380;
    wire N__39377;
    wire N__39374;
    wire N__39371;
    wire N__39368;
    wire N__39365;
    wire N__39362;
    wire N__39357;
    wire N__39356;
    wire N__39355;
    wire N__39352;
    wire N__39349;
    wire N__39346;
    wire N__39341;
    wire N__39336;
    wire N__39333;
    wire N__39330;
    wire N__39327;
    wire N__39326;
    wire N__39323;
    wire N__39320;
    wire N__39315;
    wire N__39312;
    wire N__39309;
    wire N__39306;
    wire N__39303;
    wire N__39300;
    wire N__39297;
    wire N__39294;
    wire N__39291;
    wire N__39288;
    wire N__39285;
    wire N__39282;
    wire N__39279;
    wire N__39276;
    wire N__39273;
    wire N__39272;
    wire N__39269;
    wire N__39266;
    wire N__39263;
    wire N__39260;
    wire N__39257;
    wire N__39254;
    wire N__39251;
    wire N__39248;
    wire N__39245;
    wire N__39242;
    wire N__39239;
    wire N__39236;
    wire N__39233;
    wire N__39230;
    wire N__39227;
    wire N__39222;
    wire N__39221;
    wire N__39218;
    wire N__39215;
    wire N__39214;
    wire N__39209;
    wire N__39206;
    wire N__39203;
    wire N__39198;
    wire N__39197;
    wire N__39192;
    wire N__39189;
    wire N__39188;
    wire N__39183;
    wire N__39180;
    wire N__39177;
    wire N__39176;
    wire N__39173;
    wire N__39170;
    wire N__39169;
    wire N__39166;
    wire N__39163;
    wire N__39160;
    wire N__39155;
    wire N__39150;
    wire N__39147;
    wire N__39144;
    wire N__39143;
    wire N__39142;
    wire N__39139;
    wire N__39136;
    wire N__39133;
    wire N__39130;
    wire N__39127;
    wire N__39124;
    wire N__39121;
    wire N__39118;
    wire N__39111;
    wire N__39108;
    wire N__39105;
    wire N__39104;
    wire N__39103;
    wire N__39100;
    wire N__39097;
    wire N__39094;
    wire N__39091;
    wire N__39084;
    wire N__39081;
    wire N__39078;
    wire N__39077;
    wire N__39076;
    wire N__39073;
    wire N__39070;
    wire N__39067;
    wire N__39062;
    wire N__39057;
    wire N__39056;
    wire N__39055;
    wire N__39052;
    wire N__39049;
    wire N__39046;
    wire N__39041;
    wire N__39036;
    wire N__39033;
    wire N__39030;
    wire N__39027;
    wire N__39026;
    wire N__39023;
    wire N__39020;
    wire N__39017;
    wire N__39014;
    wire N__39009;
    wire N__39006;
    wire N__39005;
    wire N__39002;
    wire N__38999;
    wire N__38996;
    wire N__38993;
    wire N__38988;
    wire N__38985;
    wire N__38982;
    wire N__38979;
    wire N__38976;
    wire N__38975;
    wire N__38972;
    wire N__38969;
    wire N__38964;
    wire N__38963;
    wire N__38962;
    wire N__38959;
    wire N__38956;
    wire N__38953;
    wire N__38946;
    wire N__38945;
    wire N__38944;
    wire N__38941;
    wire N__38938;
    wire N__38935;
    wire N__38934;
    wire N__38933;
    wire N__38932;
    wire N__38931;
    wire N__38930;
    wire N__38929;
    wire N__38928;
    wire N__38927;
    wire N__38924;
    wire N__38921;
    wire N__38918;
    wire N__38915;
    wire N__38912;
    wire N__38909;
    wire N__38906;
    wire N__38903;
    wire N__38900;
    wire N__38897;
    wire N__38894;
    wire N__38891;
    wire N__38886;
    wire N__38877;
    wire N__38868;
    wire N__38859;
    wire N__38856;
    wire N__38853;
    wire N__38850;
    wire N__38847;
    wire N__38844;
    wire N__38841;
    wire N__38838;
    wire N__38835;
    wire N__38832;
    wire N__38829;
    wire N__38828;
    wire N__38825;
    wire N__38824;
    wire N__38821;
    wire N__38814;
    wire N__38811;
    wire N__38810;
    wire N__38807;
    wire N__38804;
    wire N__38801;
    wire N__38798;
    wire N__38795;
    wire N__38790;
    wire N__38789;
    wire N__38788;
    wire N__38785;
    wire N__38780;
    wire N__38775;
    wire N__38774;
    wire N__38773;
    wire N__38772;
    wire N__38771;
    wire N__38770;
    wire N__38765;
    wire N__38764;
    wire N__38763;
    wire N__38762;
    wire N__38759;
    wire N__38754;
    wire N__38753;
    wire N__38752;
    wire N__38751;
    wire N__38750;
    wire N__38749;
    wire N__38748;
    wire N__38747;
    wire N__38746;
    wire N__38745;
    wire N__38744;
    wire N__38743;
    wire N__38742;
    wire N__38739;
    wire N__38738;
    wire N__38737;
    wire N__38734;
    wire N__38731;
    wire N__38728;
    wire N__38725;
    wire N__38722;
    wire N__38719;
    wire N__38712;
    wire N__38709;
    wire N__38706;
    wire N__38701;
    wire N__38696;
    wire N__38693;
    wire N__38688;
    wire N__38685;
    wire N__38680;
    wire N__38673;
    wire N__38670;
    wire N__38665;
    wire N__38662;
    wire N__38659;
    wire N__38654;
    wire N__38651;
    wire N__38644;
    wire N__38641;
    wire N__38640;
    wire N__38635;
    wire N__38628;
    wire N__38619;
    wire N__38616;
    wire N__38607;
    wire N__38606;
    wire N__38603;
    wire N__38602;
    wire N__38601;
    wire N__38600;
    wire N__38599;
    wire N__38598;
    wire N__38597;
    wire N__38596;
    wire N__38595;
    wire N__38594;
    wire N__38593;
    wire N__38592;
    wire N__38591;
    wire N__38590;
    wire N__38589;
    wire N__38588;
    wire N__38587;
    wire N__38586;
    wire N__38585;
    wire N__38584;
    wire N__38583;
    wire N__38582;
    wire N__38579;
    wire N__38574;
    wire N__38571;
    wire N__38570;
    wire N__38565;
    wire N__38564;
    wire N__38563;
    wire N__38562;
    wire N__38561;
    wire N__38560;
    wire N__38559;
    wire N__38558;
    wire N__38557;
    wire N__38554;
    wire N__38553;
    wire N__38552;
    wire N__38551;
    wire N__38544;
    wire N__38533;
    wire N__38528;
    wire N__38515;
    wire N__38510;
    wire N__38507;
    wire N__38506;
    wire N__38505;
    wire N__38504;
    wire N__38503;
    wire N__38502;
    wire N__38501;
    wire N__38500;
    wire N__38497;
    wire N__38494;
    wire N__38491;
    wire N__38488;
    wire N__38481;
    wire N__38474;
    wire N__38471;
    wire N__38468;
    wire N__38463;
    wire N__38460;
    wire N__38459;
    wire N__38458;
    wire N__38457;
    wire N__38456;
    wire N__38455;
    wire N__38454;
    wire N__38453;
    wire N__38452;
    wire N__38451;
    wire N__38450;
    wire N__38449;
    wire N__38448;
    wire N__38447;
    wire N__38446;
    wire N__38443;
    wire N__38438;
    wire N__38435;
    wire N__38432;
    wire N__38427;
    wire N__38422;
    wire N__38415;
    wire N__38412;
    wire N__38409;
    wire N__38408;
    wire N__38407;
    wire N__38406;
    wire N__38405;
    wire N__38404;
    wire N__38403;
    wire N__38402;
    wire N__38401;
    wire N__38400;
    wire N__38399;
    wire N__38398;
    wire N__38397;
    wire N__38394;
    wire N__38385;
    wire N__38378;
    wire N__38371;
    wire N__38364;
    wire N__38353;
    wire N__38348;
    wire N__38345;
    wire N__38342;
    wire N__38335;
    wire N__38324;
    wire N__38317;
    wire N__38308;
    wire N__38297;
    wire N__38288;
    wire N__38265;
    wire N__38264;
    wire N__38263;
    wire N__38260;
    wire N__38257;
    wire N__38254;
    wire N__38251;
    wire N__38248;
    wire N__38245;
    wire N__38238;
    wire N__38237;
    wire N__38236;
    wire N__38233;
    wire N__38230;
    wire N__38227;
    wire N__38224;
    wire N__38221;
    wire N__38218;
    wire N__38215;
    wire N__38212;
    wire N__38205;
    wire N__38202;
    wire N__38199;
    wire N__38196;
    wire N__38195;
    wire N__38192;
    wire N__38189;
    wire N__38184;
    wire N__38183;
    wire N__38182;
    wire N__38179;
    wire N__38176;
    wire N__38173;
    wire N__38168;
    wire N__38163;
    wire N__38160;
    wire N__38157;
    wire N__38154;
    wire N__38151;
    wire N__38150;
    wire N__38149;
    wire N__38146;
    wire N__38143;
    wire N__38140;
    wire N__38139;
    wire N__38136;
    wire N__38133;
    wire N__38130;
    wire N__38127;
    wire N__38124;
    wire N__38121;
    wire N__38118;
    wire N__38115;
    wire N__38106;
    wire N__38103;
    wire N__38100;
    wire N__38097;
    wire N__38096;
    wire N__38095;
    wire N__38092;
    wire N__38089;
    wire N__38086;
    wire N__38079;
    wire N__38078;
    wire N__38075;
    wire N__38072;
    wire N__38067;
    wire N__38064;
    wire N__38061;
    wire N__38058;
    wire N__38057;
    wire N__38054;
    wire N__38051;
    wire N__38050;
    wire N__38045;
    wire N__38042;
    wire N__38039;
    wire N__38034;
    wire N__38033;
    wire N__38030;
    wire N__38027;
    wire N__38024;
    wire N__38021;
    wire N__38018;
    wire N__38013;
    wire N__38010;
    wire N__38009;
    wire N__38008;
    wire N__38005;
    wire N__38002;
    wire N__37999;
    wire N__37994;
    wire N__37989;
    wire N__37988;
    wire N__37983;
    wire N__37980;
    wire N__37977;
    wire N__37974;
    wire N__37971;
    wire N__37968;
    wire N__37965;
    wire N__37962;
    wire N__37959;
    wire N__37956;
    wire N__37955;
    wire N__37954;
    wire N__37951;
    wire N__37948;
    wire N__37945;
    wire N__37942;
    wire N__37939;
    wire N__37932;
    wire N__37929;
    wire N__37926;
    wire N__37925;
    wire N__37922;
    wire N__37919;
    wire N__37916;
    wire N__37911;
    wire N__37908;
    wire N__37905;
    wire N__37904;
    wire N__37901;
    wire N__37898;
    wire N__37895;
    wire N__37890;
    wire N__37887;
    wire N__37884;
    wire N__37883;
    wire N__37880;
    wire N__37877;
    wire N__37874;
    wire N__37869;
    wire N__37866;
    wire N__37863;
    wire N__37860;
    wire N__37859;
    wire N__37856;
    wire N__37853;
    wire N__37850;
    wire N__37845;
    wire N__37844;
    wire N__37843;
    wire N__37842;
    wire N__37839;
    wire N__37836;
    wire N__37833;
    wire N__37830;
    wire N__37827;
    wire N__37824;
    wire N__37821;
    wire N__37818;
    wire N__37815;
    wire N__37812;
    wire N__37809;
    wire N__37808;
    wire N__37805;
    wire N__37802;
    wire N__37797;
    wire N__37794;
    wire N__37785;
    wire N__37784;
    wire N__37781;
    wire N__37780;
    wire N__37779;
    wire N__37776;
    wire N__37773;
    wire N__37772;
    wire N__37771;
    wire N__37766;
    wire N__37763;
    wire N__37760;
    wire N__37757;
    wire N__37754;
    wire N__37751;
    wire N__37748;
    wire N__37743;
    wire N__37736;
    wire N__37733;
    wire N__37728;
    wire N__37725;
    wire N__37722;
    wire N__37721;
    wire N__37718;
    wire N__37717;
    wire N__37714;
    wire N__37711;
    wire N__37708;
    wire N__37701;
    wire N__37698;
    wire N__37695;
    wire N__37692;
    wire N__37691;
    wire N__37690;
    wire N__37687;
    wire N__37684;
    wire N__37681;
    wire N__37678;
    wire N__37671;
    wire N__37668;
    wire N__37667;
    wire N__37664;
    wire N__37661;
    wire N__37660;
    wire N__37657;
    wire N__37654;
    wire N__37651;
    wire N__37648;
    wire N__37645;
    wire N__37638;
    wire N__37635;
    wire N__37632;
    wire N__37629;
    wire N__37626;
    wire N__37623;
    wire N__37620;
    wire N__37617;
    wire N__37614;
    wire N__37611;
    wire N__37608;
    wire N__37605;
    wire N__37602;
    wire N__37599;
    wire N__37596;
    wire N__37593;
    wire N__37590;
    wire N__37589;
    wire N__37586;
    wire N__37583;
    wire N__37582;
    wire N__37579;
    wire N__37576;
    wire N__37573;
    wire N__37572;
    wire N__37571;
    wire N__37570;
    wire N__37567;
    wire N__37564;
    wire N__37557;
    wire N__37554;
    wire N__37545;
    wire N__37542;
    wire N__37539;
    wire N__37536;
    wire N__37533;
    wire N__37532;
    wire N__37531;
    wire N__37528;
    wire N__37525;
    wire N__37524;
    wire N__37523;
    wire N__37522;
    wire N__37519;
    wire N__37514;
    wire N__37509;
    wire N__37506;
    wire N__37503;
    wire N__37498;
    wire N__37497;
    wire N__37496;
    wire N__37493;
    wire N__37488;
    wire N__37483;
    wire N__37476;
    wire N__37473;
    wire N__37472;
    wire N__37469;
    wire N__37466;
    wire N__37461;
    wire N__37458;
    wire N__37455;
    wire N__37452;
    wire N__37449;
    wire N__37446;
    wire N__37445;
    wire N__37442;
    wire N__37439;
    wire N__37436;
    wire N__37431;
    wire N__37428;
    wire N__37425;
    wire N__37422;
    wire N__37419;
    wire N__37416;
    wire N__37413;
    wire N__37410;
    wire N__37407;
    wire N__37404;
    wire N__37401;
    wire N__37398;
    wire N__37395;
    wire N__37392;
    wire N__37389;
    wire N__37386;
    wire N__37383;
    wire N__37380;
    wire N__37377;
    wire N__37374;
    wire N__37371;
    wire N__37368;
    wire N__37365;
    wire N__37362;
    wire N__37359;
    wire N__37356;
    wire N__37353;
    wire N__37350;
    wire N__37347;
    wire N__37344;
    wire N__37341;
    wire N__37338;
    wire N__37335;
    wire N__37332;
    wire N__37329;
    wire N__37326;
    wire N__37323;
    wire N__37320;
    wire N__37317;
    wire N__37314;
    wire N__37313;
    wire N__37312;
    wire N__37311;
    wire N__37304;
    wire N__37301;
    wire N__37296;
    wire N__37295;
    wire N__37294;
    wire N__37289;
    wire N__37286;
    wire N__37281;
    wire N__37278;
    wire N__37277;
    wire N__37276;
    wire N__37275;
    wire N__37274;
    wire N__37265;
    wire N__37262;
    wire N__37257;
    wire N__37254;
    wire N__37251;
    wire N__37250;
    wire N__37249;
    wire N__37246;
    wire N__37243;
    wire N__37240;
    wire N__37237;
    wire N__37234;
    wire N__37231;
    wire N__37228;
    wire N__37225;
    wire N__37222;
    wire N__37219;
    wire N__37216;
    wire N__37213;
    wire N__37206;
    wire N__37203;
    wire N__37200;
    wire N__37197;
    wire N__37196;
    wire N__37193;
    wire N__37190;
    wire N__37187;
    wire N__37182;
    wire N__37179;
    wire N__37176;
    wire N__37173;
    wire N__37170;
    wire N__37167;
    wire N__37164;
    wire N__37161;
    wire N__37158;
    wire N__37155;
    wire N__37152;
    wire N__37149;
    wire N__37146;
    wire N__37143;
    wire N__37140;
    wire N__37137;
    wire N__37134;
    wire N__37131;
    wire N__37128;
    wire N__37125;
    wire N__37122;
    wire N__37119;
    wire N__37116;
    wire N__37113;
    wire N__37110;
    wire N__37109;
    wire N__37106;
    wire N__37103;
    wire N__37100;
    wire N__37095;
    wire N__37092;
    wire N__37089;
    wire N__37086;
    wire N__37085;
    wire N__37082;
    wire N__37079;
    wire N__37076;
    wire N__37071;
    wire N__37068;
    wire N__37065;
    wire N__37062;
    wire N__37059;
    wire N__37058;
    wire N__37055;
    wire N__37052;
    wire N__37049;
    wire N__37044;
    wire N__37043;
    wire N__37042;
    wire N__37039;
    wire N__37036;
    wire N__37035;
    wire N__37032;
    wire N__37027;
    wire N__37024;
    wire N__37021;
    wire N__37018;
    wire N__37015;
    wire N__37010;
    wire N__37007;
    wire N__37002;
    wire N__36999;
    wire N__36998;
    wire N__36995;
    wire N__36992;
    wire N__36989;
    wire N__36986;
    wire N__36983;
    wire N__36980;
    wire N__36977;
    wire N__36972;
    wire N__36971;
    wire N__36970;
    wire N__36967;
    wire N__36964;
    wire N__36961;
    wire N__36954;
    wire N__36951;
    wire N__36950;
    wire N__36947;
    wire N__36944;
    wire N__36939;
    wire N__36936;
    wire N__36933;
    wire N__36930;
    wire N__36929;
    wire N__36926;
    wire N__36923;
    wire N__36918;
    wire N__36915;
    wire N__36912;
    wire N__36911;
    wire N__36908;
    wire N__36905;
    wire N__36904;
    wire N__36899;
    wire N__36896;
    wire N__36891;
    wire N__36888;
    wire N__36887;
    wire N__36886;
    wire N__36883;
    wire N__36880;
    wire N__36877;
    wire N__36874;
    wire N__36867;
    wire N__36864;
    wire N__36863;
    wire N__36860;
    wire N__36857;
    wire N__36854;
    wire N__36849;
    wire N__36846;
    wire N__36843;
    wire N__36842;
    wire N__36839;
    wire N__36836;
    wire N__36833;
    wire N__36828;
    wire N__36825;
    wire N__36822;
    wire N__36819;
    wire N__36818;
    wire N__36815;
    wire N__36812;
    wire N__36809;
    wire N__36804;
    wire N__36801;
    wire N__36798;
    wire N__36797;
    wire N__36794;
    wire N__36791;
    wire N__36788;
    wire N__36783;
    wire N__36780;
    wire N__36777;
    wire N__36776;
    wire N__36773;
    wire N__36770;
    wire N__36767;
    wire N__36762;
    wire N__36759;
    wire N__36756;
    wire N__36753;
    wire N__36750;
    wire N__36747;
    wire N__36746;
    wire N__36743;
    wire N__36740;
    wire N__36737;
    wire N__36732;
    wire N__36729;
    wire N__36726;
    wire N__36723;
    wire N__36720;
    wire N__36719;
    wire N__36716;
    wire N__36713;
    wire N__36710;
    wire N__36705;
    wire N__36702;
    wire N__36699;
    wire N__36698;
    wire N__36695;
    wire N__36692;
    wire N__36689;
    wire N__36684;
    wire N__36681;
    wire N__36680;
    wire N__36677;
    wire N__36674;
    wire N__36671;
    wire N__36666;
    wire N__36663;
    wire N__36660;
    wire N__36657;
    wire N__36654;
    wire N__36653;
    wire N__36650;
    wire N__36647;
    wire N__36644;
    wire N__36639;
    wire N__36636;
    wire N__36633;
    wire N__36630;
    wire N__36627;
    wire N__36624;
    wire N__36621;
    wire N__36618;
    wire N__36615;
    wire N__36612;
    wire N__36609;
    wire N__36606;
    wire N__36605;
    wire N__36602;
    wire N__36599;
    wire N__36596;
    wire N__36591;
    wire N__36588;
    wire N__36585;
    wire N__36582;
    wire N__36579;
    wire N__36576;
    wire N__36573;
    wire N__36570;
    wire N__36569;
    wire N__36568;
    wire N__36565;
    wire N__36562;
    wire N__36559;
    wire N__36556;
    wire N__36553;
    wire N__36546;
    wire N__36545;
    wire N__36542;
    wire N__36539;
    wire N__36536;
    wire N__36533;
    wire N__36530;
    wire N__36525;
    wire N__36522;
    wire N__36519;
    wire N__36516;
    wire N__36513;
    wire N__36512;
    wire N__36507;
    wire N__36504;
    wire N__36501;
    wire N__36498;
    wire N__36495;
    wire N__36492;
    wire N__36489;
    wire N__36486;
    wire N__36485;
    wire N__36482;
    wire N__36481;
    wire N__36478;
    wire N__36475;
    wire N__36472;
    wire N__36467;
    wire N__36466;
    wire N__36465;
    wire N__36462;
    wire N__36459;
    wire N__36454;
    wire N__36451;
    wire N__36448;
    wire N__36441;
    wire N__36438;
    wire N__36435;
    wire N__36432;
    wire N__36429;
    wire N__36426;
    wire N__36423;
    wire N__36420;
    wire N__36417;
    wire N__36414;
    wire N__36411;
    wire N__36408;
    wire N__36405;
    wire N__36402;
    wire N__36399;
    wire N__36396;
    wire N__36393;
    wire N__36392;
    wire N__36389;
    wire N__36386;
    wire N__36383;
    wire N__36380;
    wire N__36377;
    wire N__36374;
    wire N__36371;
    wire N__36368;
    wire N__36365;
    wire N__36362;
    wire N__36359;
    wire N__36354;
    wire N__36351;
    wire N__36348;
    wire N__36345;
    wire N__36344;
    wire N__36341;
    wire N__36338;
    wire N__36335;
    wire N__36332;
    wire N__36331;
    wire N__36328;
    wire N__36325;
    wire N__36322;
    wire N__36315;
    wire N__36312;
    wire N__36309;
    wire N__36306;
    wire N__36303;
    wire N__36302;
    wire N__36301;
    wire N__36298;
    wire N__36293;
    wire N__36288;
    wire N__36287;
    wire N__36284;
    wire N__36281;
    wire N__36278;
    wire N__36277;
    wire N__36274;
    wire N__36271;
    wire N__36268;
    wire N__36263;
    wire N__36258;
    wire N__36257;
    wire N__36256;
    wire N__36253;
    wire N__36250;
    wire N__36247;
    wire N__36244;
    wire N__36237;
    wire N__36234;
    wire N__36231;
    wire N__36228;
    wire N__36225;
    wire N__36222;
    wire N__36219;
    wire N__36216;
    wire N__36215;
    wire N__36214;
    wire N__36211;
    wire N__36208;
    wire N__36205;
    wire N__36198;
    wire N__36197;
    wire N__36196;
    wire N__36193;
    wire N__36190;
    wire N__36187;
    wire N__36182;
    wire N__36179;
    wire N__36176;
    wire N__36171;
    wire N__36170;
    wire N__36167;
    wire N__36166;
    wire N__36165;
    wire N__36162;
    wire N__36159;
    wire N__36156;
    wire N__36153;
    wire N__36150;
    wire N__36147;
    wire N__36144;
    wire N__36139;
    wire N__36136;
    wire N__36129;
    wire N__36128;
    wire N__36125;
    wire N__36122;
    wire N__36117;
    wire N__36114;
    wire N__36111;
    wire N__36108;
    wire N__36105;
    wire N__36102;
    wire N__36099;
    wire N__36096;
    wire N__36093;
    wire N__36090;
    wire N__36087;
    wire N__36084;
    wire N__36081;
    wire N__36080;
    wire N__36077;
    wire N__36074;
    wire N__36071;
    wire N__36068;
    wire N__36065;
    wire N__36062;
    wire N__36059;
    wire N__36056;
    wire N__36053;
    wire N__36050;
    wire N__36047;
    wire N__36044;
    wire N__36041;
    wire N__36038;
    wire N__36035;
    wire N__36032;
    wire N__36029;
    wire N__36024;
    wire N__36021;
    wire N__36018;
    wire N__36015;
    wire N__36012;
    wire N__36009;
    wire N__36006;
    wire N__36003;
    wire N__36000;
    wire N__35997;
    wire N__35996;
    wire N__35993;
    wire N__35990;
    wire N__35989;
    wire N__35984;
    wire N__35981;
    wire N__35978;
    wire N__35975;
    wire N__35972;
    wire N__35967;
    wire N__35964;
    wire N__35961;
    wire N__35958;
    wire N__35955;
    wire N__35952;
    wire N__35949;
    wire N__35946;
    wire N__35943;
    wire N__35940;
    wire N__35937;
    wire N__35934;
    wire N__35931;
    wire N__35928;
    wire N__35925;
    wire N__35922;
    wire N__35921;
    wire N__35918;
    wire N__35915;
    wire N__35912;
    wire N__35909;
    wire N__35906;
    wire N__35903;
    wire N__35900;
    wire N__35897;
    wire N__35894;
    wire N__35891;
    wire N__35888;
    wire N__35883;
    wire N__35880;
    wire N__35877;
    wire N__35876;
    wire N__35875;
    wire N__35874;
    wire N__35873;
    wire N__35872;
    wire N__35871;
    wire N__35870;
    wire N__35867;
    wire N__35866;
    wire N__35865;
    wire N__35862;
    wire N__35861;
    wire N__35860;
    wire N__35859;
    wire N__35852;
    wire N__35847;
    wire N__35844;
    wire N__35841;
    wire N__35834;
    wire N__35829;
    wire N__35826;
    wire N__35811;
    wire N__35808;
    wire N__35807;
    wire N__35804;
    wire N__35801;
    wire N__35800;
    wire N__35795;
    wire N__35794;
    wire N__35793;
    wire N__35792;
    wire N__35791;
    wire N__35788;
    wire N__35785;
    wire N__35784;
    wire N__35783;
    wire N__35782;
    wire N__35781;
    wire N__35778;
    wire N__35777;
    wire N__35776;
    wire N__35775;
    wire N__35768;
    wire N__35763;
    wire N__35752;
    wire N__35745;
    wire N__35736;
    wire N__35735;
    wire N__35734;
    wire N__35733;
    wire N__35732;
    wire N__35731;
    wire N__35728;
    wire N__35725;
    wire N__35720;
    wire N__35717;
    wire N__35714;
    wire N__35711;
    wire N__35710;
    wire N__35709;
    wire N__35708;
    wire N__35707;
    wire N__35706;
    wire N__35703;
    wire N__35698;
    wire N__35695;
    wire N__35692;
    wire N__35689;
    wire N__35686;
    wire N__35681;
    wire N__35678;
    wire N__35675;
    wire N__35672;
    wire N__35667;
    wire N__35664;
    wire N__35661;
    wire N__35658;
    wire N__35643;
    wire N__35640;
    wire N__35637;
    wire N__35634;
    wire N__35631;
    wire N__35630;
    wire N__35629;
    wire N__35626;
    wire N__35623;
    wire N__35620;
    wire N__35617;
    wire N__35614;
    wire N__35607;
    wire N__35604;
    wire N__35603;
    wire N__35602;
    wire N__35599;
    wire N__35596;
    wire N__35593;
    wire N__35590;
    wire N__35587;
    wire N__35584;
    wire N__35581;
    wire N__35578;
    wire N__35571;
    wire N__35570;
    wire N__35569;
    wire N__35562;
    wire N__35561;
    wire N__35560;
    wire N__35559;
    wire N__35558;
    wire N__35557;
    wire N__35556;
    wire N__35555;
    wire N__35552;
    wire N__35547;
    wire N__35544;
    wire N__35539;
    wire N__35538;
    wire N__35537;
    wire N__35534;
    wire N__35533;
    wire N__35530;
    wire N__35525;
    wire N__35520;
    wire N__35511;
    wire N__35510;
    wire N__35509;
    wire N__35508;
    wire N__35505;
    wire N__35502;
    wire N__35499;
    wire N__35496;
    wire N__35489;
    wire N__35478;
    wire N__35475;
    wire N__35472;
    wire N__35469;
    wire N__35466;
    wire N__35463;
    wire N__35460;
    wire N__35457;
    wire N__35456;
    wire N__35453;
    wire N__35450;
    wire N__35445;
    wire N__35442;
    wire N__35439;
    wire N__35436;
    wire N__35433;
    wire N__35430;
    wire N__35427;
    wire N__35424;
    wire N__35423;
    wire N__35420;
    wire N__35417;
    wire N__35414;
    wire N__35411;
    wire N__35408;
    wire N__35403;
    wire N__35400;
    wire N__35397;
    wire N__35394;
    wire N__35393;
    wire N__35392;
    wire N__35389;
    wire N__35384;
    wire N__35379;
    wire N__35376;
    wire N__35375;
    wire N__35374;
    wire N__35371;
    wire N__35368;
    wire N__35365;
    wire N__35362;
    wire N__35357;
    wire N__35352;
    wire N__35349;
    wire N__35346;
    wire N__35343;
    wire N__35340;
    wire N__35337;
    wire N__35336;
    wire N__35335;
    wire N__35332;
    wire N__35329;
    wire N__35326;
    wire N__35323;
    wire N__35316;
    wire N__35313;
    wire N__35310;
    wire N__35309;
    wire N__35306;
    wire N__35303;
    wire N__35300;
    wire N__35299;
    wire N__35296;
    wire N__35293;
    wire N__35290;
    wire N__35287;
    wire N__35280;
    wire N__35279;
    wire N__35276;
    wire N__35273;
    wire N__35270;
    wire N__35267;
    wire N__35264;
    wire N__35261;
    wire N__35256;
    wire N__35253;
    wire N__35250;
    wire N__35247;
    wire N__35246;
    wire N__35243;
    wire N__35240;
    wire N__35237;
    wire N__35234;
    wire N__35231;
    wire N__35226;
    wire N__35223;
    wire N__35220;
    wire N__35217;
    wire N__35214;
    wire N__35211;
    wire N__35210;
    wire N__35207;
    wire N__35206;
    wire N__35203;
    wire N__35200;
    wire N__35197;
    wire N__35192;
    wire N__35187;
    wire N__35184;
    wire N__35181;
    wire N__35178;
    wire N__35175;
    wire N__35172;
    wire N__35169;
    wire N__35166;
    wire N__35163;
    wire N__35160;
    wire N__35159;
    wire N__35156;
    wire N__35153;
    wire N__35148;
    wire N__35145;
    wire N__35144;
    wire N__35141;
    wire N__35138;
    wire N__35135;
    wire N__35130;
    wire N__35129;
    wire N__35126;
    wire N__35123;
    wire N__35120;
    wire N__35115;
    wire N__35112;
    wire N__35109;
    wire N__35106;
    wire N__35103;
    wire N__35100;
    wire N__35097;
    wire N__35094;
    wire N__35091;
    wire N__35088;
    wire N__35085;
    wire N__35082;
    wire N__35079;
    wire N__35076;
    wire N__35073;
    wire N__35070;
    wire N__35069;
    wire N__35066;
    wire N__35063;
    wire N__35060;
    wire N__35057;
    wire N__35052;
    wire N__35049;
    wire N__35046;
    wire N__35045;
    wire N__35044;
    wire N__35041;
    wire N__35038;
    wire N__35035;
    wire N__35030;
    wire N__35025;
    wire N__35022;
    wire N__35021;
    wire N__35018;
    wire N__35015;
    wire N__35010;
    wire N__35009;
    wire N__35008;
    wire N__35005;
    wire N__35000;
    wire N__34999;
    wire N__34998;
    wire N__34993;
    wire N__34990;
    wire N__34987;
    wire N__34984;
    wire N__34981;
    wire N__34978;
    wire N__34971;
    wire N__34968;
    wire N__34967;
    wire N__34964;
    wire N__34961;
    wire N__34960;
    wire N__34957;
    wire N__34954;
    wire N__34951;
    wire N__34948;
    wire N__34941;
    wire N__34940;
    wire N__34939;
    wire N__34934;
    wire N__34931;
    wire N__34928;
    wire N__34923;
    wire N__34920;
    wire N__34919;
    wire N__34918;
    wire N__34915;
    wire N__34912;
    wire N__34909;
    wire N__34902;
    wire N__34899;
    wire N__34896;
    wire N__34893;
    wire N__34892;
    wire N__34889;
    wire N__34886;
    wire N__34881;
    wire N__34880;
    wire N__34879;
    wire N__34874;
    wire N__34871;
    wire N__34866;
    wire N__34863;
    wire N__34860;
    wire N__34859;
    wire N__34856;
    wire N__34855;
    wire N__34852;
    wire N__34851;
    wire N__34848;
    wire N__34845;
    wire N__34842;
    wire N__34839;
    wire N__34836;
    wire N__34833;
    wire N__34830;
    wire N__34827;
    wire N__34822;
    wire N__34819;
    wire N__34816;
    wire N__34813;
    wire N__34806;
    wire N__34805;
    wire N__34804;
    wire N__34801;
    wire N__34798;
    wire N__34795;
    wire N__34788;
    wire N__34785;
    wire N__34782;
    wire N__34779;
    wire N__34776;
    wire N__34773;
    wire N__34770;
    wire N__34769;
    wire N__34768;
    wire N__34765;
    wire N__34760;
    wire N__34755;
    wire N__34752;
    wire N__34751;
    wire N__34750;
    wire N__34747;
    wire N__34742;
    wire N__34737;
    wire N__34734;
    wire N__34731;
    wire N__34728;
    wire N__34725;
    wire N__34722;
    wire N__34719;
    wire N__34716;
    wire N__34715;
    wire N__34714;
    wire N__34711;
    wire N__34708;
    wire N__34705;
    wire N__34702;
    wire N__34697;
    wire N__34694;
    wire N__34693;
    wire N__34690;
    wire N__34687;
    wire N__34684;
    wire N__34677;
    wire N__34674;
    wire N__34671;
    wire N__34668;
    wire N__34665;
    wire N__34664;
    wire N__34661;
    wire N__34658;
    wire N__34655;
    wire N__34652;
    wire N__34647;
    wire N__34644;
    wire N__34643;
    wire N__34640;
    wire N__34637;
    wire N__34634;
    wire N__34629;
    wire N__34626;
    wire N__34625;
    wire N__34622;
    wire N__34619;
    wire N__34616;
    wire N__34611;
    wire N__34610;
    wire N__34607;
    wire N__34604;
    wire N__34601;
    wire N__34596;
    wire N__34593;
    wire N__34592;
    wire N__34589;
    wire N__34586;
    wire N__34583;
    wire N__34578;
    wire N__34575;
    wire N__34572;
    wire N__34571;
    wire N__34568;
    wire N__34565;
    wire N__34562;
    wire N__34557;
    wire N__34554;
    wire N__34553;
    wire N__34550;
    wire N__34547;
    wire N__34542;
    wire N__34539;
    wire N__34536;
    wire N__34533;
    wire N__34532;
    wire N__34529;
    wire N__34526;
    wire N__34523;
    wire N__34518;
    wire N__34517;
    wire N__34514;
    wire N__34511;
    wire N__34508;
    wire N__34503;
    wire N__34500;
    wire N__34497;
    wire N__34494;
    wire N__34491;
    wire N__34488;
    wire N__34487;
    wire N__34484;
    wire N__34481;
    wire N__34480;
    wire N__34477;
    wire N__34474;
    wire N__34471;
    wire N__34466;
    wire N__34461;
    wire N__34458;
    wire N__34455;
    wire N__34452;
    wire N__34449;
    wire N__34446;
    wire N__34443;
    wire N__34440;
    wire N__34437;
    wire N__34436;
    wire N__34433;
    wire N__34430;
    wire N__34429;
    wire N__34426;
    wire N__34423;
    wire N__34422;
    wire N__34419;
    wire N__34414;
    wire N__34411;
    wire N__34404;
    wire N__34401;
    wire N__34398;
    wire N__34397;
    wire N__34394;
    wire N__34393;
    wire N__34390;
    wire N__34387;
    wire N__34384;
    wire N__34377;
    wire N__34374;
    wire N__34373;
    wire N__34370;
    wire N__34369;
    wire N__34366;
    wire N__34363;
    wire N__34360;
    wire N__34359;
    wire N__34354;
    wire N__34351;
    wire N__34348;
    wire N__34341;
    wire N__34338;
    wire N__34337;
    wire N__34334;
    wire N__34333;
    wire N__34330;
    wire N__34327;
    wire N__34326;
    wire N__34323;
    wire N__34318;
    wire N__34315;
    wire N__34308;
    wire N__34305;
    wire N__34302;
    wire N__34301;
    wire N__34298;
    wire N__34297;
    wire N__34296;
    wire N__34293;
    wire N__34290;
    wire N__34285;
    wire N__34278;
    wire N__34275;
    wire N__34274;
    wire N__34273;
    wire N__34270;
    wire N__34267;
    wire N__34262;
    wire N__34257;
    wire N__34254;
    wire N__34253;
    wire N__34252;
    wire N__34249;
    wire N__34244;
    wire N__34239;
    wire N__34236;
    wire N__34233;
    wire N__34230;
    wire N__34227;
    wire N__34224;
    wire N__34221;
    wire N__34218;
    wire N__34215;
    wire N__34212;
    wire N__34209;
    wire N__34206;
    wire N__34203;
    wire N__34200;
    wire N__34197;
    wire N__34194;
    wire N__34193;
    wire N__34190;
    wire N__34187;
    wire N__34184;
    wire N__34181;
    wire N__34178;
    wire N__34175;
    wire N__34172;
    wire N__34169;
    wire N__34166;
    wire N__34163;
    wire N__34160;
    wire N__34157;
    wire N__34154;
    wire N__34153;
    wire N__34150;
    wire N__34147;
    wire N__34144;
    wire N__34141;
    wire N__34138;
    wire N__34131;
    wire N__34128;
    wire N__34125;
    wire N__34122;
    wire N__34119;
    wire N__34116;
    wire N__34113;
    wire N__34110;
    wire N__34107;
    wire N__34104;
    wire N__34101;
    wire N__34098;
    wire N__34095;
    wire N__34092;
    wire N__34091;
    wire N__34088;
    wire N__34085;
    wire N__34082;
    wire N__34079;
    wire N__34076;
    wire N__34073;
    wire N__34070;
    wire N__34067;
    wire N__34064;
    wire N__34061;
    wire N__34058;
    wire N__34055;
    wire N__34052;
    wire N__34049;
    wire N__34046;
    wire N__34045;
    wire N__34042;
    wire N__34039;
    wire N__34036;
    wire N__34033;
    wire N__34030;
    wire N__34023;
    wire N__34020;
    wire N__34017;
    wire N__34014;
    wire N__34011;
    wire N__34008;
    wire N__34005;
    wire N__34002;
    wire N__33999;
    wire N__33996;
    wire N__33993;
    wire N__33990;
    wire N__33987;
    wire N__33984;
    wire N__33981;
    wire N__33978;
    wire N__33977;
    wire N__33974;
    wire N__33971;
    wire N__33968;
    wire N__33965;
    wire N__33962;
    wire N__33959;
    wire N__33956;
    wire N__33953;
    wire N__33950;
    wire N__33947;
    wire N__33944;
    wire N__33941;
    wire N__33938;
    wire N__33937;
    wire N__33934;
    wire N__33931;
    wire N__33928;
    wire N__33925;
    wire N__33922;
    wire N__33915;
    wire N__33912;
    wire N__33909;
    wire N__33906;
    wire N__33903;
    wire N__33900;
    wire N__33897;
    wire N__33894;
    wire N__33891;
    wire N__33888;
    wire N__33885;
    wire N__33882;
    wire N__33879;
    wire N__33876;
    wire N__33873;
    wire N__33870;
    wire N__33867;
    wire N__33864;
    wire N__33863;
    wire N__33860;
    wire N__33857;
    wire N__33854;
    wire N__33851;
    wire N__33848;
    wire N__33845;
    wire N__33842;
    wire N__33839;
    wire N__33836;
    wire N__33835;
    wire N__33832;
    wire N__33829;
    wire N__33826;
    wire N__33821;
    wire N__33816;
    wire N__33813;
    wire N__33810;
    wire N__33807;
    wire N__33804;
    wire N__33803;
    wire N__33800;
    wire N__33797;
    wire N__33796;
    wire N__33791;
    wire N__33788;
    wire N__33783;
    wire N__33780;
    wire N__33777;
    wire N__33776;
    wire N__33773;
    wire N__33772;
    wire N__33769;
    wire N__33766;
    wire N__33761;
    wire N__33756;
    wire N__33753;
    wire N__33750;
    wire N__33747;
    wire N__33744;
    wire N__33741;
    wire N__33738;
    wire N__33735;
    wire N__33732;
    wire N__33729;
    wire N__33726;
    wire N__33723;
    wire N__33720;
    wire N__33717;
    wire N__33714;
    wire N__33713;
    wire N__33710;
    wire N__33707;
    wire N__33704;
    wire N__33701;
    wire N__33698;
    wire N__33695;
    wire N__33692;
    wire N__33689;
    wire N__33686;
    wire N__33683;
    wire N__33680;
    wire N__33677;
    wire N__33674;
    wire N__33673;
    wire N__33670;
    wire N__33667;
    wire N__33664;
    wire N__33659;
    wire N__33654;
    wire N__33651;
    wire N__33648;
    wire N__33645;
    wire N__33642;
    wire N__33639;
    wire N__33636;
    wire N__33633;
    wire N__33630;
    wire N__33627;
    wire N__33624;
    wire N__33621;
    wire N__33618;
    wire N__33615;
    wire N__33612;
    wire N__33611;
    wire N__33608;
    wire N__33605;
    wire N__33602;
    wire N__33599;
    wire N__33596;
    wire N__33593;
    wire N__33590;
    wire N__33587;
    wire N__33584;
    wire N__33581;
    wire N__33578;
    wire N__33575;
    wire N__33572;
    wire N__33571;
    wire N__33568;
    wire N__33565;
    wire N__33562;
    wire N__33559;
    wire N__33556;
    wire N__33549;
    wire N__33546;
    wire N__33543;
    wire N__33540;
    wire N__33537;
    wire N__33534;
    wire N__33531;
    wire N__33528;
    wire N__33525;
    wire N__33522;
    wire N__33519;
    wire N__33516;
    wire N__33513;
    wire N__33510;
    wire N__33507;
    wire N__33504;
    wire N__33501;
    wire N__33500;
    wire N__33497;
    wire N__33494;
    wire N__33491;
    wire N__33488;
    wire N__33485;
    wire N__33482;
    wire N__33479;
    wire N__33476;
    wire N__33473;
    wire N__33470;
    wire N__33467;
    wire N__33464;
    wire N__33461;
    wire N__33460;
    wire N__33457;
    wire N__33454;
    wire N__33451;
    wire N__33448;
    wire N__33445;
    wire N__33438;
    wire N__33435;
    wire N__33432;
    wire N__33429;
    wire N__33426;
    wire N__33423;
    wire N__33420;
    wire N__33417;
    wire N__33414;
    wire N__33411;
    wire N__33408;
    wire N__33405;
    wire N__33402;
    wire N__33399;
    wire N__33396;
    wire N__33393;
    wire N__33390;
    wire N__33389;
    wire N__33386;
    wire N__33383;
    wire N__33380;
    wire N__33377;
    wire N__33374;
    wire N__33371;
    wire N__33368;
    wire N__33365;
    wire N__33362;
    wire N__33359;
    wire N__33356;
    wire N__33353;
    wire N__33350;
    wire N__33349;
    wire N__33346;
    wire N__33343;
    wire N__33340;
    wire N__33337;
    wire N__33334;
    wire N__33327;
    wire N__33324;
    wire N__33321;
    wire N__33318;
    wire N__33315;
    wire N__33312;
    wire N__33309;
    wire N__33306;
    wire N__33303;
    wire N__33300;
    wire N__33297;
    wire N__33294;
    wire N__33291;
    wire N__33288;
    wire N__33285;
    wire N__33282;
    wire N__33279;
    wire N__33276;
    wire N__33275;
    wire N__33272;
    wire N__33269;
    wire N__33266;
    wire N__33263;
    wire N__33260;
    wire N__33257;
    wire N__33254;
    wire N__33251;
    wire N__33248;
    wire N__33247;
    wire N__33244;
    wire N__33241;
    wire N__33238;
    wire N__33235;
    wire N__33232;
    wire N__33225;
    wire N__33222;
    wire N__33219;
    wire N__33216;
    wire N__33213;
    wire N__33210;
    wire N__33207;
    wire N__33204;
    wire N__33201;
    wire N__33198;
    wire N__33195;
    wire N__33192;
    wire N__33189;
    wire N__33186;
    wire N__33183;
    wire N__33182;
    wire N__33179;
    wire N__33176;
    wire N__33173;
    wire N__33170;
    wire N__33167;
    wire N__33164;
    wire N__33161;
    wire N__33158;
    wire N__33155;
    wire N__33152;
    wire N__33149;
    wire N__33146;
    wire N__33143;
    wire N__33142;
    wire N__33139;
    wire N__33136;
    wire N__33133;
    wire N__33130;
    wire N__33127;
    wire N__33120;
    wire N__33117;
    wire N__33114;
    wire N__33113;
    wire N__33110;
    wire N__33107;
    wire N__33104;
    wire N__33101;
    wire N__33098;
    wire N__33097;
    wire N__33092;
    wire N__33089;
    wire N__33084;
    wire N__33083;
    wire N__33080;
    wire N__33079;
    wire N__33076;
    wire N__33073;
    wire N__33070;
    wire N__33067;
    wire N__33064;
    wire N__33061;
    wire N__33056;
    wire N__33053;
    wire N__33048;
    wire N__33045;
    wire N__33042;
    wire N__33041;
    wire N__33040;
    wire N__33037;
    wire N__33032;
    wire N__33027;
    wire N__33024;
    wire N__33023;
    wire N__33020;
    wire N__33017;
    wire N__33016;
    wire N__33013;
    wire N__33010;
    wire N__33007;
    wire N__33004;
    wire N__32997;
    wire N__32996;
    wire N__32995;
    wire N__32992;
    wire N__32989;
    wire N__32986;
    wire N__32983;
    wire N__32976;
    wire N__32975;
    wire N__32972;
    wire N__32971;
    wire N__32968;
    wire N__32965;
    wire N__32962;
    wire N__32955;
    wire N__32952;
    wire N__32949;
    wire N__32946;
    wire N__32943;
    wire N__32940;
    wire N__32937;
    wire N__32934;
    wire N__32931;
    wire N__32928;
    wire N__32925;
    wire N__32922;
    wire N__32919;
    wire N__32916;
    wire N__32913;
    wire N__32910;
    wire N__32907;
    wire N__32904;
    wire N__32901;
    wire N__32900;
    wire N__32897;
    wire N__32894;
    wire N__32891;
    wire N__32888;
    wire N__32885;
    wire N__32882;
    wire N__32879;
    wire N__32876;
    wire N__32873;
    wire N__32870;
    wire N__32867;
    wire N__32864;
    wire N__32861;
    wire N__32858;
    wire N__32855;
    wire N__32852;
    wire N__32849;
    wire N__32844;
    wire N__32841;
    wire N__32838;
    wire N__32835;
    wire N__32832;
    wire N__32829;
    wire N__32826;
    wire N__32823;
    wire N__32820;
    wire N__32817;
    wire N__32816;
    wire N__32815;
    wire N__32810;
    wire N__32807;
    wire N__32804;
    wire N__32801;
    wire N__32796;
    wire N__32793;
    wire N__32790;
    wire N__32787;
    wire N__32786;
    wire N__32783;
    wire N__32780;
    wire N__32779;
    wire N__32776;
    wire N__32773;
    wire N__32770;
    wire N__32763;
    wire N__32760;
    wire N__32757;
    wire N__32756;
    wire N__32753;
    wire N__32750;
    wire N__32749;
    wire N__32746;
    wire N__32743;
    wire N__32740;
    wire N__32737;
    wire N__32734;
    wire N__32727;
    wire N__32726;
    wire N__32723;
    wire N__32720;
    wire N__32719;
    wire N__32716;
    wire N__32713;
    wire N__32710;
    wire N__32707;
    wire N__32704;
    wire N__32697;
    wire N__32694;
    wire N__32691;
    wire N__32688;
    wire N__32687;
    wire N__32684;
    wire N__32683;
    wire N__32680;
    wire N__32677;
    wire N__32674;
    wire N__32667;
    wire N__32664;
    wire N__32661;
    wire N__32660;
    wire N__32659;
    wire N__32656;
    wire N__32651;
    wire N__32646;
    wire N__32643;
    wire N__32640;
    wire N__32637;
    wire N__32634;
    wire N__32631;
    wire N__32628;
    wire N__32625;
    wire N__32622;
    wire N__32619;
    wire N__32616;
    wire N__32613;
    wire N__32610;
    wire N__32607;
    wire N__32604;
    wire N__32601;
    wire N__32600;
    wire N__32597;
    wire N__32594;
    wire N__32591;
    wire N__32588;
    wire N__32585;
    wire N__32580;
    wire N__32577;
    wire N__32574;
    wire N__32571;
    wire N__32568;
    wire N__32565;
    wire N__32562;
    wire N__32561;
    wire N__32558;
    wire N__32555;
    wire N__32554;
    wire N__32551;
    wire N__32548;
    wire N__32545;
    wire N__32538;
    wire N__32535;
    wire N__32532;
    wire N__32529;
    wire N__32526;
    wire N__32525;
    wire N__32522;
    wire N__32519;
    wire N__32518;
    wire N__32513;
    wire N__32510;
    wire N__32507;
    wire N__32502;
    wire N__32499;
    wire N__32496;
    wire N__32493;
    wire N__32490;
    wire N__32489;
    wire N__32486;
    wire N__32483;
    wire N__32480;
    wire N__32477;
    wire N__32472;
    wire N__32469;
    wire N__32468;
    wire N__32465;
    wire N__32462;
    wire N__32461;
    wire N__32458;
    wire N__32455;
    wire N__32452;
    wire N__32449;
    wire N__32446;
    wire N__32439;
    wire N__32436;
    wire N__32433;
    wire N__32430;
    wire N__32427;
    wire N__32424;
    wire N__32421;
    wire N__32420;
    wire N__32415;
    wire N__32412;
    wire N__32411;
    wire N__32408;
    wire N__32405;
    wire N__32402;
    wire N__32399;
    wire N__32396;
    wire N__32391;
    wire N__32390;
    wire N__32387;
    wire N__32384;
    wire N__32381;
    wire N__32378;
    wire N__32377;
    wire N__32372;
    wire N__32369;
    wire N__32364;
    wire N__32361;
    wire N__32358;
    wire N__32355;
    wire N__32352;
    wire N__32349;
    wire N__32346;
    wire N__32343;
    wire N__32340;
    wire N__32337;
    wire N__32334;
    wire N__32331;
    wire N__32328;
    wire N__32327;
    wire N__32324;
    wire N__32321;
    wire N__32318;
    wire N__32313;
    wire N__32310;
    wire N__32307;
    wire N__32306;
    wire N__32305;
    wire N__32302;
    wire N__32299;
    wire N__32296;
    wire N__32293;
    wire N__32290;
    wire N__32283;
    wire N__32280;
    wire N__32277;
    wire N__32274;
    wire N__32271;
    wire N__32270;
    wire N__32267;
    wire N__32264;
    wire N__32261;
    wire N__32256;
    wire N__32255;
    wire N__32252;
    wire N__32249;
    wire N__32246;
    wire N__32245;
    wire N__32242;
    wire N__32239;
    wire N__32236;
    wire N__32233;
    wire N__32226;
    wire N__32223;
    wire N__32220;
    wire N__32217;
    wire N__32216;
    wire N__32215;
    wire N__32212;
    wire N__32207;
    wire N__32202;
    wire N__32199;
    wire N__32196;
    wire N__32195;
    wire N__32192;
    wire N__32189;
    wire N__32184;
    wire N__32181;
    wire N__32178;
    wire N__32175;
    wire N__32174;
    wire N__32171;
    wire N__32168;
    wire N__32163;
    wire N__32162;
    wire N__32159;
    wire N__32156;
    wire N__32153;
    wire N__32148;
    wire N__32145;
    wire N__32142;
    wire N__32141;
    wire N__32138;
    wire N__32135;
    wire N__32132;
    wire N__32129;
    wire N__32128;
    wire N__32125;
    wire N__32122;
    wire N__32119;
    wire N__32116;
    wire N__32113;
    wire N__32106;
    wire N__32103;
    wire N__32100;
    wire N__32097;
    wire N__32094;
    wire N__32091;
    wire N__32090;
    wire N__32089;
    wire N__32086;
    wire N__32083;
    wire N__32080;
    wire N__32073;
    wire N__32070;
    wire N__32069;
    wire N__32066;
    wire N__32063;
    wire N__32060;
    wire N__32057;
    wire N__32054;
    wire N__32049;
    wire N__32046;
    wire N__32043;
    wire N__32042;
    wire N__32039;
    wire N__32036;
    wire N__32033;
    wire N__32030;
    wire N__32025;
    wire N__32022;
    wire N__32019;
    wire N__32016;
    wire N__32013;
    wire N__32010;
    wire N__32007;
    wire N__32004;
    wire N__32001;
    wire N__31998;
    wire N__31995;
    wire N__31992;
    wire N__31991;
    wire N__31990;
    wire N__31987;
    wire N__31982;
    wire N__31979;
    wire N__31974;
    wire N__31971;
    wire N__31968;
    wire N__31967;
    wire N__31966;
    wire N__31963;
    wire N__31958;
    wire N__31953;
    wire N__31950;
    wire N__31947;
    wire N__31944;
    wire N__31941;
    wire N__31938;
    wire N__31935;
    wire N__31932;
    wire N__31929;
    wire N__31928;
    wire N__31925;
    wire N__31922;
    wire N__31919;
    wire N__31914;
    wire N__31911;
    wire N__31908;
    wire N__31905;
    wire N__31902;
    wire N__31899;
    wire N__31896;
    wire N__31895;
    wire N__31892;
    wire N__31889;
    wire N__31884;
    wire N__31881;
    wire N__31878;
    wire N__31875;
    wire N__31872;
    wire N__31871;
    wire N__31868;
    wire N__31865;
    wire N__31860;
    wire N__31859;
    wire N__31856;
    wire N__31853;
    wire N__31850;
    wire N__31845;
    wire N__31844;
    wire N__31841;
    wire N__31838;
    wire N__31833;
    wire N__31832;
    wire N__31829;
    wire N__31826;
    wire N__31821;
    wire N__31818;
    wire N__31817;
    wire N__31814;
    wire N__31811;
    wire N__31808;
    wire N__31803;
    wire N__31802;
    wire N__31799;
    wire N__31796;
    wire N__31791;
    wire N__31788;
    wire N__31785;
    wire N__31784;
    wire N__31781;
    wire N__31778;
    wire N__31773;
    wire N__31772;
    wire N__31769;
    wire N__31766;
    wire N__31761;
    wire N__31760;
    wire N__31757;
    wire N__31754;
    wire N__31751;
    wire N__31746;
    wire N__31745;
    wire N__31742;
    wire N__31739;
    wire N__31734;
    wire N__31731;
    wire N__31728;
    wire N__31727;
    wire N__31724;
    wire N__31721;
    wire N__31718;
    wire N__31715;
    wire N__31710;
    wire N__31707;
    wire N__31704;
    wire N__31701;
    wire N__31698;
    wire N__31695;
    wire N__31692;
    wire N__31689;
    wire N__31686;
    wire N__31683;
    wire N__31680;
    wire N__31677;
    wire N__31674;
    wire N__31671;
    wire N__31668;
    wire N__31665;
    wire N__31662;
    wire N__31661;
    wire N__31658;
    wire N__31655;
    wire N__31652;
    wire N__31649;
    wire N__31646;
    wire N__31643;
    wire N__31640;
    wire N__31635;
    wire N__31632;
    wire N__31629;
    wire N__31626;
    wire N__31625;
    wire N__31624;
    wire N__31621;
    wire N__31620;
    wire N__31619;
    wire N__31618;
    wire N__31617;
    wire N__31614;
    wire N__31611;
    wire N__31610;
    wire N__31609;
    wire N__31608;
    wire N__31605;
    wire N__31602;
    wire N__31601;
    wire N__31600;
    wire N__31597;
    wire N__31594;
    wire N__31591;
    wire N__31590;
    wire N__31589;
    wire N__31588;
    wire N__31587;
    wire N__31586;
    wire N__31585;
    wire N__31584;
    wire N__31583;
    wire N__31582;
    wire N__31581;
    wire N__31580;
    wire N__31577;
    wire N__31570;
    wire N__31567;
    wire N__31562;
    wire N__31549;
    wire N__31540;
    wire N__31537;
    wire N__31526;
    wire N__31521;
    wire N__31518;
    wire N__31513;
    wire N__31502;
    wire N__31497;
    wire N__31494;
    wire N__31493;
    wire N__31490;
    wire N__31487;
    wire N__31484;
    wire N__31481;
    wire N__31478;
    wire N__31475;
    wire N__31470;
    wire N__31467;
    wire N__31464;
    wire N__31461;
    wire N__31458;
    wire N__31455;
    wire N__31452;
    wire N__31449;
    wire N__31448;
    wire N__31447;
    wire N__31444;
    wire N__31439;
    wire N__31434;
    wire N__31431;
    wire N__31428;
    wire N__31425;
    wire N__31422;
    wire N__31419;
    wire N__31416;
    wire N__31413;
    wire N__31410;
    wire N__31407;
    wire N__31404;
    wire N__31401;
    wire N__31398;
    wire N__31395;
    wire N__31392;
    wire N__31389;
    wire N__31386;
    wire N__31383;
    wire N__31380;
    wire N__31377;
    wire N__31374;
    wire N__31371;
    wire N__31368;
    wire N__31367;
    wire N__31366;
    wire N__31363;
    wire N__31360;
    wire N__31357;
    wire N__31350;
    wire N__31347;
    wire N__31344;
    wire N__31341;
    wire N__31338;
    wire N__31335;
    wire N__31332;
    wire N__31329;
    wire N__31326;
    wire N__31323;
    wire N__31320;
    wire N__31319;
    wire N__31318;
    wire N__31315;
    wire N__31312;
    wire N__31309;
    wire N__31306;
    wire N__31299;
    wire N__31298;
    wire N__31295;
    wire N__31294;
    wire N__31291;
    wire N__31288;
    wire N__31285;
    wire N__31282;
    wire N__31279;
    wire N__31276;
    wire N__31273;
    wire N__31270;
    wire N__31263;
    wire N__31260;
    wire N__31257;
    wire N__31254;
    wire N__31253;
    wire N__31252;
    wire N__31249;
    wire N__31246;
    wire N__31243;
    wire N__31238;
    wire N__31233;
    wire N__31230;
    wire N__31227;
    wire N__31224;
    wire N__31221;
    wire N__31218;
    wire N__31215;
    wire N__31212;
    wire N__31209;
    wire N__31206;
    wire N__31203;
    wire N__31200;
    wire N__31199;
    wire N__31198;
    wire N__31195;
    wire N__31190;
    wire N__31185;
    wire N__31184;
    wire N__31181;
    wire N__31178;
    wire N__31175;
    wire N__31172;
    wire N__31171;
    wire N__31166;
    wire N__31163;
    wire N__31158;
    wire N__31155;
    wire N__31154;
    wire N__31151;
    wire N__31148;
    wire N__31145;
    wire N__31140;
    wire N__31137;
    wire N__31134;
    wire N__31131;
    wire N__31128;
    wire N__31125;
    wire N__31122;
    wire N__31121;
    wire N__31118;
    wire N__31115;
    wire N__31112;
    wire N__31109;
    wire N__31106;
    wire N__31103;
    wire N__31098;
    wire N__31095;
    wire N__31092;
    wire N__31091;
    wire N__31088;
    wire N__31085;
    wire N__31082;
    wire N__31081;
    wire N__31078;
    wire N__31075;
    wire N__31072;
    wire N__31069;
    wire N__31062;
    wire N__31059;
    wire N__31056;
    wire N__31053;
    wire N__31050;
    wire N__31047;
    wire N__31046;
    wire N__31045;
    wire N__31040;
    wire N__31037;
    wire N__31034;
    wire N__31031;
    wire N__31030;
    wire N__31029;
    wire N__31028;
    wire N__31025;
    wire N__31022;
    wire N__31017;
    wire N__31014;
    wire N__31011;
    wire N__31006;
    wire N__30999;
    wire N__30996;
    wire N__30995;
    wire N__30992;
    wire N__30989;
    wire N__30984;
    wire N__30983;
    wire N__30982;
    wire N__30981;
    wire N__30980;
    wire N__30979;
    wire N__30976;
    wire N__30973;
    wire N__30970;
    wire N__30969;
    wire N__30968;
    wire N__30967;
    wire N__30966;
    wire N__30965;
    wire N__30964;
    wire N__30963;
    wire N__30962;
    wire N__30959;
    wire N__30956;
    wire N__30955;
    wire N__30944;
    wire N__30937;
    wire N__30932;
    wire N__30929;
    wire N__30920;
    wire N__30909;
    wire N__30908;
    wire N__30905;
    wire N__30902;
    wire N__30897;
    wire N__30894;
    wire N__30893;
    wire N__30890;
    wire N__30889;
    wire N__30886;
    wire N__30883;
    wire N__30880;
    wire N__30873;
    wire N__30872;
    wire N__30869;
    wire N__30866;
    wire N__30863;
    wire N__30862;
    wire N__30857;
    wire N__30854;
    wire N__30849;
    wire N__30846;
    wire N__30845;
    wire N__30842;
    wire N__30841;
    wire N__30838;
    wire N__30835;
    wire N__30832;
    wire N__30827;
    wire N__30822;
    wire N__30819;
    wire N__30816;
    wire N__30813;
    wire N__30810;
    wire N__30807;
    wire N__30806;
    wire N__30805;
    wire N__30802;
    wire N__30799;
    wire N__30796;
    wire N__30793;
    wire N__30790;
    wire N__30787;
    wire N__30780;
    wire N__30779;
    wire N__30778;
    wire N__30775;
    wire N__30772;
    wire N__30769;
    wire N__30766;
    wire N__30763;
    wire N__30760;
    wire N__30757;
    wire N__30754;
    wire N__30749;
    wire N__30746;
    wire N__30741;
    wire N__30738;
    wire N__30735;
    wire N__30732;
    wire N__30729;
    wire N__30726;
    wire N__30723;
    wire N__30722;
    wire N__30721;
    wire N__30718;
    wire N__30715;
    wire N__30712;
    wire N__30709;
    wire N__30706;
    wire N__30703;
    wire N__30700;
    wire N__30697;
    wire N__30694;
    wire N__30689;
    wire N__30686;
    wire N__30681;
    wire N__30678;
    wire N__30677;
    wire N__30674;
    wire N__30671;
    wire N__30668;
    wire N__30665;
    wire N__30662;
    wire N__30657;
    wire N__30654;
    wire N__30651;
    wire N__30648;
    wire N__30645;
    wire N__30642;
    wire N__30639;
    wire N__30636;
    wire N__30633;
    wire N__30630;
    wire N__30627;
    wire N__30624;
    wire N__30621;
    wire N__30620;
    wire N__30617;
    wire N__30614;
    wire N__30609;
    wire N__30608;
    wire N__30605;
    wire N__30602;
    wire N__30601;
    wire N__30598;
    wire N__30595;
    wire N__30592;
    wire N__30589;
    wire N__30586;
    wire N__30579;
    wire N__30576;
    wire N__30573;
    wire N__30570;
    wire N__30567;
    wire N__30564;
    wire N__30561;
    wire N__30558;
    wire N__30555;
    wire N__30552;
    wire N__30549;
    wire N__30546;
    wire N__30543;
    wire N__30542;
    wire N__30539;
    wire N__30536;
    wire N__30533;
    wire N__30530;
    wire N__30527;
    wire N__30526;
    wire N__30523;
    wire N__30520;
    wire N__30517;
    wire N__30514;
    wire N__30507;
    wire N__30504;
    wire N__30501;
    wire N__30498;
    wire N__30495;
    wire N__30492;
    wire N__30489;
    wire N__30486;
    wire N__30483;
    wire N__30480;
    wire N__30477;
    wire N__30474;
    wire N__30471;
    wire N__30468;
    wire N__30465;
    wire N__30462;
    wire N__30459;
    wire N__30456;
    wire N__30453;
    wire N__30450;
    wire N__30447;
    wire N__30444;
    wire N__30441;
    wire N__30438;
    wire N__30435;
    wire N__30432;
    wire N__30429;
    wire N__30426;
    wire N__30423;
    wire N__30422;
    wire N__30419;
    wire N__30416;
    wire N__30413;
    wire N__30408;
    wire N__30407;
    wire N__30404;
    wire N__30401;
    wire N__30396;
    wire N__30393;
    wire N__30392;
    wire N__30389;
    wire N__30386;
    wire N__30383;
    wire N__30378;
    wire N__30377;
    wire N__30374;
    wire N__30371;
    wire N__30366;
    wire N__30363;
    wire N__30360;
    wire N__30359;
    wire N__30356;
    wire N__30353;
    wire N__30348;
    wire N__30345;
    wire N__30342;
    wire N__30339;
    wire N__30336;
    wire N__30333;
    wire N__30330;
    wire N__30327;
    wire N__30324;
    wire N__30321;
    wire N__30318;
    wire N__30315;
    wire N__30312;
    wire N__30309;
    wire N__30306;
    wire N__30303;
    wire N__30300;
    wire N__30297;
    wire N__30294;
    wire N__30291;
    wire N__30288;
    wire N__30285;
    wire N__30282;
    wire N__30279;
    wire N__30278;
    wire N__30275;
    wire N__30274;
    wire N__30271;
    wire N__30268;
    wire N__30265;
    wire N__30262;
    wire N__30259;
    wire N__30256;
    wire N__30251;
    wire N__30246;
    wire N__30243;
    wire N__30240;
    wire N__30237;
    wire N__30236;
    wire N__30233;
    wire N__30230;
    wire N__30227;
    wire N__30222;
    wire N__30219;
    wire N__30216;
    wire N__30213;
    wire N__30210;
    wire N__30209;
    wire N__30206;
    wire N__30203;
    wire N__30198;
    wire N__30197;
    wire N__30194;
    wire N__30191;
    wire N__30186;
    wire N__30185;
    wire N__30182;
    wire N__30179;
    wire N__30176;
    wire N__30171;
    wire N__30170;
    wire N__30167;
    wire N__30164;
    wire N__30159;
    wire N__30156;
    wire N__30153;
    wire N__30150;
    wire N__30147;
    wire N__30144;
    wire N__30143;
    wire N__30140;
    wire N__30137;
    wire N__30132;
    wire N__30129;
    wire N__30126;
    wire N__30123;
    wire N__30120;
    wire N__30117;
    wire N__30114;
    wire N__30111;
    wire N__30110;
    wire N__30109;
    wire N__30108;
    wire N__30107;
    wire N__30106;
    wire N__30105;
    wire N__30104;
    wire N__30103;
    wire N__30102;
    wire N__30101;
    wire N__30100;
    wire N__30099;
    wire N__30098;
    wire N__30097;
    wire N__30096;
    wire N__30095;
    wire N__30094;
    wire N__30093;
    wire N__30090;
    wire N__30075;
    wire N__30074;
    wire N__30073;
    wire N__30072;
    wire N__30069;
    wire N__30066;
    wire N__30049;
    wire N__30046;
    wire N__30045;
    wire N__30042;
    wire N__30039;
    wire N__30032;
    wire N__30031;
    wire N__30026;
    wire N__30023;
    wire N__30020;
    wire N__30017;
    wire N__30016;
    wire N__30011;
    wire N__30008;
    wire N__30007;
    wire N__30004;
    wire N__30001;
    wire N__29998;
    wire N__29995;
    wire N__29990;
    wire N__29987;
    wire N__29984;
    wire N__29981;
    wire N__29978;
    wire N__29973;
    wire N__29968;
    wire N__29963;
    wire N__29952;
    wire N__29951;
    wire N__29948;
    wire N__29947;
    wire N__29946;
    wire N__29943;
    wire N__29942;
    wire N__29941;
    wire N__29934;
    wire N__29931;
    wire N__29928;
    wire N__29925;
    wire N__29922;
    wire N__29919;
    wire N__29914;
    wire N__29911;
    wire N__29910;
    wire N__29909;
    wire N__29908;
    wire N__29907;
    wire N__29904;
    wire N__29899;
    wire N__29894;
    wire N__29889;
    wire N__29880;
    wire N__29879;
    wire N__29878;
    wire N__29877;
    wire N__29876;
    wire N__29875;
    wire N__29874;
    wire N__29873;
    wire N__29872;
    wire N__29855;
    wire N__29854;
    wire N__29853;
    wire N__29852;
    wire N__29851;
    wire N__29848;
    wire N__29847;
    wire N__29846;
    wire N__29845;
    wire N__29844;
    wire N__29841;
    wire N__29840;
    wire N__29823;
    wire N__29822;
    wire N__29821;
    wire N__29820;
    wire N__29819;
    wire N__29816;
    wire N__29813;
    wire N__29810;
    wire N__29807;
    wire N__29804;
    wire N__29801;
    wire N__29798;
    wire N__29795;
    wire N__29794;
    wire N__29793;
    wire N__29792;
    wire N__29791;
    wire N__29790;
    wire N__29787;
    wire N__29782;
    wire N__29777;
    wire N__29774;
    wire N__29771;
    wire N__29768;
    wire N__29767;
    wire N__29760;
    wire N__29755;
    wire N__29750;
    wire N__29747;
    wire N__29742;
    wire N__29739;
    wire N__29736;
    wire N__29731;
    wire N__29718;
    wire N__29715;
    wire N__29712;
    wire N__29711;
    wire N__29708;
    wire N__29705;
    wire N__29702;
    wire N__29699;
    wire N__29694;
    wire N__29691;
    wire N__29688;
    wire N__29687;
    wire N__29686;
    wire N__29683;
    wire N__29680;
    wire N__29677;
    wire N__29670;
    wire N__29667;
    wire N__29666;
    wire N__29663;
    wire N__29660;
    wire N__29657;
    wire N__29654;
    wire N__29649;
    wire N__29646;
    wire N__29643;
    wire N__29642;
    wire N__29639;
    wire N__29636;
    wire N__29631;
    wire N__29628;
    wire N__29625;
    wire N__29622;
    wire N__29621;
    wire N__29618;
    wire N__29615;
    wire N__29610;
    wire N__29607;
    wire N__29604;
    wire N__29601;
    wire N__29600;
    wire N__29597;
    wire N__29594;
    wire N__29589;
    wire N__29586;
    wire N__29583;
    wire N__29582;
    wire N__29579;
    wire N__29576;
    wire N__29571;
    wire N__29568;
    wire N__29565;
    wire N__29564;
    wire N__29561;
    wire N__29558;
    wire N__29553;
    wire N__29550;
    wire N__29547;
    wire N__29544;
    wire N__29541;
    wire N__29540;
    wire N__29537;
    wire N__29534;
    wire N__29529;
    wire N__29526;
    wire N__29523;
    wire N__29520;
    wire N__29519;
    wire N__29516;
    wire N__29513;
    wire N__29508;
    wire N__29505;
    wire N__29502;
    wire N__29501;
    wire N__29498;
    wire N__29495;
    wire N__29492;
    wire N__29489;
    wire N__29484;
    wire N__29481;
    wire N__29478;
    wire N__29475;
    wire N__29474;
    wire N__29471;
    wire N__29468;
    wire N__29463;
    wire N__29460;
    wire N__29457;
    wire N__29456;
    wire N__29453;
    wire N__29452;
    wire N__29449;
    wire N__29446;
    wire N__29443;
    wire N__29440;
    wire N__29437;
    wire N__29430;
    wire N__29429;
    wire N__29428;
    wire N__29425;
    wire N__29422;
    wire N__29419;
    wire N__29416;
    wire N__29413;
    wire N__29410;
    wire N__29407;
    wire N__29402;
    wire N__29399;
    wire N__29394;
    wire N__29393;
    wire N__29392;
    wire N__29391;
    wire N__29390;
    wire N__29387;
    wire N__29386;
    wire N__29385;
    wire N__29384;
    wire N__29383;
    wire N__29382;
    wire N__29381;
    wire N__29380;
    wire N__29375;
    wire N__29374;
    wire N__29373;
    wire N__29372;
    wire N__29369;
    wire N__29366;
    wire N__29365;
    wire N__29364;
    wire N__29363;
    wire N__29362;
    wire N__29357;
    wire N__29354;
    wire N__29349;
    wire N__29344;
    wire N__29341;
    wire N__29338;
    wire N__29337;
    wire N__29336;
    wire N__29335;
    wire N__29334;
    wire N__29333;
    wire N__29332;
    wire N__29329;
    wire N__29328;
    wire N__29327;
    wire N__29326;
    wire N__29325;
    wire N__29324;
    wire N__29323;
    wire N__29320;
    wire N__29313;
    wire N__29308;
    wire N__29303;
    wire N__29298;
    wire N__29295;
    wire N__29292;
    wire N__29287;
    wire N__29284;
    wire N__29277;
    wire N__29272;
    wire N__29263;
    wire N__29256;
    wire N__29249;
    wire N__29246;
    wire N__29241;
    wire N__29236;
    wire N__29217;
    wire N__29214;
    wire N__29213;
    wire N__29210;
    wire N__29207;
    wire N__29202;
    wire N__29201;
    wire N__29198;
    wire N__29195;
    wire N__29192;
    wire N__29189;
    wire N__29188;
    wire N__29185;
    wire N__29182;
    wire N__29179;
    wire N__29176;
    wire N__29173;
    wire N__29166;
    wire N__29163;
    wire N__29160;
    wire N__29157;
    wire N__29154;
    wire N__29151;
    wire N__29148;
    wire N__29145;
    wire N__29142;
    wire N__29141;
    wire N__29140;
    wire N__29139;
    wire N__29138;
    wire N__29137;
    wire N__29136;
    wire N__29135;
    wire N__29134;
    wire N__29131;
    wire N__29128;
    wire N__29125;
    wire N__29122;
    wire N__29119;
    wire N__29118;
    wire N__29117;
    wire N__29116;
    wire N__29115;
    wire N__29114;
    wire N__29097;
    wire N__29094;
    wire N__29093;
    wire N__29092;
    wire N__29091;
    wire N__29088;
    wire N__29085;
    wire N__29084;
    wire N__29083;
    wire N__29082;
    wire N__29081;
    wire N__29080;
    wire N__29077;
    wire N__29074;
    wire N__29071;
    wire N__29070;
    wire N__29067;
    wire N__29064;
    wire N__29047;
    wire N__29034;
    wire N__29031;
    wire N__29028;
    wire N__29023;
    wire N__29020;
    wire N__29017;
    wire N__29014;
    wire N__29007;
    wire N__29004;
    wire N__29001;
    wire N__28998;
    wire N__28995;
    wire N__28994;
    wire N__28991;
    wire N__28990;
    wire N__28987;
    wire N__28984;
    wire N__28981;
    wire N__28978;
    wire N__28971;
    wire N__28968;
    wire N__28965;
    wire N__28962;
    wire N__28961;
    wire N__28960;
    wire N__28957;
    wire N__28952;
    wire N__28947;
    wire N__28944;
    wire N__28941;
    wire N__28940;
    wire N__28937;
    wire N__28934;
    wire N__28933;
    wire N__28930;
    wire N__28927;
    wire N__28924;
    wire N__28921;
    wire N__28918;
    wire N__28911;
    wire N__28908;
    wire N__28907;
    wire N__28904;
    wire N__28901;
    wire N__28900;
    wire N__28897;
    wire N__28892;
    wire N__28887;
    wire N__28886;
    wire N__28883;
    wire N__28880;
    wire N__28879;
    wire N__28876;
    wire N__28873;
    wire N__28870;
    wire N__28863;
    wire N__28862;
    wire N__28859;
    wire N__28856;
    wire N__28851;
    wire N__28848;
    wire N__28847;
    wire N__28846;
    wire N__28843;
    wire N__28840;
    wire N__28839;
    wire N__28836;
    wire N__28833;
    wire N__28830;
    wire N__28827;
    wire N__28826;
    wire N__28823;
    wire N__28816;
    wire N__28813;
    wire N__28806;
    wire N__28803;
    wire N__28802;
    wire N__28801;
    wire N__28798;
    wire N__28795;
    wire N__28792;
    wire N__28787;
    wire N__28786;
    wire N__28785;
    wire N__28782;
    wire N__28779;
    wire N__28774;
    wire N__28771;
    wire N__28764;
    wire N__28761;
    wire N__28758;
    wire N__28755;
    wire N__28752;
    wire N__28749;
    wire N__28746;
    wire N__28745;
    wire N__28742;
    wire N__28739;
    wire N__28738;
    wire N__28735;
    wire N__28732;
    wire N__28729;
    wire N__28722;
    wire N__28719;
    wire N__28716;
    wire N__28713;
    wire N__28710;
    wire N__28709;
    wire N__28708;
    wire N__28705;
    wire N__28702;
    wire N__28699;
    wire N__28698;
    wire N__28697;
    wire N__28692;
    wire N__28689;
    wire N__28686;
    wire N__28683;
    wire N__28680;
    wire N__28677;
    wire N__28674;
    wire N__28665;
    wire N__28664;
    wire N__28661;
    wire N__28658;
    wire N__28655;
    wire N__28650;
    wire N__28647;
    wire N__28644;
    wire N__28643;
    wire N__28640;
    wire N__28637;
    wire N__28632;
    wire N__28631;
    wire N__28628;
    wire N__28627;
    wire N__28626;
    wire N__28623;
    wire N__28622;
    wire N__28621;
    wire N__28618;
    wire N__28615;
    wire N__28614;
    wire N__28611;
    wire N__28610;
    wire N__28607;
    wire N__28604;
    wire N__28603;
    wire N__28602;
    wire N__28599;
    wire N__28596;
    wire N__28593;
    wire N__28590;
    wire N__28587;
    wire N__28584;
    wire N__28579;
    wire N__28576;
    wire N__28575;
    wire N__28572;
    wire N__28571;
    wire N__28568;
    wire N__28563;
    wire N__28560;
    wire N__28555;
    wire N__28550;
    wire N__28547;
    wire N__28544;
    wire N__28541;
    wire N__28538;
    wire N__28533;
    wire N__28528;
    wire N__28525;
    wire N__28520;
    wire N__28511;
    wire N__28508;
    wire N__28505;
    wire N__28502;
    wire N__28499;
    wire N__28494;
    wire N__28491;
    wire N__28488;
    wire N__28485;
    wire N__28482;
    wire N__28481;
    wire N__28478;
    wire N__28475;
    wire N__28472;
    wire N__28467;
    wire N__28464;
    wire N__28461;
    wire N__28458;
    wire N__28455;
    wire N__28452;
    wire N__28449;
    wire N__28446;
    wire N__28443;
    wire N__28440;
    wire N__28437;
    wire N__28434;
    wire N__28433;
    wire N__28432;
    wire N__28429;
    wire N__28426;
    wire N__28423;
    wire N__28418;
    wire N__28415;
    wire N__28412;
    wire N__28407;
    wire N__28404;
    wire N__28403;
    wire N__28400;
    wire N__28397;
    wire N__28392;
    wire N__28389;
    wire N__28386;
    wire N__28383;
    wire N__28380;
    wire N__28377;
    wire N__28374;
    wire N__28371;
    wire N__28368;
    wire N__28365;
    wire N__28362;
    wire N__28359;
    wire N__28356;
    wire N__28353;
    wire N__28350;
    wire N__28347;
    wire N__28344;
    wire N__28341;
    wire N__28338;
    wire N__28337;
    wire N__28334;
    wire N__28331;
    wire N__28328;
    wire N__28325;
    wire N__28320;
    wire N__28317;
    wire N__28314;
    wire N__28313;
    wire N__28312;
    wire N__28309;
    wire N__28306;
    wire N__28303;
    wire N__28300;
    wire N__28297;
    wire N__28292;
    wire N__28287;
    wire N__28284;
    wire N__28283;
    wire N__28280;
    wire N__28277;
    wire N__28272;
    wire N__28269;
    wire N__28268;
    wire N__28267;
    wire N__28266;
    wire N__28265;
    wire N__28262;
    wire N__28257;
    wire N__28256;
    wire N__28255;
    wire N__28254;
    wire N__28251;
    wire N__28248;
    wire N__28247;
    wire N__28246;
    wire N__28245;
    wire N__28244;
    wire N__28241;
    wire N__28240;
    wire N__28239;
    wire N__28238;
    wire N__28237;
    wire N__28234;
    wire N__28227;
    wire N__28224;
    wire N__28221;
    wire N__28216;
    wire N__28215;
    wire N__28214;
    wire N__28213;
    wire N__28212;
    wire N__28211;
    wire N__28210;
    wire N__28205;
    wire N__28202;
    wire N__28195;
    wire N__28192;
    wire N__28191;
    wire N__28190;
    wire N__28189;
    wire N__28188;
    wire N__28187;
    wire N__28186;
    wire N__28185;
    wire N__28180;
    wire N__28173;
    wire N__28160;
    wire N__28157;
    wire N__28150;
    wire N__28145;
    wire N__28138;
    wire N__28133;
    wire N__28132;
    wire N__28131;
    wire N__28130;
    wire N__28127;
    wire N__28122;
    wire N__28117;
    wire N__28112;
    wire N__28109;
    wire N__28102;
    wire N__28089;
    wire N__28088;
    wire N__28085;
    wire N__28082;
    wire N__28079;
    wire N__28078;
    wire N__28075;
    wire N__28072;
    wire N__28069;
    wire N__28062;
    wire N__28059;
    wire N__28056;
    wire N__28053;
    wire N__28050;
    wire N__28047;
    wire N__28046;
    wire N__28043;
    wire N__28040;
    wire N__28035;
    wire N__28034;
    wire N__28031;
    wire N__28028;
    wire N__28023;
    wire N__28020;
    wire N__28019;
    wire N__28016;
    wire N__28013;
    wire N__28010;
    wire N__28007;
    wire N__28002;
    wire N__28001;
    wire N__28000;
    wire N__27999;
    wire N__27998;
    wire N__27997;
    wire N__27992;
    wire N__27991;
    wire N__27990;
    wire N__27989;
    wire N__27988;
    wire N__27985;
    wire N__27982;
    wire N__27981;
    wire N__27980;
    wire N__27979;
    wire N__27978;
    wire N__27977;
    wire N__27976;
    wire N__27975;
    wire N__27974;
    wire N__27973;
    wire N__27968;
    wire N__27967;
    wire N__27966;
    wire N__27965;
    wire N__27964;
    wire N__27961;
    wire N__27952;
    wire N__27947;
    wire N__27940;
    wire N__27937;
    wire N__27928;
    wire N__27925;
    wire N__27922;
    wire N__27917;
    wire N__27914;
    wire N__27911;
    wire N__27906;
    wire N__27899;
    wire N__27894;
    wire N__27887;
    wire N__27884;
    wire N__27883;
    wire N__27880;
    wire N__27877;
    wire N__27870;
    wire N__27867;
    wire N__27858;
    wire N__27857;
    wire N__27856;
    wire N__27855;
    wire N__27852;
    wire N__27851;
    wire N__27850;
    wire N__27849;
    wire N__27848;
    wire N__27847;
    wire N__27844;
    wire N__27843;
    wire N__27842;
    wire N__27841;
    wire N__27840;
    wire N__27839;
    wire N__27836;
    wire N__27835;
    wire N__27834;
    wire N__27833;
    wire N__27832;
    wire N__27831;
    wire N__27828;
    wire N__27827;
    wire N__27826;
    wire N__27825;
    wire N__27824;
    wire N__27823;
    wire N__27822;
    wire N__27821;
    wire N__27820;
    wire N__27817;
    wire N__27812;
    wire N__27807;
    wire N__27806;
    wire N__27805;
    wire N__27804;
    wire N__27803;
    wire N__27802;
    wire N__27801;
    wire N__27800;
    wire N__27797;
    wire N__27796;
    wire N__27795;
    wire N__27794;
    wire N__27793;
    wire N__27792;
    wire N__27791;
    wire N__27790;
    wire N__27787;
    wire N__27784;
    wire N__27779;
    wire N__27778;
    wire N__27773;
    wire N__27760;
    wire N__27759;
    wire N__27758;
    wire N__27757;
    wire N__27756;
    wire N__27755;
    wire N__27752;
    wire N__27747;
    wire N__27742;
    wire N__27733;
    wire N__27726;
    wire N__27725;
    wire N__27724;
    wire N__27723;
    wire N__27722;
    wire N__27721;
    wire N__27708;
    wire N__27705;
    wire N__27700;
    wire N__27687;
    wire N__27684;
    wire N__27679;
    wire N__27676;
    wire N__27671;
    wire N__27670;
    wire N__27669;
    wire N__27668;
    wire N__27665;
    wire N__27662;
    wire N__27659;
    wire N__27658;
    wire N__27657;
    wire N__27656;
    wire N__27655;
    wire N__27652;
    wire N__27651;
    wire N__27650;
    wire N__27647;
    wire N__27646;
    wire N__27645;
    wire N__27644;
    wire N__27639;
    wire N__27632;
    wire N__27631;
    wire N__27630;
    wire N__27629;
    wire N__27628;
    wire N__27621;
    wire N__27616;
    wire N__27613;
    wire N__27610;
    wire N__27601;
    wire N__27596;
    wire N__27589;
    wire N__27574;
    wire N__27571;
    wire N__27566;
    wire N__27557;
    wire N__27552;
    wire N__27543;
    wire N__27526;
    wire N__27513;
    wire N__27512;
    wire N__27509;
    wire N__27504;
    wire N__27501;
    wire N__27500;
    wire N__27497;
    wire N__27494;
    wire N__27489;
    wire N__27486;
    wire N__27483;
    wire N__27482;
    wire N__27481;
    wire N__27478;
    wire N__27473;
    wire N__27470;
    wire N__27465;
    wire N__27462;
    wire N__27459;
    wire N__27458;
    wire N__27455;
    wire N__27452;
    wire N__27449;
    wire N__27446;
    wire N__27445;
    wire N__27442;
    wire N__27439;
    wire N__27436;
    wire N__27429;
    wire N__27426;
    wire N__27425;
    wire N__27422;
    wire N__27421;
    wire N__27418;
    wire N__27415;
    wire N__27412;
    wire N__27409;
    wire N__27406;
    wire N__27403;
    wire N__27400;
    wire N__27397;
    wire N__27390;
    wire N__27387;
    wire N__27384;
    wire N__27383;
    wire N__27380;
    wire N__27377;
    wire N__27374;
    wire N__27373;
    wire N__27370;
    wire N__27367;
    wire N__27364;
    wire N__27361;
    wire N__27354;
    wire N__27351;
    wire N__27350;
    wire N__27347;
    wire N__27344;
    wire N__27341;
    wire N__27338;
    wire N__27333;
    wire N__27330;
    wire N__27329;
    wire N__27326;
    wire N__27325;
    wire N__27322;
    wire N__27319;
    wire N__27316;
    wire N__27313;
    wire N__27310;
    wire N__27307;
    wire N__27304;
    wire N__27301;
    wire N__27294;
    wire N__27293;
    wire N__27290;
    wire N__27287;
    wire N__27284;
    wire N__27281;
    wire N__27276;
    wire N__27273;
    wire N__27272;
    wire N__27269;
    wire N__27266;
    wire N__27263;
    wire N__27260;
    wire N__27259;
    wire N__27256;
    wire N__27253;
    wire N__27250;
    wire N__27247;
    wire N__27244;
    wire N__27237;
    wire N__27234;
    wire N__27231;
    wire N__27230;
    wire N__27227;
    wire N__27224;
    wire N__27223;
    wire N__27220;
    wire N__27217;
    wire N__27214;
    wire N__27211;
    wire N__27208;
    wire N__27201;
    wire N__27198;
    wire N__27195;
    wire N__27192;
    wire N__27189;
    wire N__27186;
    wire N__27183;
    wire N__27180;
    wire N__27179;
    wire N__27176;
    wire N__27173;
    wire N__27170;
    wire N__27167;
    wire N__27162;
    wire N__27159;
    wire N__27156;
    wire N__27153;
    wire N__27150;
    wire N__27149;
    wire N__27146;
    wire N__27143;
    wire N__27138;
    wire N__27137;
    wire N__27134;
    wire N__27131;
    wire N__27128;
    wire N__27123;
    wire N__27120;
    wire N__27117;
    wire N__27114;
    wire N__27113;
    wire N__27110;
    wire N__27107;
    wire N__27104;
    wire N__27101;
    wire N__27100;
    wire N__27097;
    wire N__27094;
    wire N__27091;
    wire N__27088;
    wire N__27085;
    wire N__27078;
    wire N__27077;
    wire N__27074;
    wire N__27071;
    wire N__27070;
    wire N__27067;
    wire N__27064;
    wire N__27061;
    wire N__27060;
    wire N__27057;
    wire N__27054;
    wire N__27053;
    wire N__27050;
    wire N__27047;
    wire N__27044;
    wire N__27041;
    wire N__27038;
    wire N__27033;
    wire N__27024;
    wire N__27021;
    wire N__27018;
    wire N__27017;
    wire N__27016;
    wire N__27015;
    wire N__27014;
    wire N__27011;
    wire N__27006;
    wire N__27001;
    wire N__26998;
    wire N__26995;
    wire N__26992;
    wire N__26985;
    wire N__26982;
    wire N__26979;
    wire N__26976;
    wire N__26975;
    wire N__26972;
    wire N__26969;
    wire N__26964;
    wire N__26961;
    wire N__26958;
    wire N__26957;
    wire N__26954;
    wire N__26951;
    wire N__26946;
    wire N__26945;
    wire N__26942;
    wire N__26941;
    wire N__26940;
    wire N__26937;
    wire N__26934;
    wire N__26931;
    wire N__26930;
    wire N__26929;
    wire N__26926;
    wire N__26923;
    wire N__26918;
    wire N__26915;
    wire N__26912;
    wire N__26909;
    wire N__26908;
    wire N__26901;
    wire N__26900;
    wire N__26897;
    wire N__26894;
    wire N__26891;
    wire N__26888;
    wire N__26885;
    wire N__26880;
    wire N__26873;
    wire N__26868;
    wire N__26865;
    wire N__26864;
    wire N__26863;
    wire N__26860;
    wire N__26857;
    wire N__26856;
    wire N__26855;
    wire N__26854;
    wire N__26853;
    wire N__26850;
    wire N__26845;
    wire N__26842;
    wire N__26839;
    wire N__26836;
    wire N__26833;
    wire N__26830;
    wire N__26827;
    wire N__26824;
    wire N__26819;
    wire N__26816;
    wire N__26813;
    wire N__26810;
    wire N__26805;
    wire N__26796;
    wire N__26793;
    wire N__26792;
    wire N__26789;
    wire N__26786;
    wire N__26781;
    wire N__26778;
    wire N__26777;
    wire N__26774;
    wire N__26771;
    wire N__26766;
    wire N__26763;
    wire N__26760;
    wire N__26759;
    wire N__26756;
    wire N__26753;
    wire N__26748;
    wire N__26745;
    wire N__26742;
    wire N__26739;
    wire N__26738;
    wire N__26735;
    wire N__26732;
    wire N__26727;
    wire N__26724;
    wire N__26721;
    wire N__26720;
    wire N__26717;
    wire N__26714;
    wire N__26709;
    wire N__26706;
    wire N__26705;
    wire N__26702;
    wire N__26699;
    wire N__26694;
    wire N__26691;
    wire N__26690;
    wire N__26687;
    wire N__26684;
    wire N__26681;
    wire N__26676;
    wire N__26673;
    wire N__26670;
    wire N__26669;
    wire N__26666;
    wire N__26663;
    wire N__26660;
    wire N__26655;
    wire N__26652;
    wire N__26649;
    wire N__26648;
    wire N__26645;
    wire N__26642;
    wire N__26639;
    wire N__26634;
    wire N__26631;
    wire N__26630;
    wire N__26627;
    wire N__26624;
    wire N__26621;
    wire N__26616;
    wire N__26613;
    wire N__26610;
    wire N__26609;
    wire N__26606;
    wire N__26603;
    wire N__26600;
    wire N__26595;
    wire N__26592;
    wire N__26589;
    wire N__26586;
    wire N__26585;
    wire N__26584;
    wire N__26581;
    wire N__26578;
    wire N__26575;
    wire N__26572;
    wire N__26565;
    wire N__26562;
    wire N__26559;
    wire N__26556;
    wire N__26553;
    wire N__26550;
    wire N__26547;
    wire N__26544;
    wire N__26541;
    wire N__26538;
    wire N__26535;
    wire N__26532;
    wire N__26529;
    wire N__26526;
    wire N__26523;
    wire N__26520;
    wire N__26517;
    wire N__26516;
    wire N__26513;
    wire N__26510;
    wire N__26505;
    wire N__26502;
    wire N__26499;
    wire N__26496;
    wire N__26493;
    wire N__26490;
    wire N__26487;
    wire N__26486;
    wire N__26485;
    wire N__26482;
    wire N__26477;
    wire N__26472;
    wire N__26469;
    wire N__26466;
    wire N__26465;
    wire N__26462;
    wire N__26461;
    wire N__26458;
    wire N__26455;
    wire N__26450;
    wire N__26445;
    wire N__26442;
    wire N__26441;
    wire N__26438;
    wire N__26435;
    wire N__26432;
    wire N__26431;
    wire N__26426;
    wire N__26423;
    wire N__26418;
    wire N__26415;
    wire N__26412;
    wire N__26409;
    wire N__26408;
    wire N__26405;
    wire N__26402;
    wire N__26401;
    wire N__26398;
    wire N__26395;
    wire N__26392;
    wire N__26385;
    wire N__26384;
    wire N__26383;
    wire N__26380;
    wire N__26375;
    wire N__26370;
    wire N__26369;
    wire N__26366;
    wire N__26365;
    wire N__26358;
    wire N__26355;
    wire N__26354;
    wire N__26351;
    wire N__26348;
    wire N__26347;
    wire N__26342;
    wire N__26339;
    wire N__26336;
    wire N__26333;
    wire N__26328;
    wire N__26327;
    wire N__26324;
    wire N__26323;
    wire N__26316;
    wire N__26313;
    wire N__26310;
    wire N__26307;
    wire N__26304;
    wire N__26301;
    wire N__26300;
    wire N__26297;
    wire N__26294;
    wire N__26291;
    wire N__26288;
    wire N__26285;
    wire N__26282;
    wire N__26281;
    wire N__26278;
    wire N__26275;
    wire N__26272;
    wire N__26265;
    wire N__26264;
    wire N__26263;
    wire N__26260;
    wire N__26255;
    wire N__26250;
    wire N__26247;
    wire N__26244;
    wire N__26241;
    wire N__26238;
    wire N__26235;
    wire N__26234;
    wire N__26231;
    wire N__26228;
    wire N__26225;
    wire N__26222;
    wire N__26221;
    wire N__26216;
    wire N__26213;
    wire N__26208;
    wire N__26207;
    wire N__26204;
    wire N__26201;
    wire N__26198;
    wire N__26195;
    wire N__26194;
    wire N__26189;
    wire N__26186;
    wire N__26181;
    wire N__26178;
    wire N__26175;
    wire N__26174;
    wire N__26173;
    wire N__26170;
    wire N__26165;
    wire N__26160;
    wire N__26157;
    wire N__26156;
    wire N__26153;
    wire N__26150;
    wire N__26147;
    wire N__26142;
    wire N__26139;
    wire N__26136;
    wire N__26133;
    wire N__26130;
    wire N__26127;
    wire N__26126;
    wire N__26123;
    wire N__26122;
    wire N__26119;
    wire N__26116;
    wire N__26113;
    wire N__26110;
    wire N__26107;
    wire N__26100;
    wire N__26097;
    wire N__26094;
    wire N__26091;
    wire N__26090;
    wire N__26087;
    wire N__26084;
    wire N__26081;
    wire N__26080;
    wire N__26077;
    wire N__26074;
    wire N__26071;
    wire N__26068;
    wire N__26061;
    wire N__26060;
    wire N__26057;
    wire N__26054;
    wire N__26051;
    wire N__26048;
    wire N__26043;
    wire N__26040;
    wire N__26037;
    wire N__26034;
    wire N__26031;
    wire N__26028;
    wire N__26025;
    wire N__26022;
    wire N__26019;
    wire N__26016;
    wire N__26013;
    wire N__26010;
    wire N__26007;
    wire N__26004;
    wire N__26003;
    wire N__26000;
    wire N__25997;
    wire N__25996;
    wire N__25993;
    wire N__25990;
    wire N__25987;
    wire N__25980;
    wire N__25977;
    wire N__25974;
    wire N__25971;
    wire N__25970;
    wire N__25969;
    wire N__25966;
    wire N__25963;
    wire N__25960;
    wire N__25957;
    wire N__25954;
    wire N__25947;
    wire N__25946;
    wire N__25943;
    wire N__25942;
    wire N__25939;
    wire N__25934;
    wire N__25929;
    wire N__25928;
    wire N__25927;
    wire N__25924;
    wire N__25919;
    wire N__25914;
    wire N__25911;
    wire N__25908;
    wire N__25907;
    wire N__25904;
    wire N__25901;
    wire N__25896;
    wire N__25893;
    wire N__25890;
    wire N__25887;
    wire N__25884;
    wire N__25881;
    wire N__25878;
    wire N__25875;
    wire N__25872;
    wire N__25869;
    wire N__25866;
    wire N__25863;
    wire N__25862;
    wire N__25861;
    wire N__25858;
    wire N__25855;
    wire N__25852;
    wire N__25845;
    wire N__25842;
    wire N__25839;
    wire N__25836;
    wire N__25833;
    wire N__25830;
    wire N__25827;
    wire N__25824;
    wire N__25821;
    wire N__25818;
    wire N__25817;
    wire N__25814;
    wire N__25811;
    wire N__25806;
    wire N__25803;
    wire N__25800;
    wire N__25799;
    wire N__25796;
    wire N__25793;
    wire N__25790;
    wire N__25787;
    wire N__25782;
    wire N__25779;
    wire N__25778;
    wire N__25775;
    wire N__25772;
    wire N__25769;
    wire N__25766;
    wire N__25763;
    wire N__25762;
    wire N__25759;
    wire N__25756;
    wire N__25753;
    wire N__25748;
    wire N__25743;
    wire N__25740;
    wire N__25739;
    wire N__25736;
    wire N__25735;
    wire N__25732;
    wire N__25729;
    wire N__25726;
    wire N__25723;
    wire N__25720;
    wire N__25717;
    wire N__25716;
    wire N__25715;
    wire N__25712;
    wire N__25709;
    wire N__25706;
    wire N__25701;
    wire N__25692;
    wire N__25689;
    wire N__25686;
    wire N__25683;
    wire N__25680;
    wire N__25677;
    wire N__25676;
    wire N__25673;
    wire N__25670;
    wire N__25667;
    wire N__25664;
    wire N__25659;
    wire N__25658;
    wire N__25655;
    wire N__25652;
    wire N__25647;
    wire N__25644;
    wire N__25643;
    wire N__25640;
    wire N__25637;
    wire N__25634;
    wire N__25631;
    wire N__25628;
    wire N__25625;
    wire N__25620;
    wire N__25619;
    wire N__25616;
    wire N__25613;
    wire N__25608;
    wire N__25605;
    wire N__25604;
    wire N__25601;
    wire N__25598;
    wire N__25595;
    wire N__25592;
    wire N__25587;
    wire N__25586;
    wire N__25583;
    wire N__25580;
    wire N__25575;
    wire N__25572;
    wire N__25571;
    wire N__25568;
    wire N__25565;
    wire N__25562;
    wire N__25559;
    wire N__25554;
    wire N__25553;
    wire N__25550;
    wire N__25549;
    wire N__25546;
    wire N__25543;
    wire N__25540;
    wire N__25535;
    wire N__25530;
    wire N__25529;
    wire N__25526;
    wire N__25525;
    wire N__25522;
    wire N__25519;
    wire N__25516;
    wire N__25513;
    wire N__25506;
    wire N__25503;
    wire N__25500;
    wire N__25497;
    wire N__25494;
    wire N__25491;
    wire N__25488;
    wire N__25487;
    wire N__25486;
    wire N__25483;
    wire N__25478;
    wire N__25475;
    wire N__25470;
    wire N__25469;
    wire N__25468;
    wire N__25465;
    wire N__25462;
    wire N__25459;
    wire N__25456;
    wire N__25449;
    wire N__25448;
    wire N__25445;
    wire N__25442;
    wire N__25437;
    wire N__25434;
    wire N__25431;
    wire N__25430;
    wire N__25427;
    wire N__25424;
    wire N__25419;
    wire N__25418;
    wire N__25415;
    wire N__25412;
    wire N__25409;
    wire N__25404;
    wire N__25401;
    wire N__25398;
    wire N__25397;
    wire N__25394;
    wire N__25391;
    wire N__25388;
    wire N__25385;
    wire N__25380;
    wire N__25379;
    wire N__25376;
    wire N__25373;
    wire N__25368;
    wire N__25365;
    wire N__25364;
    wire N__25363;
    wire N__25360;
    wire N__25357;
    wire N__25354;
    wire N__25351;
    wire N__25344;
    wire N__25343;
    wire N__25340;
    wire N__25337;
    wire N__25332;
    wire N__25329;
    wire N__25328;
    wire N__25325;
    wire N__25322;
    wire N__25317;
    wire N__25316;
    wire N__25315;
    wire N__25310;
    wire N__25307;
    wire N__25302;
    wire N__25301;
    wire N__25300;
    wire N__25297;
    wire N__25294;
    wire N__25291;
    wire N__25288;
    wire N__25281;
    wire N__25278;
    wire N__25277;
    wire N__25276;
    wire N__25273;
    wire N__25270;
    wire N__25267;
    wire N__25260;
    wire N__25259;
    wire N__25258;
    wire N__25255;
    wire N__25252;
    wire N__25249;
    wire N__25246;
    wire N__25239;
    wire N__25238;
    wire N__25235;
    wire N__25234;
    wire N__25231;
    wire N__25228;
    wire N__25225;
    wire N__25222;
    wire N__25215;
    wire N__25214;
    wire N__25213;
    wire N__25210;
    wire N__25207;
    wire N__25204;
    wire N__25201;
    wire N__25194;
    wire N__25193;
    wire N__25190;
    wire N__25189;
    wire N__25186;
    wire N__25183;
    wire N__25180;
    wire N__25177;
    wire N__25174;
    wire N__25167;
    wire N__25166;
    wire N__25165;
    wire N__25162;
    wire N__25157;
    wire N__25154;
    wire N__25149;
    wire N__25148;
    wire N__25147;
    wire N__25142;
    wire N__25139;
    wire N__25134;
    wire N__25133;
    wire N__25130;
    wire N__25127;
    wire N__25126;
    wire N__25121;
    wire N__25118;
    wire N__25115;
    wire N__25112;
    wire N__25107;
    wire N__25104;
    wire N__25101;
    wire N__25100;
    wire N__25097;
    wire N__25094;
    wire N__25089;
    wire N__25086;
    wire N__25083;
    wire N__25080;
    wire N__25077;
    wire N__25074;
    wire N__25073;
    wire N__25072;
    wire N__25069;
    wire N__25066;
    wire N__25063;
    wire N__25060;
    wire N__25057;
    wire N__25054;
    wire N__25047;
    wire N__25046;
    wire N__25045;
    wire N__25042;
    wire N__25037;
    wire N__25034;
    wire N__25029;
    wire N__25028;
    wire N__25027;
    wire N__25024;
    wire N__25019;
    wire N__25016;
    wire N__25011;
    wire N__25008;
    wire N__25005;
    wire N__25002;
    wire N__24999;
    wire N__24998;
    wire N__24993;
    wire N__24990;
    wire N__24989;
    wire N__24986;
    wire N__24983;
    wire N__24980;
    wire N__24975;
    wire N__24972;
    wire N__24969;
    wire N__24966;
    wire N__24963;
    wire N__24960;
    wire N__24957;
    wire N__24954;
    wire N__24951;
    wire N__24950;
    wire N__24945;
    wire N__24942;
    wire N__24941;
    wire N__24940;
    wire N__24939;
    wire N__24936;
    wire N__24935;
    wire N__24932;
    wire N__24929;
    wire N__24928;
    wire N__24927;
    wire N__24926;
    wire N__24919;
    wire N__24918;
    wire N__24915;
    wire N__24912;
    wire N__24909;
    wire N__24908;
    wire N__24905;
    wire N__24904;
    wire N__24903;
    wire N__24900;
    wire N__24897;
    wire N__24894;
    wire N__24891;
    wire N__24888;
    wire N__24885;
    wire N__24878;
    wire N__24875;
    wire N__24868;
    wire N__24855;
    wire N__24854;
    wire N__24853;
    wire N__24852;
    wire N__24851;
    wire N__24850;
    wire N__24847;
    wire N__24846;
    wire N__24843;
    wire N__24842;
    wire N__24841;
    wire N__24840;
    wire N__24839;
    wire N__24834;
    wire N__24829;
    wire N__24828;
    wire N__24825;
    wire N__24822;
    wire N__24819;
    wire N__24816;
    wire N__24809;
    wire N__24804;
    wire N__24801;
    wire N__24786;
    wire N__24783;
    wire N__24780;
    wire N__24777;
    wire N__24776;
    wire N__24773;
    wire N__24770;
    wire N__24767;
    wire N__24764;
    wire N__24759;
    wire N__24756;
    wire N__24753;
    wire N__24750;
    wire N__24749;
    wire N__24746;
    wire N__24743;
    wire N__24742;
    wire N__24739;
    wire N__24736;
    wire N__24733;
    wire N__24730;
    wire N__24727;
    wire N__24720;
    wire N__24717;
    wire N__24714;
    wire N__24713;
    wire N__24710;
    wire N__24707;
    wire N__24702;
    wire N__24699;
    wire N__24698;
    wire N__24693;
    wire N__24690;
    wire N__24687;
    wire N__24684;
    wire N__24681;
    wire N__24680;
    wire N__24677;
    wire N__24674;
    wire N__24669;
    wire N__24666;
    wire N__24663;
    wire N__24660;
    wire N__24659;
    wire N__24658;
    wire N__24655;
    wire N__24650;
    wire N__24645;
    wire N__24642;
    wire N__24641;
    wire N__24638;
    wire N__24635;
    wire N__24632;
    wire N__24629;
    wire N__24624;
    wire N__24623;
    wire N__24620;
    wire N__24617;
    wire N__24616;
    wire N__24615;
    wire N__24612;
    wire N__24607;
    wire N__24606;
    wire N__24603;
    wire N__24598;
    wire N__24595;
    wire N__24592;
    wire N__24587;
    wire N__24582;
    wire N__24579;
    wire N__24576;
    wire N__24573;
    wire N__24570;
    wire N__24567;
    wire N__24564;
    wire N__24561;
    wire N__24558;
    wire N__24555;
    wire N__24552;
    wire N__24549;
    wire N__24546;
    wire N__24543;
    wire N__24540;
    wire N__24537;
    wire N__24534;
    wire N__24531;
    wire N__24528;
    wire N__24525;
    wire N__24522;
    wire N__24521;
    wire N__24520;
    wire N__24517;
    wire N__24514;
    wire N__24511;
    wire N__24508;
    wire N__24505;
    wire N__24498;
    wire N__24497;
    wire N__24494;
    wire N__24493;
    wire N__24492;
    wire N__24487;
    wire N__24484;
    wire N__24481;
    wire N__24474;
    wire N__24473;
    wire N__24472;
    wire N__24467;
    wire N__24464;
    wire N__24461;
    wire N__24458;
    wire N__24453;
    wire N__24450;
    wire N__24447;
    wire N__24444;
    wire N__24441;
    wire N__24440;
    wire N__24439;
    wire N__24438;
    wire N__24437;
    wire N__24430;
    wire N__24427;
    wire N__24424;
    wire N__24417;
    wire N__24416;
    wire N__24413;
    wire N__24412;
    wire N__24409;
    wire N__24406;
    wire N__24401;
    wire N__24396;
    wire N__24393;
    wire N__24392;
    wire N__24389;
    wire N__24386;
    wire N__24381;
    wire N__24378;
    wire N__24375;
    wire N__24372;
    wire N__24369;
    wire N__24366;
    wire N__24363;
    wire N__24360;
    wire N__24357;
    wire N__24354;
    wire N__24353;
    wire N__24350;
    wire N__24347;
    wire N__24346;
    wire N__24343;
    wire N__24340;
    wire N__24337;
    wire N__24330;
    wire N__24327;
    wire N__24326;
    wire N__24323;
    wire N__24320;
    wire N__24317;
    wire N__24314;
    wire N__24313;
    wire N__24308;
    wire N__24305;
    wire N__24300;
    wire N__24297;
    wire N__24294;
    wire N__24291;
    wire N__24290;
    wire N__24287;
    wire N__24284;
    wire N__24283;
    wire N__24280;
    wire N__24277;
    wire N__24274;
    wire N__24271;
    wire N__24264;
    wire N__24261;
    wire N__24258;
    wire N__24257;
    wire N__24254;
    wire N__24253;
    wire N__24250;
    wire N__24247;
    wire N__24244;
    wire N__24237;
    wire N__24234;
    wire N__24231;
    wire N__24228;
    wire N__24227;
    wire N__24226;
    wire N__24223;
    wire N__24218;
    wire N__24213;
    wire N__24210;
    wire N__24207;
    wire N__24204;
    wire N__24201;
    wire N__24198;
    wire N__24195;
    wire N__24192;
    wire N__24191;
    wire N__24188;
    wire N__24185;
    wire N__24180;
    wire N__24177;
    wire N__24174;
    wire N__24171;
    wire N__24168;
    wire N__24165;
    wire N__24162;
    wire N__24159;
    wire N__24156;
    wire N__24155;
    wire N__24152;
    wire N__24149;
    wire N__24146;
    wire N__24143;
    wire N__24138;
    wire N__24135;
    wire N__24132;
    wire N__24131;
    wire N__24130;
    wire N__24127;
    wire N__24124;
    wire N__24121;
    wire N__24118;
    wire N__24115;
    wire N__24112;
    wire N__24109;
    wire N__24106;
    wire N__24099;
    wire N__24096;
    wire N__24093;
    wire N__24090;
    wire N__24087;
    wire N__24084;
    wire N__24081;
    wire N__24078;
    wire N__24075;
    wire N__24072;
    wire N__24069;
    wire N__24066;
    wire N__24063;
    wire N__24060;
    wire N__24057;
    wire N__24054;
    wire N__24051;
    wire N__24050;
    wire N__24047;
    wire N__24044;
    wire N__24039;
    wire N__24036;
    wire N__24033;
    wire N__24030;
    wire N__24029;
    wire N__24028;
    wire N__24025;
    wire N__24020;
    wire N__24017;
    wire N__24012;
    wire N__24009;
    wire N__24006;
    wire N__24005;
    wire N__24004;
    wire N__24001;
    wire N__23996;
    wire N__23993;
    wire N__23988;
    wire N__23985;
    wire N__23982;
    wire N__23981;
    wire N__23978;
    wire N__23975;
    wire N__23974;
    wire N__23971;
    wire N__23968;
    wire N__23965;
    wire N__23962;
    wire N__23955;
    wire N__23952;
    wire N__23949;
    wire N__23946;
    wire N__23943;
    wire N__23940;
    wire N__23937;
    wire N__23934;
    wire N__23931;
    wire N__23928;
    wire N__23925;
    wire N__23922;
    wire N__23919;
    wire N__23916;
    wire N__23913;
    wire N__23910;
    wire N__23909;
    wire N__23906;
    wire N__23903;
    wire N__23902;
    wire N__23899;
    wire N__23896;
    wire N__23893;
    wire N__23890;
    wire N__23883;
    wire N__23880;
    wire N__23877;
    wire N__23874;
    wire N__23871;
    wire N__23868;
    wire N__23865;
    wire N__23862;
    wire N__23859;
    wire N__23856;
    wire N__23853;
    wire N__23850;
    wire N__23847;
    wire N__23844;
    wire N__23841;
    wire N__23838;
    wire N__23835;
    wire N__23832;
    wire N__23831;
    wire N__23830;
    wire N__23827;
    wire N__23822;
    wire N__23819;
    wire N__23814;
    wire N__23811;
    wire N__23808;
    wire N__23805;
    wire N__23802;
    wire N__23799;
    wire N__23796;
    wire N__23793;
    wire N__23790;
    wire N__23789;
    wire N__23784;
    wire N__23781;
    wire N__23778;
    wire N__23775;
    wire N__23774;
    wire N__23769;
    wire N__23766;
    wire N__23765;
    wire N__23760;
    wire N__23757;
    wire N__23754;
    wire N__23751;
    wire N__23748;
    wire N__23745;
    wire N__23742;
    wire N__23739;
    wire N__23736;
    wire N__23733;
    wire N__23730;
    wire N__23727;
    wire N__23724;
    wire N__23723;
    wire N__23720;
    wire N__23717;
    wire N__23714;
    wire N__23711;
    wire N__23706;
    wire N__23703;
    wire N__23700;
    wire N__23697;
    wire N__23694;
    wire N__23691;
    wire N__23688;
    wire N__23685;
    wire N__23682;
    wire N__23679;
    wire N__23676;
    wire N__23673;
    wire N__23670;
    wire N__23667;
    wire N__23664;
    wire N__23661;
    wire N__23658;
    wire N__23657;
    wire N__23654;
    wire N__23651;
    wire N__23646;
    wire N__23643;
    wire N__23642;
    wire N__23637;
    wire N__23634;
    wire N__23631;
    wire N__23628;
    wire N__23625;
    wire N__23622;
    wire N__23619;
    wire N__23616;
    wire N__23613;
    wire N__23610;
    wire N__23607;
    wire N__23604;
    wire N__23601;
    wire N__23598;
    wire N__23595;
    wire N__23592;
    wire N__23589;
    wire N__23586;
    wire N__23583;
    wire N__23580;
    wire N__23577;
    wire N__23574;
    wire N__23571;
    wire N__23568;
    wire N__23565;
    wire N__23562;
    wire N__23561;
    wire N__23560;
    wire N__23557;
    wire N__23554;
    wire N__23551;
    wire N__23548;
    wire N__23545;
    wire N__23538;
    wire N__23535;
    wire N__23534;
    wire N__23531;
    wire N__23528;
    wire N__23527;
    wire N__23524;
    wire N__23519;
    wire N__23514;
    wire N__23513;
    wire N__23510;
    wire N__23509;
    wire N__23504;
    wire N__23501;
    wire N__23496;
    wire N__23493;
    wire N__23490;
    wire N__23489;
    wire N__23486;
    wire N__23483;
    wire N__23482;
    wire N__23479;
    wire N__23476;
    wire N__23473;
    wire N__23466;
    wire N__23465;
    wire N__23462;
    wire N__23461;
    wire N__23458;
    wire N__23453;
    wire N__23448;
    wire N__23447;
    wire N__23444;
    wire N__23443;
    wire N__23438;
    wire N__23435;
    wire N__23432;
    wire N__23429;
    wire N__23424;
    wire N__23423;
    wire N__23420;
    wire N__23417;
    wire N__23416;
    wire N__23413;
    wire N__23408;
    wire N__23403;
    wire N__23400;
    wire N__23397;
    wire N__23394;
    wire N__23391;
    wire N__23388;
    wire N__23385;
    wire N__23382;
    wire N__23379;
    wire N__23376;
    wire N__23373;
    wire N__23370;
    wire N__23367;
    wire N__23364;
    wire N__23361;
    wire N__23358;
    wire N__23355;
    wire N__23352;
    wire N__23349;
    wire N__23348;
    wire N__23345;
    wire N__23342;
    wire N__23337;
    wire N__23334;
    wire N__23331;
    wire N__23330;
    wire N__23327;
    wire N__23324;
    wire N__23323;
    wire N__23320;
    wire N__23315;
    wire N__23314;
    wire N__23313;
    wire N__23308;
    wire N__23303;
    wire N__23298;
    wire N__23297;
    wire N__23294;
    wire N__23291;
    wire N__23288;
    wire N__23285;
    wire N__23284;
    wire N__23281;
    wire N__23278;
    wire N__23275;
    wire N__23268;
    wire N__23265;
    wire N__23262;
    wire N__23259;
    wire N__23258;
    wire N__23257;
    wire N__23254;
    wire N__23251;
    wire N__23248;
    wire N__23245;
    wire N__23242;
    wire N__23235;
    wire N__23232;
    wire N__23229;
    wire N__23228;
    wire N__23227;
    wire N__23224;
    wire N__23221;
    wire N__23218;
    wire N__23215;
    wire N__23212;
    wire N__23209;
    wire N__23202;
    wire N__23201;
    wire N__23200;
    wire N__23197;
    wire N__23194;
    wire N__23191;
    wire N__23184;
    wire N__23181;
    wire N__23178;
    wire N__23175;
    wire N__23172;
    wire N__23169;
    wire N__23166;
    wire N__23163;
    wire N__23160;
    wire N__23159;
    wire N__23158;
    wire N__23155;
    wire N__23150;
    wire N__23145;
    wire N__23142;
    wire N__23139;
    wire N__23138;
    wire N__23137;
    wire N__23134;
    wire N__23131;
    wire N__23128;
    wire N__23125;
    wire N__23122;
    wire N__23117;
    wire N__23114;
    wire N__23109;
    wire N__23106;
    wire N__23103;
    wire N__23100;
    wire N__23099;
    wire N__23096;
    wire N__23093;
    wire N__23092;
    wire N__23089;
    wire N__23086;
    wire N__23083;
    wire N__23080;
    wire N__23073;
    wire N__23070;
    wire N__23067;
    wire N__23064;
    wire N__23061;
    wire N__23060;
    wire N__23057;
    wire N__23054;
    wire N__23053;
    wire N__23050;
    wire N__23047;
    wire N__23044;
    wire N__23037;
    wire N__23034;
    wire N__23031;
    wire N__23030;
    wire N__23027;
    wire N__23024;
    wire N__23023;
    wire N__23020;
    wire N__23015;
    wire N__23010;
    wire N__23009;
    wire N__23008;
    wire N__23007;
    wire N__23006;
    wire N__23005;
    wire N__23002;
    wire N__22999;
    wire N__22998;
    wire N__22995;
    wire N__22992;
    wire N__22989;
    wire N__22980;
    wire N__22971;
    wire N__22970;
    wire N__22969;
    wire N__22968;
    wire N__22967;
    wire N__22964;
    wire N__22961;
    wire N__22960;
    wire N__22957;
    wire N__22954;
    wire N__22951;
    wire N__22950;
    wire N__22949;
    wire N__22948;
    wire N__22945;
    wire N__22942;
    wire N__22939;
    wire N__22936;
    wire N__22925;
    wire N__22916;
    wire N__22913;
    wire N__22910;
    wire N__22907;
    wire N__22902;
    wire N__22901;
    wire N__22898;
    wire N__22895;
    wire N__22892;
    wire N__22887;
    wire N__22886;
    wire N__22883;
    wire N__22880;
    wire N__22875;
    wire N__22874;
    wire N__22871;
    wire N__22868;
    wire N__22865;
    wire N__22862;
    wire N__22857;
    wire N__22854;
    wire N__22853;
    wire N__22850;
    wire N__22847;
    wire N__22846;
    wire N__22843;
    wire N__22840;
    wire N__22837;
    wire N__22834;
    wire N__22831;
    wire N__22824;
    wire N__22821;
    wire N__22818;
    wire N__22815;
    wire N__22814;
    wire N__22811;
    wire N__22808;
    wire N__22803;
    wire N__22800;
    wire N__22799;
    wire N__22796;
    wire N__22793;
    wire N__22792;
    wire N__22789;
    wire N__22786;
    wire N__22783;
    wire N__22780;
    wire N__22773;
    wire N__22770;
    wire N__22767;
    wire N__22766;
    wire N__22763;
    wire N__22760;
    wire N__22755;
    wire N__22754;
    wire N__22749;
    wire N__22746;
    wire N__22743;
    wire N__22740;
    wire N__22739;
    wire N__22734;
    wire N__22731;
    wire N__22730;
    wire N__22725;
    wire N__22722;
    wire N__22721;
    wire N__22716;
    wire N__22713;
    wire N__22710;
    wire N__22707;
    wire N__22706;
    wire N__22703;
    wire N__22700;
    wire N__22695;
    wire N__22694;
    wire N__22693;
    wire N__22692;
    wire N__22691;
    wire N__22688;
    wire N__22687;
    wire N__22686;
    wire N__22685;
    wire N__22684;
    wire N__22683;
    wire N__22680;
    wire N__22679;
    wire N__22678;
    wire N__22677;
    wire N__22674;
    wire N__22671;
    wire N__22670;
    wire N__22663;
    wire N__22660;
    wire N__22653;
    wire N__22652;
    wire N__22649;
    wire N__22646;
    wire N__22645;
    wire N__22644;
    wire N__22641;
    wire N__22640;
    wire N__22639;
    wire N__22636;
    wire N__22635;
    wire N__22632;
    wire N__22627;
    wire N__22620;
    wire N__22617;
    wire N__22614;
    wire N__22611;
    wire N__22610;
    wire N__22609;
    wire N__22606;
    wire N__22605;
    wire N__22604;
    wire N__22603;
    wire N__22600;
    wire N__22597;
    wire N__22594;
    wire N__22587;
    wire N__22580;
    wire N__22573;
    wire N__22560;
    wire N__22545;
    wire N__22544;
    wire N__22541;
    wire N__22538;
    wire N__22535;
    wire N__22532;
    wire N__22527;
    wire N__22526;
    wire N__22523;
    wire N__22520;
    wire N__22517;
    wire N__22516;
    wire N__22513;
    wire N__22512;
    wire N__22509;
    wire N__22506;
    wire N__22503;
    wire N__22500;
    wire N__22491;
    wire N__22488;
    wire N__22487;
    wire N__22484;
    wire N__22481;
    wire N__22476;
    wire N__22473;
    wire N__22470;
    wire N__22469;
    wire N__22464;
    wire N__22461;
    wire N__22458;
    wire N__22455;
    wire N__22452;
    wire N__22449;
    wire N__22446;
    wire N__22443;
    wire N__22440;
    wire N__22437;
    wire N__22434;
    wire N__22431;
    wire N__22428;
    wire N__22425;
    wire N__22422;
    wire N__22421;
    wire N__22418;
    wire N__22415;
    wire N__22414;
    wire N__22413;
    wire N__22412;
    wire N__22411;
    wire N__22410;
    wire N__22409;
    wire N__22406;
    wire N__22405;
    wire N__22404;
    wire N__22403;
    wire N__22402;
    wire N__22401;
    wire N__22400;
    wire N__22399;
    wire N__22398;
    wire N__22383;
    wire N__22380;
    wire N__22379;
    wire N__22378;
    wire N__22377;
    wire N__22376;
    wire N__22375;
    wire N__22370;
    wire N__22361;
    wire N__22356;
    wire N__22353;
    wire N__22352;
    wire N__22351;
    wire N__22350;
    wire N__22347;
    wire N__22344;
    wire N__22343;
    wire N__22342;
    wire N__22341;
    wire N__22340;
    wire N__22339;
    wire N__22338;
    wire N__22337;
    wire N__22336;
    wire N__22333;
    wire N__22332;
    wire N__22331;
    wire N__22328;
    wire N__22327;
    wire N__22324;
    wire N__22321;
    wire N__22314;
    wire N__22311;
    wire N__22308;
    wire N__22305;
    wire N__22302;
    wire N__22297;
    wire N__22284;
    wire N__22269;
    wire N__22262;
    wire N__22257;
    wire N__22242;
    wire N__22239;
    wire N__22236;
    wire N__22235;
    wire N__22232;
    wire N__22229;
    wire N__22224;
    wire N__22223;
    wire N__22222;
    wire N__22221;
    wire N__22220;
    wire N__22219;
    wire N__22218;
    wire N__22217;
    wire N__22216;
    wire N__22215;
    wire N__22198;
    wire N__22197;
    wire N__22196;
    wire N__22195;
    wire N__22194;
    wire N__22193;
    wire N__22192;
    wire N__22189;
    wire N__22188;
    wire N__22187;
    wire N__22186;
    wire N__22183;
    wire N__22182;
    wire N__22181;
    wire N__22180;
    wire N__22179;
    wire N__22178;
    wire N__22177;
    wire N__22176;
    wire N__22175;
    wire N__22174;
    wire N__22173;
    wire N__22170;
    wire N__22169;
    wire N__22168;
    wire N__22157;
    wire N__22156;
    wire N__22155;
    wire N__22154;
    wire N__22153;
    wire N__22152;
    wire N__22149;
    wire N__22146;
    wire N__22141;
    wire N__22138;
    wire N__22135;
    wire N__22130;
    wire N__22125;
    wire N__22116;
    wire N__22115;
    wire N__22112;
    wire N__22111;
    wire N__22108;
    wire N__22105;
    wire N__22102;
    wire N__22099;
    wire N__22098;
    wire N__22097;
    wire N__22096;
    wire N__22095;
    wire N__22094;
    wire N__22091;
    wire N__22080;
    wire N__22077;
    wire N__22074;
    wire N__22069;
    wire N__22068;
    wire N__22067;
    wire N__22066;
    wire N__22063;
    wire N__22058;
    wire N__22055;
    wire N__22052;
    wire N__22047;
    wire N__22044;
    wire N__22039;
    wire N__22034;
    wire N__22025;
    wire N__22014;
    wire N__22007;
    wire N__22000;
    wire N__21981;
    wire N__21978;
    wire N__21975;
    wire N__21972;
    wire N__21969;
    wire N__21966;
    wire N__21963;
    wire N__21962;
    wire N__21959;
    wire N__21956;
    wire N__21953;
    wire N__21948;
    wire N__21945;
    wire N__21942;
    wire N__21941;
    wire N__21938;
    wire N__21935;
    wire N__21930;
    wire N__21927;
    wire N__21924;
    wire N__21921;
    wire N__21918;
    wire N__21915;
    wire N__21912;
    wire N__21909;
    wire N__21906;
    wire N__21903;
    wire N__21900;
    wire N__21897;
    wire N__21894;
    wire N__21891;
    wire N__21888;
    wire N__21885;
    wire N__21882;
    wire N__21879;
    wire N__21876;
    wire N__21873;
    wire N__21870;
    wire N__21869;
    wire N__21866;
    wire N__21863;
    wire N__21858;
    wire N__21855;
    wire N__21852;
    wire N__21849;
    wire N__21846;
    wire N__21843;
    wire N__21840;
    wire N__21837;
    wire N__21834;
    wire N__21831;
    wire N__21830;
    wire N__21827;
    wire N__21824;
    wire N__21819;
    wire N__21816;
    wire N__21815;
    wire N__21812;
    wire N__21809;
    wire N__21804;
    wire N__21801;
    wire N__21800;
    wire N__21797;
    wire N__21794;
    wire N__21789;
    wire N__21786;
    wire N__21785;
    wire N__21782;
    wire N__21779;
    wire N__21774;
    wire N__21771;
    wire N__21770;
    wire N__21767;
    wire N__21764;
    wire N__21759;
    wire N__21756;
    wire N__21755;
    wire N__21752;
    wire N__21749;
    wire N__21746;
    wire N__21741;
    wire N__21738;
    wire N__21735;
    wire N__21732;
    wire N__21729;
    wire N__21726;
    wire N__21723;
    wire N__21722;
    wire N__21719;
    wire N__21716;
    wire N__21715;
    wire N__21714;
    wire N__21713;
    wire N__21710;
    wire N__21707;
    wire N__21704;
    wire N__21701;
    wire N__21698;
    wire N__21695;
    wire N__21692;
    wire N__21689;
    wire N__21686;
    wire N__21683;
    wire N__21678;
    wire N__21671;
    wire N__21666;
    wire N__21663;
    wire N__21660;
    wire N__21657;
    wire N__21654;
    wire N__21651;
    wire N__21650;
    wire N__21647;
    wire N__21644;
    wire N__21641;
    wire N__21638;
    wire N__21633;
    wire N__21630;
    wire N__21627;
    wire N__21626;
    wire N__21625;
    wire N__21622;
    wire N__21621;
    wire N__21620;
    wire N__21619;
    wire N__21618;
    wire N__21617;
    wire N__21616;
    wire N__21613;
    wire N__21612;
    wire N__21609;
    wire N__21608;
    wire N__21607;
    wire N__21604;
    wire N__21601;
    wire N__21598;
    wire N__21595;
    wire N__21592;
    wire N__21587;
    wire N__21576;
    wire N__21569;
    wire N__21558;
    wire N__21557;
    wire N__21556;
    wire N__21555;
    wire N__21554;
    wire N__21553;
    wire N__21552;
    wire N__21547;
    wire N__21544;
    wire N__21543;
    wire N__21542;
    wire N__21541;
    wire N__21540;
    wire N__21539;
    wire N__21536;
    wire N__21533;
    wire N__21528;
    wire N__21523;
    wire N__21512;
    wire N__21501;
    wire N__21498;
    wire N__21497;
    wire N__21496;
    wire N__21493;
    wire N__21490;
    wire N__21487;
    wire N__21484;
    wire N__21479;
    wire N__21474;
    wire N__21471;
    wire N__21468;
    wire N__21465;
    wire N__21462;
    wire N__21459;
    wire N__21458;
    wire N__21455;
    wire N__21452;
    wire N__21449;
    wire N__21446;
    wire N__21441;
    wire N__21440;
    wire N__21437;
    wire N__21436;
    wire N__21429;
    wire N__21426;
    wire N__21423;
    wire N__21420;
    wire N__21417;
    wire N__21416;
    wire N__21413;
    wire N__21410;
    wire N__21405;
    wire N__21402;
    wire N__21399;
    wire N__21398;
    wire N__21395;
    wire N__21394;
    wire N__21391;
    wire N__21388;
    wire N__21385;
    wire N__21378;
    wire N__21377;
    wire N__21374;
    wire N__21371;
    wire N__21368;
    wire N__21367;
    wire N__21364;
    wire N__21361;
    wire N__21358;
    wire N__21351;
    wire N__21348;
    wire N__21345;
    wire N__21342;
    wire N__21339;
    wire N__21336;
    wire N__21333;
    wire N__21330;
    wire N__21329;
    wire N__21328;
    wire N__21323;
    wire N__21320;
    wire N__21315;
    wire N__21314;
    wire N__21311;
    wire N__21308;
    wire N__21307;
    wire N__21304;
    wire N__21301;
    wire N__21298;
    wire N__21295;
    wire N__21288;
    wire N__21287;
    wire N__21284;
    wire N__21281;
    wire N__21278;
    wire N__21277;
    wire N__21274;
    wire N__21271;
    wire N__21268;
    wire N__21261;
    wire N__21258;
    wire N__21255;
    wire N__21252;
    wire N__21249;
    wire N__21246;
    wire N__21243;
    wire N__21240;
    wire N__21237;
    wire N__21236;
    wire N__21233;
    wire N__21230;
    wire N__21225;
    wire N__21222;
    wire N__21219;
    wire N__21218;
    wire N__21215;
    wire N__21212;
    wire N__21211;
    wire N__21206;
    wire N__21203;
    wire N__21198;
    wire N__21197;
    wire N__21196;
    wire N__21193;
    wire N__21190;
    wire N__21187;
    wire N__21184;
    wire N__21179;
    wire N__21174;
    wire N__21173;
    wire N__21170;
    wire N__21169;
    wire N__21166;
    wire N__21165;
    wire N__21164;
    wire N__21163;
    wire N__21162;
    wire N__21161;
    wire N__21156;
    wire N__21155;
    wire N__21154;
    wire N__21153;
    wire N__21152;
    wire N__21151;
    wire N__21150;
    wire N__21149;
    wire N__21142;
    wire N__21137;
    wire N__21134;
    wire N__21131;
    wire N__21126;
    wire N__21115;
    wire N__21102;
    wire N__21101;
    wire N__21100;
    wire N__21097;
    wire N__21092;
    wire N__21089;
    wire N__21084;
    wire N__21083;
    wire N__21082;
    wire N__21079;
    wire N__21074;
    wire N__21069;
    wire N__21068;
    wire N__21067;
    wire N__21064;
    wire N__21061;
    wire N__21058;
    wire N__21055;
    wire N__21050;
    wire N__21045;
    wire N__21044;
    wire N__21043;
    wire N__21042;
    wire N__21041;
    wire N__21040;
    wire N__21039;
    wire N__21038;
    wire N__21035;
    wire N__21032;
    wire N__21031;
    wire N__21030;
    wire N__21029;
    wire N__21028;
    wire N__21027;
    wire N__21026;
    wire N__21025;
    wire N__21018;
    wire N__21011;
    wire N__21008;
    wire N__21005;
    wire N__20996;
    wire N__20989;
    wire N__20976;
    wire N__20975;
    wire N__20974;
    wire N__20971;
    wire N__20970;
    wire N__20969;
    wire N__20968;
    wire N__20965;
    wire N__20962;
    wire N__20961;
    wire N__20960;
    wire N__20959;
    wire N__20952;
    wire N__20951;
    wire N__20950;
    wire N__20949;
    wire N__20946;
    wire N__20935;
    wire N__20932;
    wire N__20925;
    wire N__20924;
    wire N__20923;
    wire N__20922;
    wire N__20921;
    wire N__20918;
    wire N__20915;
    wire N__20910;
    wire N__20903;
    wire N__20900;
    wire N__20895;
    wire N__20892;
    wire N__20887;
    wire N__20880;
    wire N__20877;
    wire N__20876;
    wire N__20873;
    wire N__20872;
    wire N__20869;
    wire N__20866;
    wire N__20863;
    wire N__20856;
    wire N__20855;
    wire N__20854;
    wire N__20851;
    wire N__20846;
    wire N__20841;
    wire N__20838;
    wire N__20835;
    wire N__20834;
    wire N__20831;
    wire N__20830;
    wire N__20827;
    wire N__20824;
    wire N__20821;
    wire N__20814;
    wire N__20811;
    wire N__20810;
    wire N__20807;
    wire N__20804;
    wire N__20801;
    wire N__20798;
    wire N__20795;
    wire N__20790;
    wire N__20787;
    wire N__20786;
    wire N__20783;
    wire N__20780;
    wire N__20775;
    wire N__20774;
    wire N__20771;
    wire N__20768;
    wire N__20767;
    wire N__20764;
    wire N__20759;
    wire N__20754;
    wire N__20753;
    wire N__20752;
    wire N__20751;
    wire N__20750;
    wire N__20749;
    wire N__20748;
    wire N__20745;
    wire N__20744;
    wire N__20743;
    wire N__20742;
    wire N__20735;
    wire N__20730;
    wire N__20729;
    wire N__20728;
    wire N__20727;
    wire N__20726;
    wire N__20725;
    wire N__20718;
    wire N__20713;
    wire N__20712;
    wire N__20711;
    wire N__20706;
    wire N__20697;
    wire N__20694;
    wire N__20691;
    wire N__20688;
    wire N__20687;
    wire N__20686;
    wire N__20685;
    wire N__20680;
    wire N__20679;
    wire N__20674;
    wire N__20673;
    wire N__20672;
    wire N__20671;
    wire N__20666;
    wire N__20663;
    wire N__20656;
    wire N__20653;
    wire N__20650;
    wire N__20647;
    wire N__20640;
    wire N__20625;
    wire N__20622;
    wire N__20619;
    wire N__20616;
    wire N__20613;
    wire N__20610;
    wire N__20609;
    wire N__20608;
    wire N__20605;
    wire N__20602;
    wire N__20599;
    wire N__20592;
    wire N__20589;
    wire N__20586;
    wire N__20583;
    wire N__20582;
    wire N__20581;
    wire N__20580;
    wire N__20579;
    wire N__20576;
    wire N__20571;
    wire N__20566;
    wire N__20559;
    wire N__20556;
    wire N__20555;
    wire N__20554;
    wire N__20551;
    wire N__20548;
    wire N__20545;
    wire N__20538;
    wire N__20535;
    wire N__20534;
    wire N__20531;
    wire N__20528;
    wire N__20525;
    wire N__20522;
    wire N__20517;
    wire N__20516;
    wire N__20513;
    wire N__20510;
    wire N__20507;
    wire N__20502;
    wire N__20499;
    wire N__20496;
    wire N__20495;
    wire N__20494;
    wire N__20491;
    wire N__20488;
    wire N__20485;
    wire N__20482;
    wire N__20479;
    wire N__20476;
    wire N__20469;
    wire N__20466;
    wire N__20463;
    wire N__20460;
    wire N__20457;
    wire N__20454;
    wire N__20451;
    wire N__20450;
    wire N__20447;
    wire N__20444;
    wire N__20441;
    wire N__20438;
    wire N__20435;
    wire N__20430;
    wire N__20429;
    wire N__20428;
    wire N__20427;
    wire N__20424;
    wire N__20419;
    wire N__20416;
    wire N__20409;
    wire N__20406;
    wire N__20403;
    wire N__20400;
    wire N__20397;
    wire N__20394;
    wire N__20393;
    wire N__20392;
    wire N__20391;
    wire N__20390;
    wire N__20389;
    wire N__20388;
    wire N__20385;
    wire N__20372;
    wire N__20367;
    wire N__20364;
    wire N__20361;
    wire N__20358;
    wire N__20355;
    wire N__20352;
    wire N__20349;
    wire N__20346;
    wire N__20345;
    wire N__20342;
    wire N__20339;
    wire N__20336;
    wire N__20333;
    wire N__20330;
    wire N__20327;
    wire N__20322;
    wire N__20319;
    wire N__20316;
    wire N__20313;
    wire N__20310;
    wire N__20307;
    wire N__20304;
    wire N__20301;
    wire N__20298;
    wire N__20295;
    wire N__20292;
    wire N__20289;
    wire N__20286;
    wire N__20283;
    wire N__20280;
    wire N__20279;
    wire N__20276;
    wire N__20273;
    wire N__20268;
    wire N__20265;
    wire N__20262;
    wire N__20259;
    wire N__20256;
    wire N__20253;
    wire N__20250;
    wire N__20249;
    wire N__20246;
    wire N__20243;
    wire N__20238;
    wire N__20237;
    wire N__20234;
    wire N__20231;
    wire N__20226;
    wire N__20225;
    wire N__20222;
    wire N__20219;
    wire N__20216;
    wire N__20211;
    wire N__20210;
    wire N__20207;
    wire N__20204;
    wire N__20199;
    wire N__20198;
    wire N__20195;
    wire N__20192;
    wire N__20189;
    wire N__20184;
    wire N__20183;
    wire N__20180;
    wire N__20177;
    wire N__20172;
    wire N__20169;
    wire N__20168;
    wire N__20165;
    wire N__20162;
    wire N__20157;
    wire N__20156;
    wire N__20153;
    wire N__20150;
    wire N__20145;
    wire N__20142;
    wire N__20139;
    wire N__20138;
    wire N__20135;
    wire N__20132;
    wire N__20127;
    wire N__20124;
    wire N__20121;
    wire N__20118;
    wire N__20115;
    wire N__20112;
    wire N__20111;
    wire N__20106;
    wire N__20103;
    wire N__20100;
    wire N__20097;
    wire N__20094;
    wire N__20091;
    wire N__20088;
    wire N__20085;
    wire N__20084;
    wire N__20079;
    wire N__20076;
    wire N__20073;
    wire N__20072;
    wire N__20067;
    wire N__20064;
    wire N__20063;
    wire N__20058;
    wire N__20055;
    wire N__20052;
    wire N__20049;
    wire N__20046;
    wire N__20043;
    wire N__20040;
    wire N__20037;
    wire N__20034;
    wire N__20033;
    wire N__20032;
    wire N__20029;
    wire N__20024;
    wire N__20019;
    wire N__20018;
    wire N__20017;
    wire N__20014;
    wire N__20011;
    wire N__20004;
    wire N__20001;
    wire N__20000;
    wire N__19999;
    wire N__19996;
    wire N__19993;
    wire N__19988;
    wire N__19985;
    wire N__19982;
    wire N__19977;
    wire N__19974;
    wire N__19973;
    wire N__19972;
    wire N__19969;
    wire N__19964;
    wire N__19959;
    wire N__19958;
    wire N__19955;
    wire N__19954;
    wire N__19951;
    wire N__19948;
    wire N__19943;
    wire N__19938;
    wire N__19935;
    wire N__19932;
    wire N__19931;
    wire N__19930;
    wire N__19927;
    wire N__19922;
    wire N__19917;
    wire N__19914;
    wire N__19911;
    wire N__19910;
    wire N__19905;
    wire N__19902;
    wire N__19899;
    wire N__19898;
    wire N__19897;
    wire N__19894;
    wire N__19889;
    wire N__19886;
    wire N__19881;
    wire N__19878;
    wire N__19875;
    wire N__19872;
    wire N__19869;
    wire N__19868;
    wire N__19867;
    wire N__19866;
    wire N__19863;
    wire N__19858;
    wire N__19855;
    wire N__19852;
    wire N__19847;
    wire N__19844;
    wire N__19839;
    wire N__19838;
    wire N__19833;
    wire N__19830;
    wire N__19827;
    wire N__19824;
    wire N__19821;
    wire N__19818;
    wire N__19815;
    wire N__19812;
    wire N__19809;
    wire N__19806;
    wire N__19803;
    wire N__19800;
    wire N__19797;
    wire N__19796;
    wire N__19795;
    wire N__19792;
    wire N__19789;
    wire N__19788;
    wire N__19787;
    wire N__19786;
    wire N__19783;
    wire N__19772;
    wire N__19767;
    wire N__19764;
    wire N__19761;
    wire N__19758;
    wire N__19755;
    wire N__19752;
    wire N__19749;
    wire N__19746;
    wire N__19743;
    wire N__19740;
    wire N__19737;
    wire N__19734;
    wire N__19733;
    wire N__19730;
    wire N__19727;
    wire N__19722;
    wire N__19719;
    wire N__19718;
    wire N__19713;
    wire N__19710;
    wire N__19707;
    wire N__19706;
    wire N__19701;
    wire N__19698;
    wire N__19695;
    wire N__19694;
    wire N__19689;
    wire N__19686;
    wire N__19683;
    wire N__19680;
    wire N__19677;
    wire N__19674;
    wire N__19671;
    wire N__19668;
    wire N__19665;
    wire N__19662;
    wire N__19661;
    wire N__19658;
    wire N__19655;
    wire N__19650;
    wire N__19647;
    wire N__19644;
    wire N__19643;
    wire N__19640;
    wire N__19637;
    wire N__19632;
    wire N__19629;
    wire N__19626;
    wire N__19623;
    wire N__19620;
    wire N__19617;
    wire N__19614;
    wire N__19613;
    wire N__19612;
    wire N__19607;
    wire N__19604;
    wire N__19599;
    wire N__19598;
    wire N__19597;
    wire N__19596;
    wire N__19589;
    wire N__19586;
    wire N__19581;
    wire N__19580;
    wire N__19579;
    wire N__19578;
    wire N__19577;
    wire N__19568;
    wire N__19565;
    wire N__19560;
    wire N__19557;
    wire N__19554;
    wire N__19551;
    wire N__19548;
    wire N__19545;
    wire N__19542;
    wire N__19539;
    wire N__19536;
    wire N__19533;
    wire N__19530;
    wire N__19527;
    wire N__19524;
    wire N__19521;
    wire N__19518;
    wire N__19515;
    wire N__19512;
    wire N__19511;
    wire N__19510;
    wire N__19509;
    wire N__19508;
    wire N__19501;
    wire N__19496;
    wire N__19491;
    wire N__19490;
    wire N__19487;
    wire N__19484;
    wire N__19479;
    wire N__19478;
    wire N__19477;
    wire N__19474;
    wire N__19471;
    wire N__19468;
    wire N__19461;
    wire N__19458;
    wire N__19457;
    wire N__19456;
    wire N__19455;
    wire N__19450;
    wire N__19447;
    wire N__19444;
    wire N__19437;
    wire N__19434;
    wire N__19431;
    wire N__19428;
    wire N__19425;
    wire N__19422;
    wire N__19419;
    wire N__19416;
    wire N__19413;
    wire N__19410;
    wire N__19407;
    wire N__19404;
    wire N__19401;
    wire N__19398;
    wire N__19395;
    wire N__19392;
    wire N__19389;
    wire N__19386;
    wire N__19383;
    wire N__19380;
    wire ICE_GPMO_2;
    wire VCCG0;
    wire INViac_raw_buf_vac_raw_buf_merged11WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged3WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged10WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged8WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged4WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged9WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged5WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged0WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged6WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged1WCLKN_net;
    wire ICE_SYSCLK;
    wire INViac_raw_buf_vac_raw_buf_merged7WCLKN_net;
    wire INViac_raw_buf_vac_raw_buf_merged2WCLKN_net;
    wire \RTD.n18092 ;
    wire RTD_SCLK;
    wire \CLK_DDS.n16974 ;
    wire bit_cnt_0_adj_1498;
    wire bit_cnt_3;
    wire bit_cnt_2;
    wire bit_cnt_1;
    wire n8_adj_1680_cascade_;
    wire n21625;
    wire \RTD.n18043_cascade_ ;
    wire \RTD.n21494 ;
    wire \RTD.n21492_cascade_ ;
    wire \RTD.n7_adj_1435 ;
    wire \RTD.bit_cnt_2 ;
    wire \RTD.bit_cnt_1 ;
    wire \RTD.bit_cnt_0 ;
    wire RTD_SDI;
    wire \RTD.n21471_cascade_ ;
    wire \RTD.n19032 ;
    wire \RTD.n4_cascade_ ;
    wire \RTD.n21387 ;
    wire \RTD.n21199_cascade_ ;
    wire \RTD.adc_state_3_N_1114_1 ;
    wire \RTD.n7_cascade_ ;
    wire \RTD.n11868 ;
    wire \RTD.n11860 ;
    wire \RTD.n8 ;
    wire adress_1;
    wire adress_2;
    wire adress_3;
    wire adress_4;
    wire adress_5;
    wire RTD_SDO;
    wire \RTD.n11915 ;
    wire n14692;
    wire \RTD.n15280 ;
    wire read_buf_10;
    wire n13212_cascade_;
    wire read_buf_15;
    wire n11856_cascade_;
    wire read_buf_14;
    wire \RTD.n12_adj_1445 ;
    wire \RTD.mode ;
    wire read_buf_4;
    wire read_buf_11;
    wire read_buf_5;
    wire read_buf_3;
    wire n19_adj_1600_cascade_;
    wire n19_adj_1597_cascade_;
    wire buf_adcdata_vac_7;
    wire cmd_rdadctmp_7_adj_1485;
    wire VAC_MISO;
    wire cmd_rdadctmp_0_adj_1492;
    wire cmd_rdadctmp_1_adj_1491;
    wire cmd_rdadctmp_2_adj_1490;
    wire bfn_5_14_0_;
    wire \ADC_VAC.n19835 ;
    wire \ADC_VAC.n19836 ;
    wire \ADC_VAC.n19837 ;
    wire \ADC_VAC.n19838 ;
    wire \ADC_VAC.n19839 ;
    wire \ADC_VAC.n19840 ;
    wire \ADC_VAC.n19841 ;
    wire \ADC_VAC.bit_cnt_4 ;
    wire \ADC_VAC.bit_cnt_3 ;
    wire \ADC_VAC.bit_cnt_1 ;
    wire \ADC_VAC.bit_cnt_2 ;
    wire \ADC_VAC.bit_cnt_6 ;
    wire \ADC_VAC.bit_cnt_0 ;
    wire \ADC_VAC.n21224_cascade_ ;
    wire \ADC_VAC.bit_cnt_7 ;
    wire \ADC_VAC.bit_cnt_5 ;
    wire \ADC_VAC.n21234_cascade_ ;
    wire \ADC_VAC.n12803 ;
    wire \ADC_VAC.n15052 ;
    wire \ADC_VAC.n21157_cascade_ ;
    wire \ADC_VAC.n21468 ;
    wire \ADC_VAC.n21158 ;
    wire \RTD.n16766 ;
    wire RTD_CS;
    wire \RTD.n14 ;
    wire \RTD.n21181_cascade_ ;
    wire \RTD.n13137_cascade_ ;
    wire \RTD.n7889 ;
    wire \RTD.bit_cnt_3 ;
    wire \RTD.n18043 ;
    wire \RTD.n19026 ;
    wire adress_6;
    wire \RTD.n9_cascade_ ;
    wire \RTD.adress_7_N_1086_7_cascade_ ;
    wire RTD_DRDY;
    wire \RTD.n11_cascade_ ;
    wire \RTD.n19_cascade_ ;
    wire \RTD.adress_7 ;
    wire \RTD.adress_7_N_1086_7 ;
    wire adress_0;
    wire n13054;
    wire \RTD.n20370 ;
    wire \RTD.cfg_buf_6 ;
    wire read_buf_9;
    wire \RTD.adc_state_1 ;
    wire \RTD.n11829 ;
    wire read_buf_8;
    wire read_buf_0;
    wire read_buf_2;
    wire n11856;
    wire read_buf_1;
    wire read_buf_12;
    wire read_buf_13;
    wire n13212;
    wire n1_adj_1592;
    wire read_buf_6;
    wire read_buf_7;
    wire buf_adcdata_iac_6;
    wire buf_adcdata_vac_4;
    wire n19_adj_1606_cascade_;
    wire buf_data_iac_4;
    wire n22_adj_1607_cascade_;
    wire cmd_rdadctmp_31_adj_1461;
    wire buf_adcdata_iac_7;
    wire cmd_rdadctmp_8_adj_1484;
    wire buf_data_iac_7;
    wire n22_adj_1598;
    wire cmd_rdadctmp_12_adj_1480;
    wire buf_adcdata_iac_4;
    wire \ADC_VAC.n17 ;
    wire VAC_SCLK;
    wire cmd_rdadctmp_26_adj_1466;
    wire cmd_rdadctmp_3_adj_1489;
    wire \ADC_VAC.n12 ;
    wire n21050;
    wire VAC_DRDY;
    wire n21050_cascade_;
    wire VAC_CS;
    wire n14_adj_1657;
    wire DTRIG_N_958_adj_1493;
    wire adc_state_1_adj_1459;
    wire cmd_rdadctmp_14;
    wire \ADC_IAC.n21458_cascade_ ;
    wire \ADC_IAC.n16 ;
    wire \ADC_IAC.bit_cnt_0 ;
    wire bfn_6_18_0_;
    wire \ADC_IAC.bit_cnt_1 ;
    wire \ADC_IAC.n19828 ;
    wire \ADC_IAC.bit_cnt_2 ;
    wire \ADC_IAC.n19829 ;
    wire \ADC_IAC.bit_cnt_3 ;
    wire \ADC_IAC.n19830 ;
    wire \ADC_IAC.bit_cnt_4 ;
    wire \ADC_IAC.n19831 ;
    wire \ADC_IAC.bit_cnt_5 ;
    wire \ADC_IAC.n19832 ;
    wire \ADC_IAC.bit_cnt_6 ;
    wire \ADC_IAC.n19833 ;
    wire \ADC_IAC.n19834 ;
    wire \ADC_IAC.bit_cnt_7 ;
    wire \ADC_IAC.n12698 ;
    wire \ADC_IAC.n12698_cascade_ ;
    wire \ADC_IAC.n15014 ;
    wire AC_ADC_SYNC;
    wire n14_adj_1662_cascade_;
    wire IAC_CS;
    wire DDS_CS1;
    wire \RTD.cfg_tmp_1 ;
    wire \RTD.cfg_tmp_2 ;
    wire \RTD.cfg_tmp_3 ;
    wire \RTD.cfg_tmp_4 ;
    wire \RTD.cfg_tmp_5 ;
    wire \RTD.cfg_tmp_6 ;
    wire \RTD.adc_state_0 ;
    wire \RTD.cfg_tmp_7 ;
    wire adc_state_2;
    wire \RTD.cfg_tmp_0 ;
    wire \RTD.n13137 ;
    wire \RTD.n15115 ;
    wire \RTD.cfg_buf_5 ;
    wire \RTD.n11_adj_1444 ;
    wire \RTD.cfg_buf_3 ;
    wire \RTD.cfg_buf_4 ;
    wire \RTD.cfg_buf_2 ;
    wire \RTD.n10 ;
    wire \RTD.n11 ;
    wire \RTD.adc_state_3 ;
    wire \RTD.n21036 ;
    wire \RTD.n21199 ;
    wire \RTD.n13090_cascade_ ;
    wire \RTD.cfg_buf_1 ;
    wire \RTD.n12 ;
    wire \RTD.cfg_buf_7 ;
    wire \RTD.n13090 ;
    wire \RTD.n21061 ;
    wire \RTD.cfg_buf_0 ;
    wire buf_readRTD_9;
    wire buf_adcdata_vdc_3;
    wire buf_adcdata_iac_3;
    wire n19_adj_1609_cascade_;
    wire buf_readRTD_14;
    wire cmd_rdadctmp_10_adj_1482;
    wire DDS_MOSI1;
    wire n20_adj_1693;
    wire n22407;
    wire buf_adcdata_vac_2;
    wire n19_adj_1612_cascade_;
    wire buf_adcdata_vac_6;
    wire buf_adcdata_vac_22;
    wire n22629;
    wire cmd_rdadctmp_14_adj_1478;
    wire cmd_rdadctmp_15_adj_1477;
    wire buf_data_iac_6;
    wire n22_adj_1601;
    wire buf_data_iac_2;
    wire n22_adj_1613;
    wire buf_readRTD_10;
    wire buf_cfgRTD_2;
    wire cmd_rdadctmp_11_adj_1481;
    wire buf_adcdata_vac_3;
    wire cmd_rdadctmp_13_adj_1479;
    wire cmd_rdadctmp_30_adj_1462;
    wire buf_adcdata_vac_9;
    wire cmd_rdadctmp_11;
    wire cmd_rdadctmp_12;
    wire cmd_rdadctmp_8;
    wire cmd_rdadctmp_17_adj_1475;
    wire cmd_rdadctmp_29_adj_1463;
    wire cmd_rdadctmp_9_adj_1483;
    wire \CLK_DDS.tmp_buf_10 ;
    wire \CLK_DDS.tmp_buf_11 ;
    wire \CLK_DDS.tmp_buf_12 ;
    wire \CLK_DDS.tmp_buf_13 ;
    wire \CLK_DDS.tmp_buf_14 ;
    wire \CLK_DDS.tmp_buf_9 ;
    wire \CLK_DDS.tmp_buf_8 ;
    wire buf_readRTD_7;
    wire n16_adj_1690;
    wire n17_adj_1691;
    wire \ADC_IAC.n12 ;
    wire \ADC_IAC.n21457 ;
    wire cmd_rdadctmp_7;
    wire cmd_rdadctmp_6;
    wire n21082;
    wire n21082_cascade_;
    wire cmd_rdadctmp_3;
    wire n12771_cascade_;
    wire cmd_rdadctmp_4;
    wire cmd_rdadctmp_5;
    wire \ADC_IAC.n17 ;
    wire DDS_MCLK1;
    wire cmd_rdadctmp_0_adj_1523;
    wire \ADC_VDC.cmd_rdadcbuf_0 ;
    wire bfn_8_6_0_;
    wire \ADC_VDC.cmd_rdadcbuf_1 ;
    wire \ADC_VDC.n19842 ;
    wire \ADC_VDC.cmd_rdadcbuf_2 ;
    wire \ADC_VDC.n19843 ;
    wire \ADC_VDC.cmd_rdadcbuf_3 ;
    wire \ADC_VDC.n19844 ;
    wire \ADC_VDC.cmd_rdadcbuf_4 ;
    wire \ADC_VDC.n19845 ;
    wire \ADC_VDC.cmd_rdadcbuf_5 ;
    wire \ADC_VDC.n19846 ;
    wire cmd_rdadctmp_6_adj_1517;
    wire \ADC_VDC.cmd_rdadcbuf_6 ;
    wire \ADC_VDC.n19847 ;
    wire \ADC_VDC.cmd_rdadcbuf_7 ;
    wire \ADC_VDC.n19848 ;
    wire \ADC_VDC.n19849 ;
    wire \ADC_VDC.cmd_rdadcbuf_8 ;
    wire bfn_8_7_0_;
    wire \ADC_VDC.cmd_rdadcbuf_9 ;
    wire \ADC_VDC.n19850 ;
    wire \ADC_VDC.cmd_rdadcbuf_10 ;
    wire \ADC_VDC.n19851 ;
    wire \ADC_VDC.n19852 ;
    wire \ADC_VDC.n19853 ;
    wire \ADC_VDC.n19854 ;
    wire cmd_rdadcbuf_14;
    wire \ADC_VDC.n19855 ;
    wire \ADC_VDC.n19856 ;
    wire \ADC_VDC.n19857 ;
    wire cmd_rdadctmp_16_adj_1507;
    wire bfn_8_8_0_;
    wire cmd_rdadctmp_17_adj_1506;
    wire \ADC_VDC.n19858 ;
    wire cmd_rdadctmp_18_adj_1505;
    wire \ADC_VDC.n19859 ;
    wire \ADC_VDC.n19860 ;
    wire \ADC_VDC.n19861 ;
    wire \ADC_VDC.n19862 ;
    wire \ADC_VDC.n19863 ;
    wire \ADC_VDC.n19864 ;
    wire \ADC_VDC.n19865 ;
    wire bfn_8_9_0_;
    wire \ADC_VDC.n19866 ;
    wire \ADC_VDC.n19867 ;
    wire \ADC_VDC.n19868 ;
    wire \ADC_VDC.n19869 ;
    wire cmd_rdadcbuf_29;
    wire \ADC_VDC.n19870 ;
    wire \ADC_VDC.n19871 ;
    wire \ADC_VDC.n19872 ;
    wire \ADC_VDC.n19873 ;
    wire bfn_8_10_0_;
    wire \ADC_VDC.n19874 ;
    wire \ADC_VDC.n19875 ;
    wire buf_adcdata_vdc_18;
    wire buf_adcdata_vac_18;
    wire n19_adj_1692;
    wire cmd_rdadctmp_13;
    wire cmd_rdadctmp_10;
    wire buf_adcdata_iac_2;
    wire buf_adcdata_vac_5;
    wire buf_adcdata_iac_5;
    wire n19_adj_1603_cascade_;
    wire n22377_cascade_;
    wire n21237;
    wire cmd_rdadctmp_28_adj_1464;
    wire tmp_buf_15_adj_1497;
    wire \CLK_DDS.tmp_buf_0 ;
    wire \CLK_DDS.tmp_buf_1 ;
    wire \CLK_DDS.tmp_buf_2 ;
    wire \CLK_DDS.tmp_buf_3 ;
    wire \CLK_DDS.tmp_buf_4 ;
    wire \CLK_DDS.tmp_buf_5 ;
    wire \CLK_DDS.tmp_buf_6 ;
    wire \CLK_DDS.tmp_buf_7 ;
    wire buf_adcdata_vac_17;
    wire \SIG_DDS.bit_cnt_1 ;
    wire \SIG_DDS.bit_cnt_2 ;
    wire \SIG_DDS.n10 ;
    wire bit_cnt_0;
    wire cmd_rdadctmp_4_adj_1488;
    wire cmd_rdadctmp_5_adj_1487;
    wire cmd_rdadctmp_6_adj_1486;
    wire cmd_rdadctmp_22;
    wire n15092;
    wire IAC_DRDY;
    wire \ADC_IAC.n21159_cascade_ ;
    wire \ADC_IAC.n21160 ;
    wire cmd_rdadctmp_1;
    wire cmd_rdadctmp_2;
    wire IAC_MISO;
    wire cmd_rdadctmp_0;
    wire DTRIG_N_958;
    wire adc_state_1;
    wire IAC_SCLK;
    wire buf_adcdata_iac_17;
    wire cmd_rdadcbuf_27;
    wire \ADC_VDC.n10309_cascade_ ;
    wire \ADC_VDC.n13276 ;
    wire cmd_rdadctmp_1_adj_1522;
    wire cmd_rdadctmp_2_adj_1521;
    wire cmd_rdadctmp_3_adj_1520;
    wire cmd_rdadctmp_4_adj_1519;
    wire cmd_rdadctmp_5_adj_1518;
    wire cmd_rdadctmp_7_adj_1516;
    wire cmd_rdadctmp_19_adj_1504;
    wire cmd_rdadctmp_8_adj_1515;
    wire cmd_rdadctmp_9_adj_1514;
    wire cmd_rdadctmp_10_adj_1513;
    wire cmd_rdadctmp_11_adj_1512;
    wire cmd_rdadctmp_12_adj_1511;
    wire cmd_rdadctmp_13_adj_1510;
    wire cmd_rdadctmp_14_adj_1509;
    wire cmd_rdadctmp_15_adj_1508;
    wire cmd_rdadcbuf_20;
    wire buf_adcdata_vdc_9;
    wire cmd_rdadcbuf_17;
    wire buf_adcdata_vdc_6;
    wire cmd_rdadcbuf_11;
    wire buf_dds1_5;
    wire cmd_rdadcbuf_21;
    wire cmd_rdadcbuf_33;
    wire buf_adcdata_vdc_22;
    wire cmd_rdadcbuf_13;
    wire buf_adcdata_vdc_2;
    wire cmd_rdadcbuf_15;
    wire buf_adcdata_vdc_4;
    wire cmd_rdadcbuf_16;
    wire buf_adcdata_vdc_5;
    wire cmd_rdadctmp_20_adj_1503;
    wire cmd_rdadctmp_21_adj_1502;
    wire \ADC_VDC.cmd_rdadcbuf_35_N_1296_34 ;
    wire \ADC_VDC.n19 ;
    wire \ADC_VDC.n21_cascade_ ;
    wire cmd_rdadcbuf_34;
    wire \ADC_VDC.n18780_cascade_ ;
    wire \ADC_VDC.n4_adj_1451 ;
    wire \ADC_VDC.n13503 ;
    wire buf_readRTD_8;
    wire buf_adcdata_vdc_16;
    wire buf_adcdata_vac_16;
    wire n22575_cascade_;
    wire buf_cfgRTD_0;
    wire n10902_cascade_;
    wire n12624_cascade_;
    wire buf_cfgRTD_3;
    wire buf_readRTD_11;
    wire n22473;
    wire bfn_9_11_0_;
    wire n19813;
    wire n19814;
    wire n19815;
    wire n19816;
    wire n19817;
    wire n19818;
    wire n19819;
    wire n19820;
    wire bfn_9_12_0_;
    wire n19821;
    wire n19822;
    wire n19823;
    wire n19824;
    wire n19825;
    wire n19826;
    wire n19827;
    wire cmd_rdadctmp_27_adj_1465;
    wire buf_adcdata_vac_19;
    wire n12493;
    wire n21705;
    wire cmd_rdadctmp_18_adj_1474;
    wire IAC_OSR1;
    wire data_idxvec_11;
    wire n26_adj_1678_cascade_;
    wire n22509;
    wire buf_dds1_2;
    wire n22476;
    wire cmd_rdadctmp_16_adj_1476;
    wire cmd_rdadctmp_25_adj_1467;
    wire cmd_rdadctmp_24_adj_1468;
    wire cmd_rdadctmp_22_adj_1470;
    wire cmd_rdadctmp_23_adj_1469;
    wire n69;
    wire cmd_rdadctmp_15;
    wire IAC_FLT1;
    wire buf_adcdata_iac_19;
    wire n22605_cascade_;
    wire buf_dds1_11;
    wire n22608;
    wire cmd_rdadctmp_27;
    wire cmd_rdadctmp_19;
    wire cmd_rdadctmp_24;
    wire cmd_rdadctmp_30;
    wire \ADC_VDC.n18780 ;
    wire \ADC_VDC.n18783_cascade_ ;
    wire \ADC_VDC.n16_adj_1450 ;
    wire \ADC_VDC.n18 ;
    wire \ADC_VDC.n18_cascade_ ;
    wire THERMOSTAT;
    wire \ADC_VDC.avg_cnt_0 ;
    wire bfn_10_6_0_;
    wire \ADC_VDC.avg_cnt_1 ;
    wire \ADC_VDC.n19877 ;
    wire \ADC_VDC.avg_cnt_2 ;
    wire \ADC_VDC.n19878 ;
    wire \ADC_VDC.n19879 ;
    wire \ADC_VDC.avg_cnt_4 ;
    wire \ADC_VDC.n19880 ;
    wire \ADC_VDC.avg_cnt_5 ;
    wire \ADC_VDC.n19881 ;
    wire \ADC_VDC.n19882 ;
    wire \ADC_VDC.avg_cnt_7 ;
    wire \ADC_VDC.n19883 ;
    wire \ADC_VDC.n19884 ;
    wire bfn_10_7_0_;
    wire \ADC_VDC.n19885 ;
    wire \ADC_VDC.avg_cnt_10 ;
    wire \ADC_VDC.n19886 ;
    wire \ADC_VDC.n19887 ;
    wire \ADC_VDC.avg_cnt_11 ;
    wire \ADC_VDC.n13463 ;
    wire \ADC_VDC.n15175 ;
    wire cmd_rdadcbuf_23;
    wire cmd_rdadcbuf_18;
    wire buf_adcdata_vdc_7;
    wire n11891_cascade_;
    wire cmd_rdadcbuf_26;
    wire cmd_rdadcbuf_25;
    wire cmd_rdadcbuf_22;
    wire buf_control_7;
    wire DDS_SCK1;
    wire buf_readRTD_15;
    wire buf_adcdata_vdc_23;
    wire n22593_cascade_;
    wire buf_adcdata_vac_23;
    wire buf_cfgRTD_6;
    wire buf_cfgRTD_7;
    wire n30_adj_1499;
    wire cmd_rdadctmp_19_adj_1473;
    wire buf_adcdata_vac_21;
    wire VAC_OSR1;
    wire buf_adcdata_vdc_10;
    wire buf_adcdata_vac_10;
    wire buf_adcdata_vdc_0;
    wire buf_adcdata_vac_0;
    wire buf_adcdata_iac_0;
    wire n19_adj_1534_cascade_;
    wire n19_adj_1652;
    wire buf_readRTD_1;
    wire buf_adcdata_vac_13;
    wire buf_readRTD_5;
    wire n19_adj_1629_cascade_;
    wire n12850;
    wire cmd_rdadctmp_21_adj_1471;
    wire n8;
    wire n10695;
    wire buf_adcdata_vdc_12;
    wire n21076;
    wire adc_state_0_adj_1460;
    wire cmd_rdadctmp_20_adj_1472;
    wire buf_adcdata_vac_12;
    wire iac_raw_buf_N_774;
    wire n21334;
    wire n22512;
    wire data_idxvec_15;
    wire buf_data_iac_23;
    wire n26_adj_1659_cascade_;
    wire n21324_cascade_;
    wire buf_adcdata_vac_15;
    wire buf_adcdata_vdc_15;
    wire n19_adj_1621;
    wire n23_adj_1658;
    wire n21323;
    wire n22371;
    wire n12_adj_1454_cascade_;
    wire acadc_trig;
    wire n21053;
    wire n21042_cascade_;
    wire n21030_cascade_;
    wire eis_end;
    wire INVacadc_trig_300C_net;
    wire n17728;
    wire n11_cascade_;
    wire acadc_dtrig_v;
    wire acadc_dtrig_i;
    wire eis_state_2_N_392_1;
    wire eis_state_2_N_392_1_cascade_;
    wire n2_adj_1696_cascade_;
    wire n22437;
    wire INVeis_state_i1C_net;
    wire cmd_rdadctmp_23;
    wire VAC_FLT1;
    wire cmd_rdadctmp_29;
    wire buf_adcdata_iac_21;
    wire cmd_rdadctmp_28;
    wire cmd_rdadctmp_25;
    wire cmd_rdadctmp_20;
    wire n12771;
    wire cmd_rdadctmp_31;
    wire buf_adcdata_iac_23;
    wire \ADC_VDC.n16 ;
    wire \ADC_VDC.n21593_cascade_ ;
    wire \ADC_VDC.n21590_cascade_ ;
    wire \ADC_VDC.n22590 ;
    wire n13324;
    wire \ADC_VDC.n7_cascade_ ;
    wire \ADC_VDC.n21193 ;
    wire cmd_rdadcbuf_19;
    wire cmd_rdadcbuf_24;
    wire buf_adcdata_vdc_13;
    wire cmd_rdadcbuf_30;
    wire buf_adcdata_vdc_19;
    wire cmd_rdadcbuf_28;
    wire buf_adcdata_vdc_17;
    wire cmd_rdadcbuf_32;
    wire buf_adcdata_vdc_21;
    wire cmd_rdadcbuf_31;
    wire buf_dds1_4;
    wire \ADC_VDC.n22587 ;
    wire \ADC_VDC.n10708 ;
    wire cmd_rdadctmp_22_adj_1501;
    wire \ADC_VDC.n10708_cascade_ ;
    wire \ADC_VDC.cmd_rdadctmp_23 ;
    wire \ADC_VDC.n5 ;
    wire \ADC_VDC.avg_cnt_9 ;
    wire \ADC_VDC.avg_cnt_8 ;
    wire \ADC_VDC.avg_cnt_6 ;
    wire \ADC_VDC.avg_cnt_3 ;
    wire \ADC_VDC.n20 ;
    wire \CLK_DDS.n13005 ;
    wire \CLK_DDS.n9_adj_1433 ;
    wire dds_state_2_adj_1494;
    wire dds_state_0_adj_1496;
    wire dds_state_1_adj_1495;
    wire \CLK_DDS.n9 ;
    wire bfn_11_7_0_;
    wire n19956;
    wire n19957;
    wire n19958;
    wire n19959;
    wire n19960;
    wire n19961;
    wire n19962;
    wire n19963;
    wire bfn_11_8_0_;
    wire n19964;
    wire n19965;
    wire n19966;
    wire n19967;
    wire n19968;
    wire n19969;
    wire n19970;
    wire n19971;
    wire bfn_11_9_0_;
    wire n19972;
    wire n19973;
    wire n19974;
    wire n19975;
    wire n19976;
    wire n19977;
    wire secclk_cnt_21;
    wire secclk_cnt_19;
    wire secclk_cnt_12;
    wire secclk_cnt_22;
    wire n14_adj_1571;
    wire n21329;
    wire IAC_FLT0;
    wire n22374;
    wire n21240;
    wire n22401;
    wire n21122;
    wire n21122_cascade_;
    wire n12610_cascade_;
    wire buf_data_iac_5;
    wire n22_adj_1604;
    wire data_idxvec_4;
    wire n26_adj_1635_cascade_;
    wire n22443_cascade_;
    wire n22446_cascade_;
    wire n30_adj_1636_cascade_;
    wire n19_adj_1634;
    wire buf_readRTD_4;
    wire buf_adcdata_iac_12;
    wire n22467_cascade_;
    wire n16_adj_1633;
    wire n22470;
    wire n22395_cascade_;
    wire req_data_cnt_8;
    wire VAC_FLT0;
    wire buf_adcdata_iac_22;
    wire n22635_cascade_;
    wire n21236;
    wire n14_adj_1578;
    wire n2_cascade_;
    wire n21501_cascade_;
    wire eis_state_2_N_392_0;
    wire n22479;
    wire eis_start;
    wire n11_adj_1632_cascade_;
    wire INVeis_state_i0C_net;
    wire n11908;
    wire eis_state_0;
    wire n21041;
    wire buf_dds1_15;
    wire buf_dds1_10;
    wire acadc_skipCount_15;
    wire n11570;
    wire EIS_SYNCCLK;
    wire IAC_CLK;
    wire buf_dds0_10;
    wire \SIG_DDS.tmp_buf_10 ;
    wire buf_dds0_11;
    wire \SIG_DDS.tmp_buf_11 ;
    wire \SIG_DDS.tmp_buf_12 ;
    wire \SIG_DDS.tmp_buf_13 ;
    wire buf_dds0_14;
    wire buf_dds0_15;
    wire \SIG_DDS.tmp_buf_14 ;
    wire buf_dds0_9;
    wire \SIG_DDS.tmp_buf_9 ;
    wire \SIG_DDS.tmp_buf_8 ;
    wire \SIG_DDS.tmp_buf_0 ;
    wire buf_dds0_1;
    wire \SIG_DDS.tmp_buf_1 ;
    wire buf_dds0_2;
    wire \SIG_DDS.tmp_buf_2 ;
    wire \SIG_DDS.tmp_buf_3 ;
    wire \SIG_DDS.tmp_buf_4 ;
    wire \SIG_DDS.tmp_buf_5 ;
    wire \ADC_VDC.n21007 ;
    wire \ADC_VDC.n21007_cascade_ ;
    wire \ADC_VDC.n4 ;
    wire \ADC_VDC.n11 ;
    wire \ADC_VDC.n65 ;
    wire \ADC_VDC.n21133 ;
    wire \ADC_VDC.n42_adj_1452 ;
    wire \ADC_VDC.n20998 ;
    wire \ADC_VDC.n11494 ;
    wire \ADC_VDC.n11494_cascade_ ;
    wire \ADC_VDC.n15 ;
    wire \ADC_VDC.n15_cascade_ ;
    wire \ADC_VDC.n21185 ;
    wire n11891;
    wire cmd_rdadcbuf_12;
    wire \ADC_VDC.n21203 ;
    wire \ADC_VDC.n21211 ;
    wire \ADC_VDC.n13368 ;
    wire secclk_cnt_20;
    wire n20048_cascade_;
    wire n14;
    wire buf_adcdata_vdc_20;
    wire buf_adcdata_vac_20;
    wire secclk_cnt_6;
    wire secclk_cnt_14;
    wire secclk_cnt_10;
    wire secclk_cnt_3;
    wire n27;
    wire secclk_cnt_2;
    wire secclk_cnt_13;
    wire secclk_cnt_7;
    wire secclk_cnt_16;
    wire n26_adj_1656;
    wire n14_adj_1552;
    wire n30;
    wire n14_adj_1574;
    wire buf_data_iac_3;
    wire n22_adj_1610;
    wire req_data_cnt_14;
    wire req_data_cnt_11;
    wire n23;
    wire n14_adj_1551;
    wire buf_dds0_4;
    wire n23_adj_1661;
    wire acadc_skipCount_14;
    wire buf_adcdata_vdc_1;
    wire buf_adcdata_vac_1;
    wire buf_adcdata_iac_20;
    wire VAC_OSR0;
    wire comm_cmd_4;
    wire n16818_cascade_;
    wire n16_adj_1628;
    wire n22365;
    wire data_idxvec_5;
    wire n26_adj_1630_cascade_;
    wire n22449_cascade_;
    wire req_data_cnt_5;
    wire n22368;
    wire n22452_cascade_;
    wire n30_adj_1631_cascade_;
    wire n9;
    wire buf_data_iac_22;
    wire data_idxvec_14;
    wire n21330;
    wire acadc_skipCount_11;
    wire n23_adj_1677;
    wire buf_dds1_9;
    wire buf_adcdata_vdc_14;
    wire buf_adcdata_vac_14;
    wire n20;
    wire n17_cascade_;
    wire n19_adj_1526;
    wire n29;
    wire data_idxvec_13;
    wire buf_dds1_3;
    wire acadc_skipCount_4;
    wire n8_adj_1560;
    wire n8_adj_1560_cascade_;
    wire data_index_9_N_212_7;
    wire n24_adj_1593;
    wire n23_adj_1591;
    wire n22_adj_1590_cascade_;
    wire n18;
    wire n30_adj_1543_cascade_;
    wire n31_adj_1537;
    wire cmd_rdadctmp_26;
    wire buf_adcdata_iac_18;
    wire acadc_skipCount_8;
    wire n14_adj_1538_cascade_;
    wire n26_adj_1525;
    wire cmd_rdadctmp_21;
    wire buf_adcdata_iac_13;
    wire acadc_skipCount_13;
    wire buf_dds0_5;
    wire buf_dds0_3;
    wire acadc_skipCount_5;
    wire n20_adj_1670;
    wire cmd_rdadctmp_16;
    wire cmd_rdadctmp_17;
    wire data_count_0;
    wire bfn_12_18_0_;
    wire data_count_1;
    wire n19765;
    wire data_count_2;
    wire n19766;
    wire data_count_3;
    wire n19767;
    wire data_count_4;
    wire n19768;
    wire data_count_5;
    wire n19769;
    wire data_count_6;
    wire n19770;
    wire data_count_7;
    wire n19771;
    wire n19772;
    wire INVdata_count_i0_i0C_net;
    wire data_count_8;
    wire bfn_12_19_0_;
    wire n19773;
    wire data_count_9;
    wire INVdata_count_i0_i8C_net;
    wire \comm_spi.n23089 ;
    wire \comm_spi.n14822 ;
    wire \comm_spi.n23089_cascade_ ;
    wire \comm_spi.n14823 ;
    wire \ADC_VDC.bit_cnt_0 ;
    wire bfn_13_6_0_;
    wire \ADC_VDC.bit_cnt_1 ;
    wire \ADC_VDC.n19918 ;
    wire \ADC_VDC.bit_cnt_2 ;
    wire \ADC_VDC.n19919 ;
    wire \ADC_VDC.bit_cnt_3 ;
    wire \ADC_VDC.n19920 ;
    wire \ADC_VDC.bit_cnt_4 ;
    wire \ADC_VDC.n19921 ;
    wire \ADC_VDC.bit_cnt_5 ;
    wire \ADC_VDC.n19922 ;
    wire \ADC_VDC.bit_cnt_6 ;
    wire \ADC_VDC.n19923 ;
    wire \ADC_VDC.n19924 ;
    wire \ADC_VDC.bit_cnt_7 ;
    wire \ADC_VDC.n15273 ;
    wire n21_adj_1594;
    wire n14899;
    wire TEST_LED;
    wire secclk_cnt_15;
    wire secclk_cnt_8;
    wire secclk_cnt_1;
    wire secclk_cnt_5;
    wire n25;
    wire secclk_cnt_18;
    wire secclk_cnt_0;
    wire secclk_cnt_11;
    wire secclk_cnt_4;
    wire n28_adj_1554;
    wire req_data_cnt_15;
    wire n24;
    wire req_data_cnt_12;
    wire n22;
    wire n14_adj_1548;
    wire \comm_spi.n23095 ;
    wire \comm_spi.data_tx_7__N_807 ;
    wire req_data_cnt_13;
    wire secclk_cnt_9;
    wire secclk_cnt_17;
    wire n10;
    wire n19_adj_1683;
    wire n20_adj_1684;
    wire buf_adcdata_vdc_11;
    wire buf_adcdata_vac_11;
    wire buf_readRTD_12;
    wire buf_cfgRTD_4;
    wire buf_dds1_13;
    wire buf_cfgRTD_5;
    wire buf_readRTD_13;
    wire n9269;
    wire n12082_cascade_;
    wire n14_adj_1573;
    wire \comm_spi.data_tx_7__N_817 ;
    wire req_data_cnt_10;
    wire n19_adj_1646;
    wire buf_readRTD_2;
    wire n16_adj_1645;
    wire n22641_cascade_;
    wire data_idxvec_2;
    wire n26_adj_1647_cascade_;
    wire acadc_skipCount_2;
    wire n22383_cascade_;
    wire req_data_cnt_2;
    wire n22644;
    wire n22386_cascade_;
    wire n30_adj_1648_cascade_;
    wire req_data_cnt_4;
    wire n18_adj_1644;
    wire buf_dds0_13;
    wire n66;
    wire buf_dds1_14;
    wire buf_dds1_1;
    wire n12662;
    wire n5_adj_1536;
    wire n7_adj_1650_cascade_;
    wire n12;
    wire SELIRNG1;
    wire n14_adj_1546;
    wire n14_adj_1549;
    wire n8_adj_1562;
    wire data_index_9_N_212_6;
    wire n17_adj_1553;
    wire AMPV_POW;
    wire data_index_9_N_212_3;
    wire eis_state_1;
    wire eis_state_2;
    wire acadc_rst;
    wire n20011;
    wire n19_adj_1616;
    wire n14_adj_1547;
    wire n8_adj_1564_cascade_;
    wire data_index_9_N_212_4;
    wire cmd_rdadctmp_9;
    wire buf_adcdata_iac_1;
    wire buf_dds1_12;
    wire buf_dds0_12;
    wire n8_adj_1566;
    wire n8_adj_1566_cascade_;
    wire \SIG_DDS.tmp_buf_6 ;
    wire \SIG_DDS.tmp_buf_7 ;
    wire \SIG_DDS.bit_cnt_3 ;
    wire \SIG_DDS.n21744 ;
    wire buf_dds1_7;
    wire acadc_skipcnt_0;
    wire bfn_13_18_0_;
    wire INVacadc_skipcnt_i0_i0C_net;
    wire n21226;
    wire n19789;
    wire n19789_THRU_CRY_0_THRU_CO;
    wire n19789_THRU_CRY_1_THRU_CO;
    wire n19789_THRU_CRY_2_THRU_CO;
    wire n19789_THRU_CRY_3_THRU_CO;
    wire n19789_THRU_CRY_4_THRU_CO;
    wire GNDG0;
    wire n19789_THRU_CRY_5_THRU_CO;
    wire n19789_THRU_CRY_6_THRU_CO;
    wire acadc_skipcnt_1;
    wire bfn_13_19_0_;
    wire acadc_skipcnt_2;
    wire n19790;
    wire acadc_skipcnt_3;
    wire n19791;
    wire acadc_skipcnt_4;
    wire n19792;
    wire acadc_skipcnt_5;
    wire n19793;
    wire acadc_skipcnt_6;
    wire n19794;
    wire acadc_skipcnt_7;
    wire n19795;
    wire acadc_skipcnt_8;
    wire n19796;
    wire n19797;
    wire INVacadc_skipcnt_i0_i1C_net;
    wire acadc_skipcnt_9;
    wire bfn_13_20_0_;
    wire n19798;
    wire acadc_skipcnt_11;
    wire n19799;
    wire n19800;
    wire acadc_skipcnt_13;
    wire n19801;
    wire acadc_skipcnt_14;
    wire n19802;
    wire n19803;
    wire acadc_skipcnt_15;
    wire INVacadc_skipcnt_i0_i9C_net;
    wire n11989;
    wire n14915;
    wire \INVcomm_spi.imiso_83_12297_12298_resetC_net ;
    wire \comm_spi.n23083 ;
    wire \comm_spi.n14846 ;
    wire \comm_spi.n14847 ;
    wire \INVADC_VDC.genclk.t_clk_24C_net ;
    wire \comm_spi.n14808 ;
    wire \comm_spi.n14809 ;
    wire \comm_spi.imosi_cascade_ ;
    wire \comm_spi.DOUT_7__N_786 ;
    wire \comm_spi.imosi_N_792 ;
    wire n12_adj_1542_cascade_;
    wire n19986_cascade_;
    wire n30_adj_1530;
    wire n33;
    wire n34_cascade_;
    wire n31;
    wire n49_cascade_;
    wire n32;
    wire \INVcomm_spi.bit_cnt_3767__i3C_net ;
    wire n19_adj_1673;
    wire n20_adj_1674;
    wire \comm_spi.bit_cnt_1 ;
    wire \comm_spi.bit_cnt_2 ;
    wire \comm_spi.bit_cnt_0 ;
    wire n14_adj_1579;
    wire n14_adj_1572;
    wire n4_adj_1637;
    wire n14_adj_1544;
    wire n14_adj_1575;
    wire n19_adj_1666;
    wire n20_adj_1667;
    wire n16_adj_1664;
    wire n17_adj_1665;
    wire n22413_cascade_;
    wire n21671;
    wire n23_adj_1668;
    wire n22569_cascade_;
    wire n21702;
    wire n22416;
    wire n22572_cascade_;
    wire n30_adj_1669_cascade_;
    wire n22404;
    wire n22380;
    wire n30_adj_1679;
    wire n8_adj_1689_cascade_;
    wire n26_adj_1595_cascade_;
    wire n18_adj_1615;
    wire n16818;
    wire n21714;
    wire n7_cascade_;
    wire n12107;
    wire iac_raw_buf_N_776;
    wire bfn_14_13_0_;
    wire n19774;
    wire data_cntvec_2;
    wire n19775;
    wire n19776;
    wire data_cntvec_4;
    wire n19777;
    wire data_cntvec_5;
    wire n19778;
    wire n19779;
    wire n19780;
    wire n19781;
    wire INVdata_cntvec_i0_i0C_net;
    wire bfn_14_14_0_;
    wire n19782;
    wire n19783;
    wire data_cntvec_11;
    wire n19784;
    wire data_cntvec_12;
    wire n19785;
    wire data_cntvec_13;
    wire n19786;
    wire data_cntvec_14;
    wire n19787;
    wire n19788;
    wire data_cntvec_15;
    wire INVdata_cntvec_i0_i8C_net;
    wire n11933;
    wire n14907;
    wire bfn_14_15_0_;
    wire n19804;
    wire n19805;
    wire data_index_3;
    wire n7_adj_1565;
    wire n19806;
    wire n19807;
    wire n19808;
    wire data_index_6;
    wire n7_adj_1561;
    wire n19809;
    wire data_index_7;
    wire n7_adj_1559;
    wire n19810;
    wire n19811;
    wire bfn_14_16_0_;
    wire n10756;
    wire n19812;
    wire buf_data_iac_1;
    wire n22_adj_1617;
    wire trig_dds1;
    wire buf_dds0_7;
    wire n21079;
    wire adc_state_0;
    wire cmd_rdadctmp_18;
    wire buf_adcdata_iac_10;
    wire n8_adj_1564;
    wire n7_adj_1563;
    wire data_index_4;
    wire n11611;
    wire buf_adcdata_iac_16;
    wire buf_dds1_8;
    wire n22389_cascade_;
    wire buf_dds0_8;
    wire data_index_5;
    wire DDS_SCK;
    wire tmp_buf_15;
    wire DDS_MOSI;
    wire data_index_9;
    wire n12624;
    wire buf_cfgRTD_1;
    wire n12610;
    wire IAC_OSR0;
    wire data_index_9_N_212_8;
    wire data_index_1;
    wire n8_adj_1570;
    wire n8_adj_1570_cascade_;
    wire n7_adj_1569;
    wire data_index_9_N_212_1;
    wire data_index_2;
    wire n8_adj_1558;
    wire n7_adj_1557;
    wire data_index_8;
    wire n8_adj_1568;
    wire n7_adj_1567;
    wire data_index_9_N_212_2;
    wire \comm_spi.n14815 ;
    wire \comm_spi.n14816 ;
    wire \INVcomm_spi.imiso_83_12297_12298_setC_net ;
    wire \comm_spi.imosi ;
    wire \comm_spi.DOUT_7__N_787 ;
    wire wdtick_cnt_0;
    wire bfn_15_5_0_;
    wire wdtick_cnt_1;
    wire n19932;
    wire wdtick_cnt_2;
    wire n19933;
    wire wdtick_cnt_3;
    wire n19934;
    wire wdtick_cnt_4;
    wire n19935;
    wire wdtick_cnt_5;
    wire n19936;
    wire wdtick_cnt_6;
    wire n19937;
    wire wdtick_cnt_7;
    wire n19938;
    wire n19939;
    wire wdtick_cnt_8;
    wire bfn_15_6_0_;
    wire wdtick_cnt_9;
    wire n19940;
    wire wdtick_cnt_10;
    wire n19941;
    wire wdtick_cnt_11;
    wire n19942;
    wire wdtick_cnt_12;
    wire n19943;
    wire wdtick_cnt_13;
    wire n19944;
    wire wdtick_cnt_14;
    wire n19945;
    wire wdtick_cnt_15;
    wire n19946;
    wire n19947;
    wire wdtick_cnt_16;
    wire bfn_15_7_0_;
    wire wdtick_cnt_17;
    wire n19948;
    wire wdtick_cnt_18;
    wire n19949;
    wire wdtick_cnt_19;
    wire n19950;
    wire wdtick_cnt_20;
    wire n19951;
    wire wdtick_cnt_21;
    wire n19952;
    wire wdtick_cnt_22;
    wire n19953;
    wire wdtick_cnt_23;
    wire n19954;
    wire n19955;
    wire n49;
    wire bfn_15_8_0_;
    wire wdtick_cnt_24;
    wire clk_RTD;
    wire n14_adj_1550;
    wire n17_adj_1672;
    wire n22461;
    wire n16_adj_1671;
    wire data_idxvec_12;
    wire n21556_cascade_;
    wire n21703;
    wire n22521;
    wire n22464;
    wire n22524_cascade_;
    wire n30_adj_1676_cascade_;
    wire n17_adj_1682;
    wire n16_adj_1681;
    wire n22485;
    wire data_idxvec_10;
    wire data_cntvec_10;
    wire n26_adj_1687_cascade_;
    wire n22455_cascade_;
    wire n24_adj_1686;
    wire n22488;
    wire n22458_cascade_;
    wire n30_adj_1688_cascade_;
    wire data_idxvec_8;
    wire data_cntvec_8;
    wire buf_data_iac_16;
    wire n26_adj_1533_cascade_;
    wire n22398;
    wire n21246_cascade_;
    wire n22392;
    wire n22578;
    wire n22581_cascade_;
    wire n22584_cascade_;
    wire buf_readRTD_3;
    wire n19_adj_1641;
    wire buf_adcdata_iac_11;
    wire n16_adj_1640;
    wire n22623_cascade_;
    wire n22626_cascade_;
    wire n30_adj_1643;
    wire data_idxvec_3;
    wire data_cntvec_3;
    wire n26_adj_1642_cascade_;
    wire req_data_cnt_3;
    wire n22425_cascade_;
    wire acadc_skipCount_3;
    wire n22428;
    wire data_index_0;
    wire n8841;
    wire n8_adj_1540;
    wire n7_adj_1539;
    wire n8_adj_1540_cascade_;
    wire data_index_9_N_212_0;
    wire buf_dds1_0;
    wire n16_cascade_;
    wire buf_adcdata_iac_8;
    wire n12596;
    wire buf_dds0_0;
    wire VDC_RNG0;
    wire n23_adj_1675;
    wire buf_dds0_6;
    wire n17705;
    wire n9342_cascade_;
    wire n17703;
    wire data_index_9_N_212_5;
    wire buf_adcdata_iac_15;
    wire n16_adj_1620;
    wire n12144;
    wire DDS_CS;
    wire \SIG_DDS.n9_adj_1434 ;
    wire n8_adj_1556;
    wire n7_adj_1555;
    wire data_index_9_N_212_9;
    wire \INVcomm_spi.MISO_48_12291_12292_resetC_net ;
    wire \comm_spi.n14818 ;
    wire \comm_spi.n14819 ;
    wire \INVcomm_spi.MISO_48_12291_12292_setC_net ;
    wire buf_data_iac_21;
    wire n21672;
    wire \ADC_VDC.n22124_cascade_ ;
    wire VDC_SCLK;
    wire VDC_CLK;
    wire buf_data_iac_20;
    wire n21557;
    wire flagcntwd;
    wire n21187_cascade_;
    wire n11605;
    wire n20578;
    wire n11576_cascade_;
    wire n12148;
    wire n11910;
    wire buf_data_iac_10;
    wire n21385;
    wire comm_buf_0_7;
    wire n21276;
    wire n22542_cascade_;
    wire n4_adj_1580;
    wire \comm_spi.data_tx_7__N_814 ;
    wire comm_tx_buf_7;
    wire \comm_spi.data_tx_7__N_806 ;
    wire \comm_spi.bit_cnt_3 ;
    wire \comm_spi.n17254 ;
    wire \INVcomm_spi.data_valid_85C_net ;
    wire n22551_cascade_;
    wire comm_buf_1_4;
    wire n4_adj_1582_cascade_;
    wire n21285_cascade_;
    wire n22554;
    wire n21474_cascade_;
    wire n12_adj_1596_cascade_;
    wire data_idxvec_9;
    wire data_cntvec_9;
    wire buf_data_iac_17;
    wire n26_adj_1694_cascade_;
    wire eis_stop;
    wire req_data_cnt_9;
    wire acadc_skipCount_9;
    wire DDS_RNG_0;
    wire n22617_cascade_;
    wire n22620_cascade_;
    wire n21360;
    wire n22410;
    wire n21361_cascade_;
    wire n30_adj_1695_cascade_;
    wire n12184;
    wire n14958;
    wire n22539;
    wire n14_adj_1541;
    wire buf_data_iac_0;
    wire n22_adj_1532;
    wire n21586;
    wire comm_buf_6_7;
    wire acadc_skipCount_6;
    wire req_data_cnt_6;
    wire n19_adj_1625;
    wire buf_readRTD_6;
    wire data_idxvec_6;
    wire data_cntvec_6;
    wire n26_adj_1626_cascade_;
    wire n22515;
    wire n16_adj_1624;
    wire buf_adcdata_iac_14;
    wire n22527;
    wire n22530_cascade_;
    wire n22518;
    wire n30_adj_1627_cascade_;
    wire data_idxvec_0;
    wire data_cntvec_0;
    wire buf_data_iac_8;
    wire n26_cascade_;
    wire n21261_cascade_;
    wire n22563_cascade_;
    wire n21257;
    wire n22566_cascade_;
    wire buf_adcdata_vdc_8;
    wire buf_adcdata_vac_8;
    wire buf_readRTD_0;
    wire n19_cascade_;
    wire n21258;
    wire acadc_skipCount_0;
    wire req_data_cnt_0;
    wire n21260;
    wire buf_adcdata_iac_9;
    wire n16_adj_1651;
    wire n22431;
    wire data_idxvec_1;
    wire data_cntvec_1;
    wire n26_adj_1653_cascade_;
    wire acadc_skipCount_1;
    wire n22497_cascade_;
    wire req_data_cnt_1;
    wire n22434;
    wire n22500_cascade_;
    wire n30_adj_1654_cascade_;
    wire n28;
    wire comm_buf_1_7;
    wire n14965;
    wire trig_dds0;
    wire \SIG_DDS.n12895 ;
    wire wdtick_flag;
    wire buf_control_0;
    wire CONT_SD;
    wire dds_state_0;
    wire dds_state_2;
    wire \SIG_DDS.n9 ;
    wire dds_state_1;
    wire \comm_spi.n14813 ;
    wire \comm_spi.n14812 ;
    wire \comm_spi.n14811 ;
    wire ICE_SPI_MISO;
    wire \ADC_VDC.n11895 ;
    wire \comm_spi.n23086 ;
    wire \comm_spi.n23086_cascade_ ;
    wire \comm_spi.n14804 ;
    wire n80;
    wire n5;
    wire \comm_spi.n23092 ;
    wire clk_cnt_1;
    wire clk_cnt_0;
    wire n17773;
    wire buf_data_vac_8;
    wire buf_data_vac_15;
    wire comm_buf_4_7;
    wire buf_data_vac_14;
    wire buf_data_vac_13;
    wire buf_data_vac_12;
    wire comm_buf_4_4;
    wire buf_data_vac_11;
    wire buf_data_vac_10;
    wire buf_data_vac_9;
    wire n14986;
    wire n21268_cascade_;
    wire n22094;
    wire n21266;
    wire n12407;
    wire n21085_cascade_;
    wire n19188;
    wire n19188_cascade_;
    wire comm_buf_0_3;
    wire n22557_cascade_;
    wire comm_buf_1_3;
    wire comm_buf_4_3;
    wire n4_adj_1583_cascade_;
    wire n22560;
    wire n21288_cascade_;
    wire n21479;
    wire n21477_cascade_;
    wire n44_cascade_;
    wire n12260;
    wire comm_buf_1_2;
    wire n1_cascade_;
    wire n2_adj_1584;
    wire comm_buf_4_2;
    wire n21528;
    wire n4_adj_1585_cascade_;
    wire n22491;
    wire n21143;
    wire n19193_cascade_;
    wire n21273;
    wire comm_buf_1_0;
    wire n22533_cascade_;
    wire comm_buf_0_0;
    wire n22536;
    wire n24_adj_1639;
    wire n21497_cascade_;
    wire n34_adj_1649_cascade_;
    wire n30_adj_1531;
    wire comm_buf_2_0;
    wire n30_adj_1599;
    wire comm_buf_2_7;
    wire n30_adj_1602;
    wire n30_adj_1605;
    wire n30_adj_1608;
    wire comm_buf_2_4;
    wire n30_adj_1611;
    wire comm_buf_2_3;
    wire n30_adj_1614;
    wire comm_buf_2_2;
    wire n30_adj_1618;
    wire n12314;
    wire n14972;
    wire comm_buf_0_2;
    wire buf_data_iac_19;
    wire n21543;
    wire SELIRNG0;
    wire n23_adj_1685;
    wire comm_buf_6_0;
    wire comm_buf_6_3;
    wire acadc_skipCount_7;
    wire req_data_cnt_7;
    wire data_idxvec_7;
    wire data_cntvec_7;
    wire buf_data_iac_15;
    wire n26_adj_1622_cascade_;
    wire comm_cmd_1;
    wire n16824;
    wire comm_length_1;
    wire n5_adj_1524;
    wire n12654;
    wire comm_buf_0_4;
    wire comm_cmd_2;
    wire n21368;
    wire n21369;
    wire n21362;
    wire n21363;
    wire n22599_cascade_;
    wire comm_cmd_3;
    wire n22602;
    wire buf_dds1_6;
    wire n68;
    wire n12048;
    wire n12048_cascade_;
    wire n16971;
    wire \comm_spi.n14805 ;
    wire \comm_spi.iclk_N_802 ;
    wire ICE_SPI_SCLK;
    wire \comm_spi.iclk_N_803 ;
    wire buf_data_vac_0;
    wire buf_data_vac_7;
    wire comm_buf_5_7;
    wire buf_data_vac_6;
    wire buf_data_vac_5;
    wire buf_data_vac_4;
    wire comm_buf_5_4;
    wire buf_data_vac_3;
    wire comm_buf_5_3;
    wire buf_data_vac_2;
    wire comm_buf_5_2;
    wire buf_data_vac_1;
    wire n12431;
    wire n14993;
    wire n11652;
    wire n2_adj_1576_cascade_;
    wire n22611;
    wire comm_state_3_N_460_3;
    wire n1348_cascade_;
    wire n21139_cascade_;
    wire n1348;
    wire n8_adj_1577;
    wire n22614;
    wire n4;
    wire n21013_cascade_;
    wire n21035;
    wire comm_length_0;
    wire n4_adj_1623;
    wire n3;
    wire n21110;
    wire n3_cascade_;
    wire n12442;
    wire n4_adj_1589;
    wire n20095_cascade_;
    wire n21013;
    wire n11619;
    wire n21588;
    wire n9342;
    wire n18070;
    wire n21033;
    wire n7_adj_1650;
    wire comm_cmd_6;
    wire comm_cmd_5;
    wire n4_adj_1455;
    wire n21147;
    wire n21219_cascade_;
    wire n21089;
    wire n21043;
    wire buf_data_vac_16;
    wire comm_rx_buf_0;
    wire comm_buf_3_0;
    wire buf_data_vac_23;
    wire comm_rx_buf_7;
    wire comm_buf_3_7;
    wire buf_data_vac_22;
    wire buf_data_vac_21;
    wire buf_data_vac_20;
    wire comm_buf_3_4;
    wire comm_rx_buf_3;
    wire buf_data_vac_19;
    wire comm_buf_3_3;
    wire buf_data_vac_18;
    wire comm_buf_3_2;
    wire comm_rx_buf_1;
    wire buf_data_vac_17;
    wire comm_buf_5_6;
    wire comm_buf_4_6;
    wire comm_buf_2_6;
    wire comm_buf_3_6;
    wire comm_buf_0_6;
    wire n22545_cascade_;
    wire comm_buf_1_6;
    wire n12353;
    wire n14979;
    wire comm_rx_buf_2;
    wire comm_buf_6_2;
    wire comm_buf_5_0;
    wire comm_buf_4_0;
    wire n4_adj_1457;
    wire comm_buf_5_1;
    wire comm_buf_4_1;
    wire comm_cmd_7;
    wire comm_buf_6_1;
    wire n4_adj_1588;
    wire n21433_cascade_;
    wire n22419_cascade_;
    wire n21085;
    wire n7_adj_1458_cascade_;
    wire n4_adj_1581;
    wire n21282_cascade_;
    wire n22548;
    wire comm_tx_buf_6;
    wire comm_buf_5_5;
    wire comm_buf_1_5;
    wire comm_buf_3_5;
    wire n17698_cascade_;
    wire n21270_cascade_;
    wire n12541;
    wire n15007;
    wire n20996_cascade_;
    wire n12_adj_1663;
    wire n20996;
    wire INVdds0_mclk_294C_net;
    wire clk_16MHz;
    wire dds0_mclk;
    wire buf_control_6;
    wire DDS_MCLK;
    wire acadc_skipcnt_10;
    wire acadc_skipCount_12;
    wire acadc_skipcnt_12;
    wire acadc_skipCount_10;
    wire n21;
    wire n11590;
    wire dds0_mclkcnt_0;
    wire bfn_18_16_0_;
    wire dds0_mclkcnt_1;
    wire n19925;
    wire dds0_mclkcnt_2;
    wire n19926;
    wire dds0_mclkcnt_3;
    wire n19927;
    wire dds0_mclkcnt_4;
    wire n19928;
    wire dds0_mclkcnt_5;
    wire n19929;
    wire n10_adj_1528;
    wire dds0_mclkcnt_6;
    wire n19930;
    wire n19931;
    wire dds0_mclkcnt_7;
    wire INVdds0_mclkcnt_i7_3772__i0C_net;
    wire n14716;
    wire ICE_SPI_MOSI;
    wire \comm_spi.imosi_N_793 ;
    wire \comm_spi.data_tx_7__N_810 ;
    wire \INVADC_VDC.genclk.div_state_i1C_net ;
    wire VDC_SDO;
    wire \ADC_VDC.adc_state_0 ;
    wire adc_state_3;
    wire adc_state_2_adj_1500;
    wire \ADC_VDC.n52_cascade_ ;
    wire \ADC_VDC.adc_state_1 ;
    wire \ADC_VDC.n11905 ;
    wire bfn_19_7_0_;
    wire \ADC_VDC.genclk.n19888 ;
    wire \ADC_VDC.genclk.n19889 ;
    wire \ADC_VDC.genclk.n19890 ;
    wire \ADC_VDC.genclk.n19891 ;
    wire \ADC_VDC.genclk.n19892 ;
    wire \ADC_VDC.genclk.n19893 ;
    wire \ADC_VDC.genclk.n19894 ;
    wire \ADC_VDC.genclk.n19895 ;
    wire \INVADC_VDC.genclk.t0off_i0C_net ;
    wire bfn_19_8_0_;
    wire \ADC_VDC.genclk.n19896 ;
    wire \ADC_VDC.genclk.n19897 ;
    wire \ADC_VDC.genclk.n19898 ;
    wire \ADC_VDC.genclk.n19899 ;
    wire \ADC_VDC.genclk.n19900 ;
    wire \ADC_VDC.genclk.n19901 ;
    wire \ADC_VDC.genclk.n19902 ;
    wire \INVADC_VDC.genclk.t0off_i8C_net ;
    wire \ADC_VDC.genclk.n11900 ;
    wire n14350;
    wire n21453;
    wire n21454_cascade_;
    wire n14_adj_1638;
    wire n21481;
    wire n12089;
    wire comm_length_2;
    wire n6541;
    wire n21154;
    wire comm_data_vld;
    wire ICE_SPI_CE0;
    wire n6401;
    wire n16821;
    wire \comm_spi.n14842 ;
    wire buf_data_iac_18;
    wire n21460;
    wire comm_buf_2_5;
    wire comm_index_2;
    wire comm_index_1;
    wire comm_buf_0_5;
    wire n22503_cascade_;
    wire comm_buf_4_5;
    wire n22506;
    wire comm_tx_buf_5;
    wire \comm_spi.data_tx_7__N_808 ;
    wire comm_rx_buf_4;
    wire comm_buf_6_4;
    wire comm_buf_3_1;
    wire comm_buf_2_1;
    wire n2_adj_1587;
    wire comm_buf_1_1;
    wire comm_buf_0_1;
    wire n1_adj_1586;
    wire comm_rx_buf_5;
    wire comm_buf_6_5;
    wire buf_data_iac_14;
    wire n21547;
    wire comm_rx_buf_6;
    wire n12477;
    wire comm_buf_6_6;
    wire comm_index_0;
    wire n8_adj_1456;
    wire comm_tx_buf_3;
    wire ICE_GPMI_0;
    wire clk_32MHz;
    wire n11600;
    wire n12433;
    wire n10_adj_1619_cascade_;
    wire comm_state_3;
    wire n12079;
    wire comm_state_2;
    wire comm_state_1;
    wire comm_state_0;
    wire n10804;
    wire \ADC_VDC.genclk.t0off_12 ;
    wire \ADC_VDC.genclk.t0off_2 ;
    wire \ADC_VDC.genclk.t0off_7 ;
    wire \ADC_VDC.genclk.t0off_10 ;
    wire \ADC_VDC.genclk.n27_cascade_ ;
    wire \ADC_VDC.genclk.n21598_cascade_ ;
    wire \ADC_VDC.genclk.n6 ;
    wire \ADC_VDC.genclk.t0off_6 ;
    wire \ADC_VDC.genclk.t0off_1 ;
    wire \ADC_VDC.genclk.t0off_4 ;
    wire \ADC_VDC.genclk.t0off_0 ;
    wire \ADC_VDC.genclk.n21600 ;
    wire \ADC_VDC.genclk.n27_adj_1449_cascade_ ;
    wire \ADC_VDC.genclk.n21597 ;
    wire \ADC_VDC.genclk.n21598 ;
    wire \ADC_VDC.genclk.n21597_cascade_ ;
    wire \INVADC_VDC.genclk.div_state_i0C_net ;
    wire \ADC_VDC.genclk.n21603 ;
    wire \ADC_VDC.genclk.t0off_13 ;
    wire \ADC_VDC.genclk.t0off_3 ;
    wire \ADC_VDC.genclk.t0off_5 ;
    wire \ADC_VDC.genclk.t0off_8 ;
    wire \ADC_VDC.genclk.n26 ;
    wire \ADC_VDC.genclk.div_state_0 ;
    wire \ADC_VDC.genclk.n28_adj_1447 ;
    wire \ADC_VDC.genclk.t0off_14 ;
    wire \ADC_VDC.genclk.t0off_9 ;
    wire \ADC_VDC.genclk.t0off_15 ;
    wire \ADC_VDC.genclk.t0off_11 ;
    wire \ADC_VDC.genclk.n28 ;
    wire \ADC_VDC.genclk.n26_adj_1448 ;
    wire \comm_spi.n23101 ;
    wire \comm_spi.n14834 ;
    wire \comm_spi.data_tx_7__N_823 ;
    wire \comm_spi.data_tx_7__N_811 ;
    wire comm_tx_buf_4;
    wire \comm_spi.data_tx_7__N_809 ;
    wire comm_tx_buf_2;
    wire \comm_spi.data_tx_7__N_829 ;
    wire \comm_spi.n23098 ;
    wire \comm_spi.n14838 ;
    wire \comm_spi.n14839 ;
    wire \comm_spi.n14843 ;
    wire \comm_spi.data_tx_7__N_820 ;
    wire \comm_spi.n23104 ;
    wire \comm_spi.n14830 ;
    wire \comm_spi.n14831 ;
    wire \comm_spi.n14835 ;
    wire \comm_spi.data_tx_7__N_826 ;
    wire buf_data_iac_13;
    wire n21456;
    wire buf_data_iac_12;
    wire n21447;
    wire buf_data_iac_9;
    wire n21512;
    wire buf_data_iac_11;
    wire comm_cmd_0;
    wire n21434;
    wire \ADC_VDC.genclk.div_state_1 ;
    wire \ADC_VDC.genclk.t0on_0 ;
    wire bfn_22_7_0_;
    wire \ADC_VDC.genclk.t0on_1 ;
    wire \ADC_VDC.genclk.n19903 ;
    wire \ADC_VDC.genclk.t0on_2 ;
    wire \ADC_VDC.genclk.n19904 ;
    wire \ADC_VDC.genclk.t0on_3 ;
    wire \ADC_VDC.genclk.n19905 ;
    wire \ADC_VDC.genclk.t0on_4 ;
    wire \ADC_VDC.genclk.n19906 ;
    wire \ADC_VDC.genclk.t0on_5 ;
    wire \ADC_VDC.genclk.n19907 ;
    wire \ADC_VDC.genclk.t0on_6 ;
    wire \ADC_VDC.genclk.n19908 ;
    wire \ADC_VDC.genclk.t0on_7 ;
    wire \ADC_VDC.genclk.n19909 ;
    wire \ADC_VDC.genclk.n19910 ;
    wire \INVADC_VDC.genclk.t0on_i0C_net ;
    wire \ADC_VDC.genclk.t0on_8 ;
    wire bfn_22_8_0_;
    wire \ADC_VDC.genclk.t0on_9 ;
    wire \ADC_VDC.genclk.n19911 ;
    wire \ADC_VDC.genclk.t0on_10 ;
    wire \ADC_VDC.genclk.n19912 ;
    wire \ADC_VDC.genclk.t0on_11 ;
    wire \ADC_VDC.genclk.n19913 ;
    wire \ADC_VDC.genclk.t0on_12 ;
    wire \ADC_VDC.genclk.n19914 ;
    wire \ADC_VDC.genclk.t0on_13 ;
    wire \ADC_VDC.genclk.n19915 ;
    wire \ADC_VDC.genclk.t0on_14 ;
    wire \ADC_VDC.genclk.n19916 ;
    wire \ADC_VDC.genclk.n19917 ;
    wire \ADC_VDC.genclk.t0on_15 ;
    wire \INVADC_VDC.genclk.t0on_i8C_net ;
    wire \ADC_VDC.genclk.div_state_1__N_1432 ;
    wire \ADC_VDC.genclk.n14894 ;
    wire \comm_spi.data_tx_7__N_835 ;
    wire \comm_spi.n14827 ;
    wire \comm_spi.n23110 ;
    wire \comm_spi.n14801 ;
    wire \comm_spi.n14826 ;
    wire \comm_spi.data_tx_7__N_812 ;
    wire \comm_spi.data_tx_7__N_832 ;
    wire comm_tx_buf_1;
    wire \comm_spi.n23107 ;
    wire CONSTANT_ONE_NET;
    wire \comm_spi.n14800 ;
    wire \comm_spi.iclk ;
    wire comm_tx_buf_0;
    wire comm_clear;
    wire \comm_spi.data_tx_7__N_813 ;
    wire _gnd_net_;

    defparam \pll_main.zim_pll_inst .DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam \pll_main.zim_pll_inst .TEST_MODE=1'b0;
    defparam \pll_main.zim_pll_inst .SHIFTREG_DIV_MODE=2'b00;
    defparam \pll_main.zim_pll_inst .PLLOUT_SELECT_PORTB="GENCLK_HALF";
    defparam \pll_main.zim_pll_inst .PLLOUT_SELECT_PORTA="GENCLK";
    defparam \pll_main.zim_pll_inst .FILTER_RANGE=3'b011;
    defparam \pll_main.zim_pll_inst .FEEDBACK_PATH="SIMPLE";
    defparam \pll_main.zim_pll_inst .FDA_RELATIVE=4'b0000;
    defparam \pll_main.zim_pll_inst .FDA_FEEDBACK=4'b0000;
    defparam \pll_main.zim_pll_inst .ENABLE_ICEGATE_PORTB=1'b0;
    defparam \pll_main.zim_pll_inst .ENABLE_ICEGATE_PORTA=1'b0;
    defparam \pll_main.zim_pll_inst .DIVR=4'b0000;
    defparam \pll_main.zim_pll_inst .DIVQ=3'b101;
    defparam \pll_main.zim_pll_inst .DIVF=7'b0011111;
    defparam \pll_main.zim_pll_inst .DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_2F_CORE \pll_main.zim_pll_inst  (
            .EXTFEEDBACK(GNDG0),
            .SDO(),
            .LOCK(),
            .PLLOUTCOREB(),
            .REFERENCECLK(N__19413),
            .RESETB(N__58773),
            .BYPASS(GNDG0),
            .PLLOUTCOREA(),
            .SDI(GNDG0),
            .PLLOUTGLOBALB(clk_16MHz),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .LATCHINPUTVALUE(GNDG0),
            .PLLOUTGLOBALA(clk_32MHz),
            .SCLK(GNDG0));
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged2_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged2_physical (
            .RDATA({dangling_wire_0,dangling_wire_1,buf_data_iac_19,dangling_wire_2,dangling_wire_3,dangling_wire_4,buf_data_vac_19,dangling_wire_5,dangling_wire_6,dangling_wire_7,buf_data_iac_18,dangling_wire_8,dangling_wire_9,dangling_wire_10,buf_data_vac_18,dangling_wire_11}),
            .RADDR({dangling_wire_12,N__41862,N__39420,N__32922,N__36093,N__41382,N__36414,N__35943,N__39879,N__39288,N__41010}),
            .WADDR({dangling_wire_13,N__33885,N__33996,N__34104,N__34212,N__33198,N__33300,N__33411,N__33522,N__33630,N__33732}),
            .MASK({dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25,dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29}),
            .WDATA({dangling_wire_30,dangling_wire_31,N__26472,dangling_wire_32,dangling_wire_33,dangling_wire_34,N__25980,dangling_wire_35,dangling_wire_36,dangling_wire_37,N__32763,dangling_wire_38,dangling_wire_39,dangling_wire_40,N__24138,dangling_wire_41}),
            .RCLKE(),
            .RCLK(N__56042),
            .RE(N__58486),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged2WCLKN_net),
            .WE(N__28614));
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged7_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged7_physical (
            .RDATA({dangling_wire_42,dangling_wire_43,buf_data_iac_9,dangling_wire_44,dangling_wire_45,dangling_wire_46,buf_data_vac_9,dangling_wire_47,dangling_wire_48,dangling_wire_49,buf_data_iac_8,dangling_wire_50,dangling_wire_51,dangling_wire_52,buf_data_vac_8,dangling_wire_53}),
            .RADDR({dangling_wire_54,N__41822,N__39380,N__32885,N__36047,N__41336,N__36377,N__35906,N__39836,N__39245,N__40967}),
            .WADDR({dangling_wire_55,N__33848,N__33956,N__34058,N__34172,N__33155,N__33266,N__33374,N__33485,N__33590,N__33692}),
            .MASK({dangling_wire_56,dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71}),
            .WDATA({dangling_wire_72,dangling_wire_73,N__43620,dangling_wire_74,dangling_wire_75,dangling_wire_76,N__23568,dangling_wire_77,dangling_wire_78,dangling_wire_79,N__41706,dangling_wire_80,dangling_wire_81,dangling_wire_82,N__43758,dangling_wire_83}),
            .RCLKE(),
            .RCLK(N__56102),
            .RE(N__58776),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged7WCLKN_net),
            .WE(N__28626));
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged1_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged1_physical (
            .RDATA({dangling_wire_84,dangling_wire_85,buf_data_iac_21,dangling_wire_86,dangling_wire_87,dangling_wire_88,buf_data_vac_21,dangling_wire_89,dangling_wire_90,dangling_wire_91,buf_data_iac_20,dangling_wire_92,dangling_wire_93,dangling_wire_94,buf_data_vac_20,dangling_wire_95}),
            .RADDR({dangling_wire_96,N__41880,N__39438,N__32940,N__36111,N__41400,N__36432,N__35961,N__39897,N__39306,N__41028}),
            .WADDR({dangling_wire_97,N__33903,N__34014,N__34122,N__34230,N__33216,N__33318,N__33429,N__33540,N__33648,N__33750}),
            .MASK({dangling_wire_98,dangling_wire_99,dangling_wire_100,dangling_wire_101,dangling_wire_102,dangling_wire_103,dangling_wire_104,dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,dangling_wire_109,dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113}),
            .WDATA({dangling_wire_114,dangling_wire_115,N__28947,dangling_wire_116,dangling_wire_117,dangling_wire_118,N__27429,dangling_wire_119,dangling_wire_120,dangling_wire_121,N__32148,dangling_wire_122,dangling_wire_123,dangling_wire_124,N__31884,dangling_wire_125}),
            .RCLKE(),
            .RCLK(N__55962),
            .RE(N__58762),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged1WCLKN_net),
            .WE(N__28631));
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged6_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged6_physical (
            .RDATA({dangling_wire_126,dangling_wire_127,buf_data_iac_11,dangling_wire_128,dangling_wire_129,dangling_wire_130,buf_data_vac_11,dangling_wire_131,dangling_wire_132,dangling_wire_133,buf_data_iac_10,dangling_wire_134,dangling_wire_135,dangling_wire_136,buf_data_vac_10,dangling_wire_137}),
            .RADDR({dangling_wire_138,N__41834,N__39392,N__32897,N__36059,N__41348,N__36389,N__35918,N__39848,N__39257,N__40979}),
            .WADDR({dangling_wire_139,N__33860,N__33968,N__34070,N__34184,N__33167,N__33276,N__33386,N__33497,N__33602,N__33704}),
            .MASK({dangling_wire_140,dangling_wire_141,dangling_wire_142,dangling_wire_143,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,dangling_wire_151,dangling_wire_152,dangling_wire_153,dangling_wire_154,dangling_wire_155}),
            .WDATA({dangling_wire_156,dangling_wire_157,N__41303,dangling_wire_158,dangling_wire_159,dangling_wire_160,N__35052,dangling_wire_161,dangling_wire_162,dangling_wire_163,N__38237,dangling_wire_164,dangling_wire_165,dangling_wire_166,N__27333,dangling_wire_167}),
            .RCLKE(),
            .RCLK(N__56100),
            .RE(N__58775),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged6WCLKN_net),
            .WE(N__28621));
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged0_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged0_physical (
            .RDATA({dangling_wire_168,dangling_wire_169,buf_data_iac_23,dangling_wire_170,dangling_wire_171,dangling_wire_172,buf_data_vac_23,dangling_wire_173,dangling_wire_174,dangling_wire_175,buf_data_iac_22,dangling_wire_176,dangling_wire_177,dangling_wire_178,buf_data_vac_22,dangling_wire_179}),
            .RADDR({dangling_wire_180,N__41886,N__39444,N__32946,N__36117,N__41406,N__36438,N__35967,N__39903,N__39312,N__41034}),
            .WADDR({dangling_wire_181,N__33909,N__34020,N__34128,N__34236,N__33222,N__33324,N__33435,N__33546,N__33654,N__33756}),
            .MASK({dangling_wire_182,dangling_wire_183,dangling_wire_184,dangling_wire_185,dangling_wire_186,dangling_wire_187,dangling_wire_188,dangling_wire_189,dangling_wire_190,dangling_wire_191,dangling_wire_192,dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197}),
            .WDATA({dangling_wire_198,dangling_wire_199,N__29201,dangling_wire_200,dangling_wire_201,dangling_wire_202,N__27120,dangling_wire_203,dangling_wire_204,dangling_wire_205,N__30779,dangling_wire_206,dangling_wire_207,dangling_wire_208,N__23109,dangling_wire_209}),
            .RCLKE(),
            .RCLK(N__55948),
            .RE(N__58763),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged0WCLKN_net),
            .WE(N__28632));
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged5_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged5_physical (
            .RDATA({dangling_wire_210,dangling_wire_211,buf_data_iac_13,dangling_wire_212,dangling_wire_213,dangling_wire_214,buf_data_vac_13,dangling_wire_215,dangling_wire_216,dangling_wire_217,buf_data_iac_12,dangling_wire_218,dangling_wire_219,dangling_wire_220,buf_data_vac_12,dangling_wire_221}),
            .RADDR({dangling_wire_222,N__41844,N__39402,N__32904,N__36071,N__41360,N__36396,N__35925,N__39860,N__39269,N__40991}),
            .WADDR({dangling_wire_223,N__33867,N__33978,N__34082,N__34194,N__33179,N__33282,N__33393,N__33504,N__33612,N__33714}),
            .MASK({dangling_wire_224,dangling_wire_225,dangling_wire_226,dangling_wire_227,dangling_wire_228,dangling_wire_229,dangling_wire_230,dangling_wire_231,dangling_wire_232,dangling_wire_233,dangling_wire_234,dangling_wire_235,dangling_wire_236,dangling_wire_237,dangling_wire_238,dangling_wire_239}),
            .WDATA({dangling_wire_240,dangling_wire_241,N__33079,dangling_wire_242,dangling_wire_243,dangling_wire_244,N__28320,dangling_wire_245,dangling_wire_246,dangling_wire_247,N__30609,dangling_wire_248,dangling_wire_249,dangling_wire_250,N__27486,dangling_wire_251}),
            .RCLKE(),
            .RCLK(N__56097),
            .RE(N__58766),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged5WCLKN_net),
            .WE(N__28610));
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged9_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged9_physical (
            .RDATA({dangling_wire_252,dangling_wire_253,buf_data_iac_5,dangling_wire_254,dangling_wire_255,dangling_wire_256,buf_data_vac_5,dangling_wire_257,dangling_wire_258,dangling_wire_259,buf_data_iac_4,dangling_wire_260,dangling_wire_261,dangling_wire_262,buf_data_vac_4,dangling_wire_263}),
            .RADDR({dangling_wire_264,N__41831,N__39389,N__32888,N__36068,N__41357,N__36380,N__35909,N__39851,N__39260,N__40982}),
            .WADDR({dangling_wire_265,N__33851,N__33965,N__34079,N__34181,N__33170,N__33263,N__33377,N__33488,N__33599,N__33701}),
            .MASK({dangling_wire_266,dangling_wire_267,dangling_wire_268,dangling_wire_269,dangling_wire_270,dangling_wire_271,dangling_wire_272,dangling_wire_273,dangling_wire_274,dangling_wire_275,dangling_wire_276,dangling_wire_277,dangling_wire_278,dangling_wire_279,dangling_wire_280,dangling_wire_281}),
            .WDATA({dangling_wire_282,dangling_wire_283,N__24237,dangling_wire_284,dangling_wire_285,dangling_wire_286,N__24264,dangling_wire_287,dangling_wire_288,dangling_wire_289,N__21315,dangling_wire_290,dangling_wire_291,dangling_wire_292,N__21288,dangling_wire_293}),
            .RCLKE(),
            .RCLK(N__55997),
            .RE(N__58758),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged9WCLKN_net),
            .WE(N__28571));
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged4_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged4_physical (
            .RDATA({dangling_wire_294,dangling_wire_295,buf_data_iac_15,dangling_wire_296,dangling_wire_297,dangling_wire_298,buf_data_vac_15,dangling_wire_299,dangling_wire_300,dangling_wire_301,buf_data_iac_14,dangling_wire_302,dangling_wire_303,dangling_wire_304,buf_data_vac_14,dangling_wire_305}),
            .RADDR({dangling_wire_306,N__41850,N__39408,N__32910,N__36081,N__41370,N__36402,N__35931,N__39867,N__39276,N__40998}),
            .WADDR({dangling_wire_307,N__33873,N__33984,N__34092,N__34200,N__33186,N__33288,N__33399,N__33510,N__33618,N__33720}),
            .MASK({dangling_wire_308,dangling_wire_309,dangling_wire_310,dangling_wire_311,dangling_wire_312,dangling_wire_313,dangling_wire_314,dangling_wire_315,dangling_wire_316,dangling_wire_317,dangling_wire_318,dangling_wire_319,dangling_wire_320,dangling_wire_321,dangling_wire_322,dangling_wire_323}),
            .WDATA({dangling_wire_324,dangling_wire_325,N__42054,dangling_wire_326,dangling_wire_327,dangling_wire_328,N__28440,dangling_wire_329,dangling_wire_330,dangling_wire_331,N__43392,dangling_wire_332,dangling_wire_333,dangling_wire_334,N__32472,dangling_wire_335}),
            .RCLKE(),
            .RCLK(N__56090),
            .RE(N__58764),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged4WCLKN_net),
            .WE(N__28575));
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged8_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged8_physical (
            .RDATA({dangling_wire_336,dangling_wire_337,buf_data_iac_7,dangling_wire_338,dangling_wire_339,dangling_wire_340,buf_data_vac_7,dangling_wire_341,dangling_wire_342,dangling_wire_343,buf_data_iac_6,dangling_wire_344,dangling_wire_345,dangling_wire_346,buf_data_vac_6,dangling_wire_347}),
            .RADDR({dangling_wire_348,N__41843,N__39401,N__32900,N__36080,N__41369,N__36392,N__35921,N__39863,N__39272,N__40994}),
            .WADDR({dangling_wire_349,N__33863,N__33977,N__34091,N__34193,N__33182,N__33275,N__33389,N__33500,N__33611,N__33713}),
            .MASK({dangling_wire_350,dangling_wire_351,dangling_wire_352,dangling_wire_353,dangling_wire_354,dangling_wire_355,dangling_wire_356,dangling_wire_357,dangling_wire_358,dangling_wire_359,dangling_wire_360,dangling_wire_361,dangling_wire_362,dangling_wire_363,dangling_wire_364,dangling_wire_365}),
            .WDATA({dangling_wire_366,dangling_wire_367,N__21405,dangling_wire_368,dangling_wire_369,dangling_wire_370,N__20040,dangling_wire_371,dangling_wire_372,dangling_wire_373,N__20841,dangling_wire_374,dangling_wire_375,dangling_wire_376,N__23142,dangling_wire_377}),
            .RCLKE(),
            .RCLK(N__55972),
            .RE(N__58774),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged8WCLKN_net),
            .WE(N__28602));
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged10_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged10_physical (
            .RDATA({dangling_wire_378,dangling_wire_379,buf_data_iac_3,dangling_wire_380,dangling_wire_381,dangling_wire_382,buf_data_vac_3,dangling_wire_383,dangling_wire_384,dangling_wire_385,buf_data_iac_2,dangling_wire_386,dangling_wire_387,dangling_wire_388,buf_data_vac_2,dangling_wire_389}),
            .RADDR({dangling_wire_390,N__41874,N__39432,N__32934,N__36105,N__41394,N__36426,N__35955,N__39891,N__39300,N__41022}),
            .WADDR({dangling_wire_391,N__33897,N__34008,N__34116,N__34224,N__33210,N__33312,N__33423,N__33534,N__33642,N__33744}),
            .MASK({dangling_wire_392,dangling_wire_393,dangling_wire_394,dangling_wire_395,dangling_wire_396,dangling_wire_397,dangling_wire_398,dangling_wire_399,dangling_wire_400,dangling_wire_401,dangling_wire_402,dangling_wire_403,dangling_wire_404,dangling_wire_405,dangling_wire_406,dangling_wire_407}),
            .WDATA({dangling_wire_408,dangling_wire_409,N__22857,dangling_wire_410,dangling_wire_411,dangling_wire_412,N__23268,dangling_wire_413,dangling_wire_414,dangling_wire_415,N__24300,dangling_wire_416,dangling_wire_417,dangling_wire_418,N__23169,dangling_wire_419}),
            .RCLKE(),
            .RCLK(N__55984),
            .RE(N__58720),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged10WCLKN_net),
            .WE(N__28627));
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged3_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged3_physical (
            .RDATA({dangling_wire_420,dangling_wire_421,buf_data_iac_17,dangling_wire_422,dangling_wire_423,dangling_wire_424,buf_data_vac_17,dangling_wire_425,dangling_wire_426,dangling_wire_427,buf_data_iac_16,dangling_wire_428,dangling_wire_429,dangling_wire_430,buf_data_vac_16,dangling_wire_431}),
            .RADDR({dangling_wire_432,N__41856,N__39414,N__32916,N__36087,N__41376,N__36408,N__35937,N__39873,N__39282,N__41004}),
            .WADDR({dangling_wire_433,N__33879,N__33990,N__34098,N__34206,N__33192,N__33294,N__33405,N__33516,N__33624,N__33726}),
            .MASK({dangling_wire_434,dangling_wire_435,dangling_wire_436,dangling_wire_437,dangling_wire_438,dangling_wire_439,dangling_wire_440,dangling_wire_441,dangling_wire_442,dangling_wire_443,dangling_wire_444,dangling_wire_445,dangling_wire_446,dangling_wire_447,dangling_wire_448,dangling_wire_449}),
            .WDATA({dangling_wire_450,dangling_wire_451,N__24759,dangling_wire_452,dangling_wire_453,dangling_wire_454,N__24528,dangling_wire_455,dangling_wire_456,dangling_wire_457,N__39143,dangling_wire_458,dangling_wire_459,dangling_wire_460,N__25782,dangling_wire_461}),
            .RCLKE(),
            .RCLK(N__56071),
            .RE(N__58728),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged3WCLKN_net),
            .WE(N__28603));
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.WRITE_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.READ_MODE=2;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_F=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_E=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_D=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_C=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_B=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_A=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_9=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_8=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_7=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_6=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_5=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_4=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_3=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_2=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_1=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    defparam iac_raw_buf_vac_raw_buf_merged11_physical.INIT_0=256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    SB_RAM40_4K iac_raw_buf_vac_raw_buf_merged11_physical (
            .RDATA({dangling_wire_462,dangling_wire_463,buf_data_iac_1,dangling_wire_464,dangling_wire_465,dangling_wire_466,buf_data_vac_1,dangling_wire_467,dangling_wire_468,dangling_wire_469,buf_data_iac_0,dangling_wire_470,dangling_wire_471,dangling_wire_472,buf_data_vac_0,dangling_wire_473}),
            .RADDR({dangling_wire_474,N__41868,N__39426,N__32928,N__36099,N__41388,N__36420,N__35949,N__39885,N__39294,N__41016}),
            .WADDR({dangling_wire_475,N__33891,N__34002,N__34110,N__34218,N__33204,N__33306,N__33417,N__33528,N__33636,N__33738}),
            .MASK({dangling_wire_476,dangling_wire_477,dangling_wire_478,dangling_wire_479,dangling_wire_480,dangling_wire_481,dangling_wire_482,dangling_wire_483,dangling_wire_484,dangling_wire_485,dangling_wire_486,dangling_wire_487,dangling_wire_488,dangling_wire_489,dangling_wire_490,dangling_wire_491}),
            .WDATA({dangling_wire_492,dangling_wire_493,N__36315,dangling_wire_494,dangling_wire_495,dangling_wire_496,N__32184,dangling_wire_497,dangling_wire_498,dangling_wire_499,N__27237,dangling_wire_500,dangling_wire_501,dangling_wire_502,N__27273,dangling_wire_503}),
            .RCLKE(),
            .RCLK(N__56012),
            .RE(N__58719),
            .WCLKE(),
            .WCLK(INViac_raw_buf_vac_raw_buf_merged11WCLKN_net),
            .WE(N__28622));
    IO_PAD ipInertedIOPad_VAC_DRDY_iopad (
            .OE(N__59914),
            .DIN(N__59913),
            .DOUT(N__59912),
            .PACKAGEPIN(VAC_DRDY));
    defparam ipInertedIOPad_VAC_DRDY_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VAC_DRDY_preio (
            .PADOEN(N__59914),
            .PADOUT(N__59913),
            .PADIN(N__59912),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(VAC_DRDY),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_FLT1_iopad (
            .OE(N__59905),
            .DIN(N__59904),
            .DOUT(N__59903),
            .PACKAGEPIN(IAC_FLT1));
    defparam ipInertedIOPad_IAC_FLT1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_FLT1_preio (
            .PADOEN(N__59905),
            .PADOUT(N__59904),
            .PADIN(N__59903),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__26502),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_SCK_iopad (
            .OE(N__59896),
            .DIN(N__59895),
            .DOUT(N__59894),
            .PACKAGEPIN(DDS_SCK));
    defparam ipInertedIOPad_DDS_SCK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_SCK_preio (
            .PADOEN(N__59896),
            .PADOUT(N__59895),
            .PADIN(N__59894),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__39036),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_166_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_166_iopad (
            .OE(N__59887),
            .DIN(N__59886),
            .DOUT(N__59885),
            .PACKAGEPIN(ICE_IOR_166));
    defparam ipInertedIOPad_ICE_IOR_166_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_166_preio (
            .PADOEN(N__59887),
            .PADOUT(N__59886),
            .PADIN(N__59885),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_119_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_119_iopad (
            .OE(N__59878),
            .DIN(N__59877),
            .DOUT(N__59876),
            .PACKAGEPIN(ICE_IOR_119));
    defparam ipInertedIOPad_ICE_IOR_119_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_119_preio (
            .PADOEN(N__59878),
            .PADOUT(N__59877),
            .PADIN(N__59876),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_MOSI_iopad (
            .OE(N__59869),
            .DIN(N__59868),
            .DOUT(N__59867),
            .PACKAGEPIN(DDS_MOSI));
    defparam ipInertedIOPad_DDS_MOSI_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_MOSI_preio (
            .PADOEN(N__59869),
            .PADOUT(N__59868),
            .PADIN(N__59867),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__38985),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_MISO_iopad (
            .OE(N__59860),
            .DIN(N__59859),
            .DOUT(N__59858),
            .PACKAGEPIN(VAC_MISO));
    defparam ipInertedIOPad_VAC_MISO_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VAC_MISO_preio (
            .PADOEN(N__59860),
            .PADOUT(N__59859),
            .PADIN(N__59858),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(VAC_MISO),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_MOSI1_iopad (
            .OE(N__59851),
            .DIN(N__59850),
            .DOUT(N__59849),
            .PACKAGEPIN(DDS_MOSI1));
    defparam ipInertedIOPad_DDS_MOSI1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_MOSI1_preio (
            .PADOEN(N__59851),
            .PADOUT(N__59850),
            .PADIN(N__59849),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__22773),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_146_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_146_iopad (
            .OE(N__59842),
            .DIN(N__59841),
            .DOUT(N__59840),
            .PACKAGEPIN(ICE_IOR_146));
    defparam ipInertedIOPad_ICE_IOR_146_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_146_preio (
            .PADOEN(N__59842),
            .PADOUT(N__59841),
            .PADIN(N__59840),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VDC_CLK_iopad (
            .OE(N__59833),
            .DIN(N__59832),
            .DOUT(N__59831),
            .PACKAGEPIN(VDC_CLK));
    defparam ipInertedIOPad_VDC_CLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VDC_CLK_preio (
            .PADOEN(N__59833),
            .PADOUT(N__59832),
            .PADIN(N__59831),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__42435),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_222_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_222_iopad (
            .OE(N__59824),
            .DIN(N__59823),
            .DOUT(N__59822),
            .PACKAGEPIN(ICE_IOT_222));
    defparam ipInertedIOPad_ICE_IOT_222_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_222_preio (
            .PADOEN(N__59824),
            .PADOUT(N__59823),
            .PADIN(N__59822),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_CS_iopad (
            .OE(N__59815),
            .DIN(N__59814),
            .DOUT(N__59813),
            .PACKAGEPIN(IAC_CS));
    defparam ipInertedIOPad_IAC_CS_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_CS_preio (
            .PADOEN(N__59815),
            .PADOUT(N__59814),
            .PADIN(N__59813),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__21879),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_18B_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_18B_iopad (
            .OE(N__59806),
            .DIN(N__59805),
            .DOUT(N__59804),
            .PACKAGEPIN(ICE_IOL_18B));
    defparam ipInertedIOPad_ICE_IOL_18B_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_18B_preio (
            .PADOEN(N__59806),
            .PADOUT(N__59805),
            .PADIN(N__59804),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_13A_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_13A_iopad (
            .OE(N__59797),
            .DIN(N__59796),
            .DOUT(N__59795),
            .PACKAGEPIN(ICE_IOL_13A));
    defparam ipInertedIOPad_ICE_IOL_13A_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_13A_preio (
            .PADOEN(N__59797),
            .PADOUT(N__59796),
            .PADIN(N__59795),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_ICE_IOB_81_iopad (
            .OE(N__59788),
            .DIN(N__59787),
            .DOUT(N__59786),
            .PACKAGEPIN(ICE_IOB_81));
    defparam ipInertedIOPad_ICE_IOB_81_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_81_preio (
            .PADOEN(N__59788),
            .PADOUT(N__59787),
            .PADIN(N__59786),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_OSR1_iopad (
            .OE(N__59779),
            .DIN(N__59778),
            .DOUT(N__59777),
            .PACKAGEPIN(VAC_OSR1));
    defparam ipInertedIOPad_VAC_OSR1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_OSR1_preio (
            .PADOEN(N__59779),
            .PADOUT(N__59778),
            .PADIN(N__59777),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__27390),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_MOSI_iopad (
            .OE(N__59770),
            .DIN(N__59769),
            .DOUT(N__59768),
            .PACKAGEPIN(IAC_MOSI));
    defparam ipInertedIOPad_IAC_MOSI_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_MOSI_preio (
            .PADOEN(N__59770),
            .PADOUT(N__59769),
            .PADIN(N__59768),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_CS1_iopad (
            .OE(N__59761),
            .DIN(N__59760),
            .DOUT(N__59759),
            .PACKAGEPIN(DDS_CS1));
    defparam ipInertedIOPad_DDS_CS1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_CS1_preio (
            .PADOEN(N__59761),
            .PADOUT(N__59760),
            .PADIN(N__59759),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__21858),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_4B_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_4B_iopad (
            .OE(N__59752),
            .DIN(N__59751),
            .DOUT(N__59750),
            .PACKAGEPIN(ICE_IOL_4B));
    defparam ipInertedIOPad_ICE_IOL_4B_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_4B_preio (
            .PADOEN(N__59752),
            .PADOUT(N__59751),
            .PADIN(N__59750),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOB_94_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOB_94_iopad (
            .OE(N__59743),
            .DIN(N__59742),
            .DOUT(N__59741),
            .PACKAGEPIN(ICE_IOB_94));
    defparam ipInertedIOPad_ICE_IOB_94_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_94_preio (
            .PADOEN(N__59743),
            .PADOUT(N__59742),
            .PADIN(N__59741),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_CS_iopad (
            .OE(N__59734),
            .DIN(N__59733),
            .DOUT(N__59732),
            .PACKAGEPIN(VAC_CS));
    defparam ipInertedIOPad_VAC_CS_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_CS_preio (
            .PADOEN(N__59734),
            .PADOUT(N__59733),
            .PADIN(N__59732),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__21660),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_CLK_iopad (
            .OE(N__59725),
            .DIN(N__59724),
            .DOUT(N__59723),
            .PACKAGEPIN(VAC_CLK));
    defparam ipInertedIOPad_VAC_CLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_CLK_preio (
            .PADOEN(N__59725),
            .PADOUT(N__59724),
            .PADIN(N__59723),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__31121),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_SPI_CE0_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_SPI_CE0_iopad (
            .OE(N__59716),
            .DIN(N__59715),
            .DOUT(N__59714),
            .PACKAGEPIN(ICE_SPI_CE0));
    defparam ipInertedIOPad_ICE_SPI_CE0_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_SPI_CE0_preio (
            .PADOEN(N__59716),
            .PADOUT(N__59715),
            .PADIN(N__59714),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(ICE_SPI_CE0),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_167_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_167_iopad (
            .OE(N__59707),
            .DIN(N__59706),
            .DOUT(N__59705),
            .PACKAGEPIN(ICE_IOR_167));
    defparam ipInertedIOPad_ICE_IOR_167_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_167_preio (
            .PADOEN(N__59707),
            .PADOUT(N__59706),
            .PADIN(N__59705),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_118_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_118_iopad (
            .OE(N__59698),
            .DIN(N__59697),
            .DOUT(N__59696),
            .PACKAGEPIN(ICE_IOR_118));
    defparam ipInertedIOPad_ICE_IOR_118_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_118_preio (
            .PADOEN(N__59698),
            .PADOUT(N__59697),
            .PADIN(N__59696),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_RTD_SDO_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_RTD_SDO_iopad (
            .OE(N__59689),
            .DIN(N__59688),
            .DOUT(N__59687),
            .PACKAGEPIN(RTD_SDO));
    defparam ipInertedIOPad_RTD_SDO_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_RTD_SDO_preio (
            .PADOEN(N__59689),
            .PADOUT(N__59688),
            .PADIN(N__59687),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(RTD_SDO),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_OSR0_iopad (
            .OE(N__59680),
            .DIN(N__59679),
            .DOUT(N__59678),
            .PACKAGEPIN(IAC_OSR0));
    defparam ipInertedIOPad_IAC_OSR0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_OSR0_preio (
            .PADOEN(N__59680),
            .PADOUT(N__59679),
            .PADIN(N__59678),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__39474),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VDC_SCLK_iopad (
            .OE(N__59671),
            .DIN(N__59670),
            .DOUT(N__59669),
            .PACKAGEPIN(VDC_SCLK));
    defparam ipInertedIOPad_VDC_SCLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VDC_SCLK_preio (
            .PADOEN(N__59671),
            .PADOUT(N__59670),
            .PADIN(N__59669),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__42462),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_FLT1_iopad (
            .OE(N__59662),
            .DIN(N__59661),
            .DOUT(N__59660),
            .PACKAGEPIN(VAC_FLT1));
    defparam ipInertedIOPad_VAC_FLT1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_FLT1_preio (
            .PADOEN(N__59662),
            .PADOUT(N__59661),
            .PADIN(N__59660),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__29007),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_SPI_MOSI_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_SPI_MOSI_iopad (
            .OE(N__59653),
            .DIN(N__59652),
            .DOUT(N__59651),
            .PACKAGEPIN(ICE_SPI_MOSI));
    defparam ipInertedIOPad_ICE_SPI_MOSI_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_SPI_MOSI_preio (
            .PADOEN(N__59653),
            .PADOUT(N__59652),
            .PADIN(N__59651),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(ICE_SPI_MOSI),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_165_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_165_iopad (
            .OE(N__59644),
            .DIN(N__59643),
            .DOUT(N__59642),
            .PACKAGEPIN(ICE_IOR_165));
    defparam ipInertedIOPad_ICE_IOR_165_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_165_preio (
            .PADOEN(N__59644),
            .PADOUT(N__59643),
            .PADIN(N__59642),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_147_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_147_iopad (
            .OE(N__59635),
            .DIN(N__59634),
            .DOUT(N__59633),
            .PACKAGEPIN(ICE_IOR_147));
    defparam ipInertedIOPad_ICE_IOR_147_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_147_preio (
            .PADOEN(N__59635),
            .PADOUT(N__59634),
            .PADIN(N__59633),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_14A_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_14A_iopad (
            .OE(N__59626),
            .DIN(N__59625),
            .DOUT(N__59624),
            .PACKAGEPIN(ICE_IOL_14A));
    defparam ipInertedIOPad_ICE_IOL_14A_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_14A_preio (
            .PADOEN(N__59626),
            .PADOUT(N__59625),
            .PADIN(N__59624),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_13B_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_13B_iopad (
            .OE(N__59617),
            .DIN(N__59616),
            .DOUT(N__59615),
            .PACKAGEPIN(ICE_IOL_13B));
    defparam ipInertedIOPad_ICE_IOL_13B_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_13B_preio (
            .PADOEN(N__59617),
            .PADOUT(N__59616),
            .PADIN(N__59615),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOB_91_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOB_91_iopad (
            .OE(N__59608),
            .DIN(N__59607),
            .DOUT(N__59606),
            .PACKAGEPIN(ICE_IOB_91));
    defparam ipInertedIOPad_ICE_IOB_91_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_91_preio (
            .PADOEN(N__59608),
            .PADOUT(N__59607),
            .PADIN(N__59606),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_GPMO_0_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_GPMO_0_iopad (
            .OE(N__59599),
            .DIN(N__59598),
            .DOUT(N__59597),
            .PACKAGEPIN(ICE_GPMO_0));
    defparam ipInertedIOPad_ICE_GPMO_0_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_GPMO_0_preio (
            .PADOEN(N__59599),
            .PADOUT(N__59598),
            .PADIN(N__59597),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_RNG_0_iopad (
            .OE(N__59590),
            .DIN(N__59589),
            .DOUT(N__59588),
            .PACKAGEPIN(DDS_RNG_0));
    defparam ipInertedIOPad_DDS_RNG_0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_RNG_0_preio (
            .PADOEN(N__59590),
            .PADOUT(N__59589),
            .PADIN(N__59588),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__42957),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VDC_RNG0_iopad (
            .OE(N__59581),
            .DIN(N__59580),
            .DOUT(N__59579),
            .PACKAGEPIN(VDC_RNG0));
    defparam ipInertedIOPad_VDC_RNG0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VDC_RNG0_preio (
            .PADOEN(N__59581),
            .PADOUT(N__59580),
            .PADIN(N__59579),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__41517),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_SPI_SCLK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_SPI_SCLK_iopad (
            .OE(N__59572),
            .DIN(N__59571),
            .DOUT(N__59570),
            .PACKAGEPIN(ICE_SPI_SCLK));
    defparam ipInertedIOPad_ICE_SPI_SCLK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_SPI_SCLK_preio (
            .PADOEN(N__59572),
            .PADOUT(N__59571),
            .PADIN(N__59570),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(ICE_SPI_SCLK),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_152_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_152_iopad (
            .OE(N__59563),
            .DIN(N__59562),
            .DOUT(N__59561),
            .PACKAGEPIN(ICE_IOR_152));
    defparam ipInertedIOPad_ICE_IOR_152_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_152_preio (
            .PADOEN(N__59563),
            .PADOUT(N__59562),
            .PADIN(N__59561),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_12A_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_12A_iopad (
            .OE(N__59554),
            .DIN(N__59553),
            .DOUT(N__59552),
            .PACKAGEPIN(ICE_IOL_12A));
    defparam ipInertedIOPad_ICE_IOL_12A_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_12A_preio (
            .PADOEN(N__59554),
            .PADOUT(N__59553),
            .PADIN(N__59552),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_RTD_DRDY_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_RTD_DRDY_iopad (
            .OE(N__59545),
            .DIN(N__59544),
            .DOUT(N__59543),
            .PACKAGEPIN(RTD_DRDY));
    defparam ipInertedIOPad_RTD_DRDY_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_RTD_DRDY_preio (
            .PADOEN(N__59545),
            .PADOUT(N__59544),
            .PADIN(N__59543),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(RTD_DRDY),
            .DIN1());
    IO_PAD ipInertedIOPad_ICE_SPI_MISO_iopad (
            .OE(N__59536),
            .DIN(N__59535),
            .DOUT(N__59534),
            .PACKAGEPIN(ICE_SPI_MISO));
    defparam ipInertedIOPad_ICE_SPI_MISO_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_ICE_SPI_MISO_preio (
            .PADOEN(N__59536),
            .PADOUT(N__59535),
            .PADIN(N__59534),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__44283),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_177_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_177_iopad (
            .OE(N__59527),
            .DIN(N__59526),
            .DOUT(N__59525),
            .PACKAGEPIN(ICE_IOT_177));
    defparam ipInertedIOPad_ICE_IOT_177_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_177_preio (
            .PADOEN(N__59527),
            .PADOUT(N__59526),
            .PADIN(N__59525),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_141_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_141_iopad (
            .OE(N__59518),
            .DIN(N__59517),
            .DOUT(N__59516),
            .PACKAGEPIN(ICE_IOR_141));
    defparam ipInertedIOPad_ICE_IOR_141_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_141_preio (
            .PADOEN(N__59518),
            .PADOUT(N__59517),
            .PADIN(N__59516),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOB_80_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOB_80_iopad (
            .OE(N__59509),
            .DIN(N__59508),
            .DOUT(N__59507),
            .PACKAGEPIN(ICE_IOB_80));
    defparam ipInertedIOPad_ICE_IOB_80_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_80_preio (
            .PADOEN(N__59509),
            .PADOUT(N__59508),
            .PADIN(N__59507),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOB_102_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOB_102_iopad (
            .OE(N__59500),
            .DIN(N__59499),
            .DOUT(N__59498),
            .PACKAGEPIN(ICE_IOB_102));
    defparam ipInertedIOPad_ICE_IOB_102_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_102_preio (
            .PADOEN(N__59500),
            .PADOUT(N__59499),
            .PADIN(N__59498),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_GPMO_2_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_GPMO_2_iopad (
            .OE(N__59491),
            .DIN(N__59490),
            .DOUT(N__59489),
            .PACKAGEPIN(ICE_GPMO_2));
    defparam ipInertedIOPad_ICE_GPMO_2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_GPMO_2_preio (
            .PADOEN(N__59491),
            .PADOUT(N__59490),
            .PADIN(N__59489),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(ICE_GPMO_2),
            .DIN1());
    IO_PAD ipInertedIOPad_ICE_GPMI_0_iopad (
            .OE(N__59482),
            .DIN(N__59481),
            .DOUT(N__59480),
            .PACKAGEPIN(ICE_GPMI_0));
    defparam ipInertedIOPad_ICE_GPMI_0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_ICE_GPMI_0_preio (
            .PADOEN(N__59482),
            .PADOUT(N__59481),
            .PADIN(N__59480),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__56118),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_MISO_iopad (
            .OE(N__59473),
            .DIN(N__59472),
            .DOUT(N__59471),
            .PACKAGEPIN(IAC_MISO));
    defparam ipInertedIOPad_IAC_MISO_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_IAC_MISO_preio (
            .PADOEN(N__59473),
            .PADOUT(N__59472),
            .PADIN(N__59471),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(IAC_MISO),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_OSR0_iopad (
            .OE(N__59464),
            .DIN(N__59463),
            .DOUT(N__59462),
            .PACKAGEPIN(VAC_OSR0));
    defparam ipInertedIOPad_VAC_OSR0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_OSR0_preio (
            .PADOEN(N__59464),
            .PADOUT(N__59463),
            .PADIN(N__59462),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__32106),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_MOSI_iopad (
            .OE(N__59455),
            .DIN(N__59454),
            .DOUT(N__59453),
            .PACKAGEPIN(VAC_MOSI));
    defparam ipInertedIOPad_VAC_MOSI_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_MOSI_preio (
            .PADOEN(N__59455),
            .PADOUT(N__59454),
            .PADIN(N__59453),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_TEST_LED_iopad (
            .OE(N__59446),
            .DIN(N__59445),
            .DOUT(N__59444),
            .PACKAGEPIN(TEST_LED));
    defparam ipInertedIOPad_TEST_LED_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_TEST_LED_preio (
            .PADOEN(N__59446),
            .PADOUT(N__59445),
            .PADIN(N__59444),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__34677),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_148_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_148_iopad (
            .OE(N__59437),
            .DIN(N__59436),
            .DOUT(N__59435),
            .PACKAGEPIN(ICE_IOR_148));
    defparam ipInertedIOPad_ICE_IOR_148_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_148_preio (
            .PADOEN(N__59437),
            .PADOUT(N__59436),
            .PADIN(N__59435),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_STAT_COMM_iopad (
            .OE(N__59428),
            .DIN(N__59427),
            .DOUT(N__59426),
            .PACKAGEPIN(STAT_COMM));
    defparam ipInertedIOPad_STAT_COMM_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_STAT_COMM_preio (
            .PADOEN(N__59428),
            .PADOUT(N__59427),
            .PADIN(N__59426),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__19398),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_SYSCLK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_SYSCLK_iopad (
            .OE(N__59419),
            .DIN(N__59418),
            .DOUT(N__59417),
            .PACKAGEPIN(ICE_SYSCLK));
    defparam ipInertedIOPad_ICE_SYSCLK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_SYSCLK_preio (
            .PADOEN(N__59419),
            .PADOUT(N__59418),
            .PADIN(N__59417),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(ICE_SYSCLK),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_161_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_161_iopad (
            .OE(N__59410),
            .DIN(N__59409),
            .DOUT(N__59408),
            .PACKAGEPIN(ICE_IOR_161));
    defparam ipInertedIOPad_ICE_IOR_161_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_161_preio (
            .PADOEN(N__59410),
            .PADOUT(N__59409),
            .PADIN(N__59408),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOB_95_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOB_95_iopad (
            .OE(N__59401),
            .DIN(N__59400),
            .DOUT(N__59399),
            .PACKAGEPIN(ICE_IOB_95));
    defparam ipInertedIOPad_ICE_IOB_95_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_95_preio (
            .PADOEN(N__59401),
            .PADOUT(N__59400),
            .PADIN(N__59399),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_ICE_IOB_82_iopad (
            .OE(N__59392),
            .DIN(N__59391),
            .DOUT(N__59390),
            .PACKAGEPIN(ICE_IOB_82));
    defparam ipInertedIOPad_ICE_IOB_82_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_82_preio (
            .PADOEN(N__59392),
            .PADOUT(N__59391),
            .PADIN(N__59390),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_ICE_IOB_104_iopad (
            .OE(N__59383),
            .DIN(N__59382),
            .DOUT(N__59381),
            .PACKAGEPIN(ICE_IOB_104));
    defparam ipInertedIOPad_ICE_IOB_104_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_104_preio (
            .PADOEN(N__59383),
            .PADOUT(N__59382),
            .PADIN(N__59381),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_CLK_iopad (
            .OE(N__59374),
            .DIN(N__59373),
            .DOUT(N__59372),
            .PACKAGEPIN(IAC_CLK));
    defparam ipInertedIOPad_IAC_CLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_CLK_preio (
            .PADOEN(N__59374),
            .PADOUT(N__59373),
            .PADIN(N__59372),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__31125),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_CS_iopad (
            .OE(N__59365),
            .DIN(N__59364),
            .DOUT(N__59363),
            .PACKAGEPIN(DDS_CS));
    defparam ipInertedIOPad_DDS_CS_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_CS_preio (
            .PADOEN(N__59365),
            .PADOUT(N__59364),
            .PADIN(N__59363),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__41949),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SELIRNG0_iopad (
            .OE(N__59356),
            .DIN(N__59355),
            .DOUT(N__59354),
            .PACKAGEPIN(SELIRNG0));
    defparam ipInertedIOPad_SELIRNG0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_SELIRNG0_preio (
            .PADOEN(N__59356),
            .PADOUT(N__59355),
            .PADIN(N__59354),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__45738),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_RTD_SDI_iopad (
            .OE(N__59347),
            .DIN(N__59346),
            .DOUT(N__59345),
            .PACKAGEPIN(RTD_SDI));
    defparam ipInertedIOPad_RTD_SDI_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_RTD_SDI_preio (
            .PADOEN(N__59347),
            .PADOUT(N__59346),
            .PADIN(N__59345),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__19560),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_221_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_221_iopad (
            .OE(N__59338),
            .DIN(N__59337),
            .DOUT(N__59336),
            .PACKAGEPIN(ICE_IOT_221));
    defparam ipInertedIOPad_ICE_IOT_221_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_221_preio (
            .PADOEN(N__59338),
            .PADOUT(N__59337),
            .PADIN(N__59336),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_197_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_197_iopad (
            .OE(N__59329),
            .DIN(N__59328),
            .DOUT(N__59327),
            .PACKAGEPIN(ICE_IOT_197));
    defparam ipInertedIOPad_ICE_IOT_197_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_197_preio (
            .PADOEN(N__59329),
            .PADOUT(N__59328),
            .PADIN(N__59327),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_MCLK_iopad (
            .OE(N__59320),
            .DIN(N__59319),
            .DOUT(N__59318),
            .PACKAGEPIN(DDS_MCLK));
    defparam ipInertedIOPad_DDS_MCLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_MCLK_preio (
            .PADOEN(N__59320),
            .PADOUT(N__59319),
            .PADIN(N__59318),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__50691),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_RTD_SCLK_iopad (
            .OE(N__59311),
            .DIN(N__59310),
            .DOUT(N__59309),
            .PACKAGEPIN(RTD_SCLK));
    defparam ipInertedIOPad_RTD_SCLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_RTD_SCLK_preio (
            .PADOEN(N__59311),
            .PADOUT(N__59310),
            .PADIN(N__59309),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__19539),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_RTD_CS_iopad (
            .OE(N__59302),
            .DIN(N__59301),
            .DOUT(N__59300),
            .PACKAGEPIN(RTD_CS));
    defparam ipInertedIOPad_RTD_CS_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_RTD_CS_preio (
            .PADOEN(N__59302),
            .PADOUT(N__59301),
            .PADIN(N__59300),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__20322),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_137_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_137_iopad (
            .OE(N__59293),
            .DIN(N__59292),
            .DOUT(N__59291),
            .PACKAGEPIN(ICE_IOR_137));
    defparam ipInertedIOPad_ICE_IOR_137_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_137_preio (
            .PADOEN(N__59293),
            .PADOUT(N__59292),
            .PADIN(N__59291),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_OSR1_iopad (
            .OE(N__59284),
            .DIN(N__59283),
            .DOUT(N__59282),
            .PACKAGEPIN(IAC_OSR1));
    defparam ipInertedIOPad_IAC_OSR1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_OSR1_preio (
            .PADOEN(N__59284),
            .PADOUT(N__59283),
            .PADIN(N__59282),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__26100),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_FLT0_iopad (
            .OE(N__59275),
            .DIN(N__59274),
            .DOUT(N__59273),
            .PACKAGEPIN(VAC_FLT0));
    defparam ipInertedIOPad_VAC_FLT0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_FLT0_preio (
            .PADOEN(N__59275),
            .PADOUT(N__59274),
            .PADIN(N__59273),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__30822),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_144_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_144_iopad (
            .OE(N__59266),
            .DIN(N__59265),
            .DOUT(N__59264),
            .PACKAGEPIN(ICE_IOR_144));
    defparam ipInertedIOPad_ICE_IOR_144_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_144_preio (
            .PADOEN(N__59266),
            .PADOUT(N__59265),
            .PADIN(N__59264),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_128_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_128_iopad (
            .OE(N__59257),
            .DIN(N__59256),
            .DOUT(N__59255),
            .PACKAGEPIN(ICE_IOR_128));
    defparam ipInertedIOPad_ICE_IOR_128_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_128_preio (
            .PADOEN(N__59257),
            .PADOUT(N__59256),
            .PADIN(N__59255),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_GPMO_1_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_GPMO_1_iopad (
            .OE(N__59248),
            .DIN(N__59247),
            .DOUT(N__59246),
            .PACKAGEPIN(ICE_GPMO_1));
    defparam ipInertedIOPad_ICE_GPMO_1_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_GPMO_1_preio (
            .PADOEN(N__59248),
            .PADOUT(N__59247),
            .PADIN(N__59246),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_SCLK_iopad (
            .OE(N__59239),
            .DIN(N__59238),
            .DOUT(N__59237),
            .PACKAGEPIN(IAC_SCLK));
    defparam ipInertedIOPad_IAC_SCLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_SCLK_preio (
            .PADOEN(N__59239),
            .PADOUT(N__59238),
            .PADIN(N__59237),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__24786),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_EIS_SYNCCLK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_EIS_SYNCCLK_iopad (
            .OE(N__59230),
            .DIN(N__59229),
            .DOUT(N__59228),
            .PACKAGEPIN(EIS_SYNCCLK));
    defparam ipInertedIOPad_EIS_SYNCCLK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_EIS_SYNCCLK_preio (
            .PADOEN(N__59230),
            .PADOUT(N__59229),
            .PADIN(N__59228),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(EIS_SYNCCLK),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_139_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_139_iopad (
            .OE(N__59221),
            .DIN(N__59220),
            .DOUT(N__59219),
            .PACKAGEPIN(ICE_IOR_139));
    defparam ipInertedIOPad_ICE_IOR_139_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_139_preio (
            .PADOEN(N__59221),
            .PADOUT(N__59220),
            .PADIN(N__59219),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_4A_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_4A_iopad (
            .OE(N__59212),
            .DIN(N__59211),
            .DOUT(N__59210),
            .PACKAGEPIN(ICE_IOL_4A));
    defparam ipInertedIOPad_ICE_IOL_4A_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_4A_preio (
            .PADOEN(N__59212),
            .PADOUT(N__59211),
            .PADIN(N__59210),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VAC_SCLK_iopad (
            .OE(N__59203),
            .DIN(N__59202),
            .DOUT(N__59201),
            .PACKAGEPIN(VAC_SCLK));
    defparam ipInertedIOPad_VAC_SCLK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VAC_SCLK_preio (
            .PADOEN(N__59203),
            .PADOUT(N__59202),
            .PADIN(N__59201),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__21468),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_THERMOSTAT_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_THERMOSTAT_iopad (
            .OE(N__59194),
            .DIN(N__59193),
            .DOUT(N__59192),
            .PACKAGEPIN(THERMOSTAT));
    defparam ipInertedIOPad_THERMOSTAT_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_THERMOSTAT_preio (
            .PADOEN(N__59194),
            .PADOUT(N__59193),
            .PADIN(N__59192),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(THERMOSTAT),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_164_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_164_iopad (
            .OE(N__59185),
            .DIN(N__59184),
            .DOUT(N__59183),
            .PACKAGEPIN(ICE_IOR_164));
    defparam ipInertedIOPad_ICE_IOR_164_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_164_preio (
            .PADOEN(N__59185),
            .PADOUT(N__59184),
            .PADIN(N__59183),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_ICE_IOB_103_iopad (
            .OE(N__59176),
            .DIN(N__59175),
            .DOUT(N__59174),
            .PACKAGEPIN(ICE_IOB_103));
    defparam ipInertedIOPad_ICE_IOB_103_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_103_preio (
            .PADOEN(N__59176),
            .PADOUT(N__59175),
            .PADIN(N__59174),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_AMPV_POW_iopad (
            .OE(N__59167),
            .DIN(N__59166),
            .DOUT(N__59165),
            .PACKAGEPIN(AMPV_POW));
    defparam ipInertedIOPad_AMPV_POW_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_AMPV_POW_preio (
            .PADOEN(N__59167),
            .PADOUT(N__59166),
            .PADIN(N__59165),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__36015),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VDC_SDO_iopad (
            .OE(N__59158),
            .DIN(N__59157),
            .DOUT(N__59156),
            .PACKAGEPIN(VDC_SDO));
    defparam ipInertedIOPad_VDC_SDO_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VDC_SDO_preio (
            .PADOEN(N__59158),
            .PADOUT(N__59157),
            .PADIN(N__59156),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(VDC_SDO),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_174_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_174_iopad (
            .OE(N__59149),
            .DIN(N__59148),
            .DOUT(N__59147),
            .PACKAGEPIN(ICE_IOT_174));
    defparam ipInertedIOPad_ICE_IOT_174_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_174_preio (
            .PADOEN(N__59149),
            .PADOUT(N__59148),
            .PADIN(N__59147),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_140_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_140_iopad (
            .OE(N__59140),
            .DIN(N__59139),
            .DOUT(N__59138),
            .PACKAGEPIN(ICE_IOR_140));
    defparam ipInertedIOPad_ICE_IOR_140_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_140_preio (
            .PADOEN(N__59140),
            .PADOUT(N__59139),
            .PADIN(N__59138),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOB_96_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOB_96_iopad (
            .OE(N__59131),
            .DIN(N__59130),
            .DOUT(N__59129),
            .PACKAGEPIN(ICE_IOB_96));
    defparam ipInertedIOPad_ICE_IOB_96_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOB_96_preio (
            .PADOEN(N__59131),
            .PADOUT(N__59130),
            .PADIN(N__59129),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_CONT_SD_iopad (
            .OE(N__59122),
            .DIN(N__59121),
            .DOUT(N__59120),
            .PACKAGEPIN(CONT_SD));
    defparam ipInertedIOPad_CONT_SD_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_CONT_SD_preio (
            .PADOEN(N__59122),
            .PADOUT(N__59121),
            .PADIN(N__59120),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__44775),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_AC_ADC_SYNC_iopad (
            .OE(N__59113),
            .DIN(N__59112),
            .DOUT(N__59111),
            .PACKAGEPIN(AC_ADC_SYNC));
    defparam ipInertedIOPad_AC_ADC_SYNC_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_AC_ADC_SYNC_preio (
            .PADOEN(N__59113),
            .PADOUT(N__59112),
            .PADIN(N__59111),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__21903),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SELIRNG1_iopad (
            .OE(N__59104),
            .DIN(N__59103),
            .DOUT(N__59102),
            .PACKAGEPIN(SELIRNG1));
    defparam ipInertedIOPad_SELIRNG1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_SELIRNG1_preio (
            .PADOEN(N__59104),
            .PADOUT(N__59103),
            .PADIN(N__59102),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__36225),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOL_12B_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOL_12B_iopad (
            .OE(N__59095),
            .DIN(N__59094),
            .DOUT(N__59093),
            .PACKAGEPIN(ICE_IOL_12B));
    defparam ipInertedIOPad_ICE_IOL_12B_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOL_12B_preio (
            .PADOEN(N__59095),
            .PADOUT(N__59094),
            .PADIN(N__59093),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_160_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_160_iopad (
            .OE(N__59086),
            .DIN(N__59085),
            .DOUT(N__59084),
            .PACKAGEPIN(ICE_IOR_160));
    defparam ipInertedIOPad_ICE_IOR_160_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_160_preio (
            .PADOEN(N__59086),
            .PADOUT(N__59085),
            .PADIN(N__59084),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_136_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_136_iopad (
            .OE(N__59077),
            .DIN(N__59076),
            .DOUT(N__59075),
            .PACKAGEPIN(ICE_IOR_136));
    defparam ipInertedIOPad_ICE_IOR_136_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_136_preio (
            .PADOEN(N__59077),
            .PADOUT(N__59076),
            .PADIN(N__59075),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_MCLK1_iopad (
            .OE(N__59068),
            .DIN(N__59067),
            .DOUT(N__59066),
            .PACKAGEPIN(DDS_MCLK1));
    defparam ipInertedIOPad_DDS_MCLK1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_MCLK1_preio (
            .PADOEN(N__59068),
            .PADOUT(N__59067),
            .PADIN(N__59066),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__23751),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_198_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_198_iopad (
            .OE(N__59059),
            .DIN(N__59058),
            .DOUT(N__59057),
            .PACKAGEPIN(ICE_IOT_198));
    defparam ipInertedIOPad_ICE_IOT_198_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_198_preio (
            .PADOEN(N__59059),
            .PADOUT(N__59058),
            .PADIN(N__59057),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_173_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_173_iopad (
            .OE(N__59050),
            .DIN(N__59049),
            .DOUT(N__59048),
            .PACKAGEPIN(ICE_IOT_173));
    defparam ipInertedIOPad_ICE_IOT_173_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_173_preio (
            .PADOEN(N__59050),
            .PADOUT(N__59049),
            .PADIN(N__59048),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_DRDY_iopad (
            .OE(N__59041),
            .DIN(N__59040),
            .DOUT(N__59039),
            .PACKAGEPIN(IAC_DRDY));
    defparam ipInertedIOPad_IAC_DRDY_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_IAC_DRDY_preio (
            .PADOEN(N__59041),
            .PADOUT(N__59040),
            .PADIN(N__59039),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(IAC_DRDY),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOT_178_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOT_178_iopad (
            .OE(N__59032),
            .DIN(N__59031),
            .DOUT(N__59030),
            .PACKAGEPIN(ICE_IOT_178));
    defparam ipInertedIOPad_ICE_IOT_178_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOT_178_preio (
            .PADOEN(N__59032),
            .PADOUT(N__59031),
            .PADIN(N__59030),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_138_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_138_iopad (
            .OE(N__59023),
            .DIN(N__59022),
            .DOUT(N__59021),
            .PACKAGEPIN(ICE_IOR_138));
    defparam ipInertedIOPad_ICE_IOR_138_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_138_preio (
            .PADOEN(N__59023),
            .PADOUT(N__59022),
            .PADIN(N__59021),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_ICE_IOR_120_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_ICE_IOR_120_iopad (
            .OE(N__59014),
            .DIN(N__59013),
            .DOUT(N__59012),
            .PACKAGEPIN(ICE_IOR_120));
    defparam ipInertedIOPad_ICE_IOR_120_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_ICE_IOR_120_preio (
            .PADOEN(N__59014),
            .PADOUT(N__59013),
            .PADIN(N__59012),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_IAC_FLT0_iopad (
            .OE(N__59005),
            .DIN(N__59004),
            .DOUT(N__59003),
            .PACKAGEPIN(IAC_FLT0));
    defparam ipInertedIOPad_IAC_FLT0_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_IAC_FLT0_preio (
            .PADOEN(N__59005),
            .PADOUT(N__59004),
            .PADIN(N__59003),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__30546),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_DDS_SCK1_iopad (
            .OE(N__58996),
            .DIN(N__58995),
            .DOUT(N__58994),
            .PACKAGEPIN(DDS_SCK1));
    defparam ipInertedIOPad_DDS_SCK1_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DDS_SCK1_preio (
            .PADOEN(N__58996),
            .PADOUT(N__58995),
            .PADIN(N__58994),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__27189),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    SRMux I__14786 (
            .O(N__58977),
            .I(N__58974));
    LocalMux I__14785 (
            .O(N__58974),
            .I(N__58969));
    SRMux I__14784 (
            .O(N__58973),
            .I(N__58965));
    SRMux I__14783 (
            .O(N__58972),
            .I(N__58962));
    Span4Mux_h I__14782 (
            .O(N__58969),
            .I(N__58959));
    SRMux I__14781 (
            .O(N__58968),
            .I(N__58956));
    LocalMux I__14780 (
            .O(N__58965),
            .I(N__58953));
    LocalMux I__14779 (
            .O(N__58962),
            .I(N__58950));
    Span4Mux_h I__14778 (
            .O(N__58959),
            .I(N__58945));
    LocalMux I__14777 (
            .O(N__58956),
            .I(N__58945));
    Span4Mux_h I__14776 (
            .O(N__58953),
            .I(N__58942));
    Span4Mux_v I__14775 (
            .O(N__58950),
            .I(N__58939));
    Span4Mux_v I__14774 (
            .O(N__58945),
            .I(N__58934));
    Span4Mux_h I__14773 (
            .O(N__58942),
            .I(N__58934));
    Span4Mux_h I__14772 (
            .O(N__58939),
            .I(N__58931));
    Odrv4 I__14771 (
            .O(N__58934),
            .I(\ADC_VDC.genclk.n14894 ));
    Odrv4 I__14770 (
            .O(N__58931),
            .I(\ADC_VDC.genclk.n14894 ));
    SRMux I__14769 (
            .O(N__58926),
            .I(N__58923));
    LocalMux I__14768 (
            .O(N__58923),
            .I(N__58920));
    Span4Mux_v I__14767 (
            .O(N__58920),
            .I(N__58917));
    Odrv4 I__14766 (
            .O(N__58917),
            .I(\comm_spi.data_tx_7__N_835 ));
    InMux I__14765 (
            .O(N__58914),
            .I(N__58911));
    LocalMux I__14764 (
            .O(N__58911),
            .I(N__58907));
    InMux I__14763 (
            .O(N__58910),
            .I(N__58904));
    Span4Mux_v I__14762 (
            .O(N__58907),
            .I(N__58899));
    LocalMux I__14761 (
            .O(N__58904),
            .I(N__58899));
    Odrv4 I__14760 (
            .O(N__58899),
            .I(\comm_spi.n14827 ));
    InMux I__14759 (
            .O(N__58896),
            .I(N__58893));
    LocalMux I__14758 (
            .O(N__58893),
            .I(N__58888));
    InMux I__14757 (
            .O(N__58892),
            .I(N__58885));
    InMux I__14756 (
            .O(N__58891),
            .I(N__58882));
    Odrv4 I__14755 (
            .O(N__58888),
            .I(\comm_spi.n23110 ));
    LocalMux I__14754 (
            .O(N__58885),
            .I(\comm_spi.n23110 ));
    LocalMux I__14753 (
            .O(N__58882),
            .I(\comm_spi.n23110 ));
    InMux I__14752 (
            .O(N__58875),
            .I(N__58871));
    InMux I__14751 (
            .O(N__58874),
            .I(N__58868));
    LocalMux I__14750 (
            .O(N__58871),
            .I(N__58863));
    LocalMux I__14749 (
            .O(N__58868),
            .I(N__58863));
    Odrv12 I__14748 (
            .O(N__58863),
            .I(\comm_spi.n14801 ));
    InMux I__14747 (
            .O(N__58860),
            .I(N__58857));
    LocalMux I__14746 (
            .O(N__58857),
            .I(N__58853));
    InMux I__14745 (
            .O(N__58856),
            .I(N__58850));
    Span4Mux_v I__14744 (
            .O(N__58853),
            .I(N__58847));
    LocalMux I__14743 (
            .O(N__58850),
            .I(N__58844));
    Odrv4 I__14742 (
            .O(N__58847),
            .I(\comm_spi.n14826 ));
    Odrv12 I__14741 (
            .O(N__58844),
            .I(\comm_spi.n14826 ));
    SRMux I__14740 (
            .O(N__58839),
            .I(N__58836));
    LocalMux I__14739 (
            .O(N__58836),
            .I(N__58833));
    Odrv4 I__14738 (
            .O(N__58833),
            .I(\comm_spi.data_tx_7__N_812 ));
    SRMux I__14737 (
            .O(N__58830),
            .I(N__58827));
    LocalMux I__14736 (
            .O(N__58827),
            .I(N__58824));
    Span4Mux_v I__14735 (
            .O(N__58824),
            .I(N__58821));
    Odrv4 I__14734 (
            .O(N__58821),
            .I(\comm_spi.data_tx_7__N_832 ));
    InMux I__14733 (
            .O(N__58818),
            .I(N__58809));
    InMux I__14732 (
            .O(N__58817),
            .I(N__58809));
    InMux I__14731 (
            .O(N__58816),
            .I(N__58809));
    LocalMux I__14730 (
            .O(N__58809),
            .I(N__58806));
    Span4Mux_v I__14729 (
            .O(N__58806),
            .I(N__58803));
    Odrv4 I__14728 (
            .O(N__58803),
            .I(comm_tx_buf_1));
    InMux I__14727 (
            .O(N__58800),
            .I(N__58797));
    LocalMux I__14726 (
            .O(N__58797),
            .I(N__58793));
    InMux I__14725 (
            .O(N__58796),
            .I(N__58790));
    Span4Mux_v I__14724 (
            .O(N__58793),
            .I(N__58784));
    LocalMux I__14723 (
            .O(N__58790),
            .I(N__58784));
    InMux I__14722 (
            .O(N__58789),
            .I(N__58781));
    Odrv4 I__14721 (
            .O(N__58784),
            .I(\comm_spi.n23107 ));
    LocalMux I__14720 (
            .O(N__58781),
            .I(\comm_spi.n23107 ));
    SRMux I__14719 (
            .O(N__58776),
            .I(N__58770));
    SRMux I__14718 (
            .O(N__58775),
            .I(N__58767));
    SRMux I__14717 (
            .O(N__58774),
            .I(N__58759));
    IoInMux I__14716 (
            .O(N__58773),
            .I(N__58755));
    LocalMux I__14715 (
            .O(N__58770),
            .I(N__58738));
    LocalMux I__14714 (
            .O(N__58767),
            .I(N__58738));
    SRMux I__14713 (
            .O(N__58766),
            .I(N__58735));
    InMux I__14712 (
            .O(N__58765),
            .I(N__58732));
    SRMux I__14711 (
            .O(N__58764),
            .I(N__58729));
    SRMux I__14710 (
            .O(N__58763),
            .I(N__58725));
    SRMux I__14709 (
            .O(N__58762),
            .I(N__58722));
    LocalMux I__14708 (
            .O(N__58759),
            .I(N__58712));
    SRMux I__14707 (
            .O(N__58758),
            .I(N__58709));
    LocalMux I__14706 (
            .O(N__58755),
            .I(N__58699));
    CascadeMux I__14705 (
            .O(N__58754),
            .I(N__58696));
    CascadeMux I__14704 (
            .O(N__58753),
            .I(N__58692));
    CascadeMux I__14703 (
            .O(N__58752),
            .I(N__58688));
    CascadeMux I__14702 (
            .O(N__58751),
            .I(N__58684));
    CascadeMux I__14701 (
            .O(N__58750),
            .I(N__58680));
    CascadeMux I__14700 (
            .O(N__58749),
            .I(N__58676));
    CascadeMux I__14699 (
            .O(N__58748),
            .I(N__58672));
    CascadeMux I__14698 (
            .O(N__58747),
            .I(N__58668));
    CascadeMux I__14697 (
            .O(N__58746),
            .I(N__58665));
    CascadeMux I__14696 (
            .O(N__58745),
            .I(N__58661));
    CascadeMux I__14695 (
            .O(N__58744),
            .I(N__58657));
    CascadeMux I__14694 (
            .O(N__58743),
            .I(N__58653));
    Span4Mux_v I__14693 (
            .O(N__58738),
            .I(N__58644));
    LocalMux I__14692 (
            .O(N__58735),
            .I(N__58644));
    LocalMux I__14691 (
            .O(N__58732),
            .I(N__58644));
    LocalMux I__14690 (
            .O(N__58729),
            .I(N__58644));
    SRMux I__14689 (
            .O(N__58728),
            .I(N__58641));
    LocalMux I__14688 (
            .O(N__58725),
            .I(N__58636));
    LocalMux I__14687 (
            .O(N__58722),
            .I(N__58636));
    InMux I__14686 (
            .O(N__58721),
            .I(N__58633));
    SRMux I__14685 (
            .O(N__58720),
            .I(N__58630));
    SRMux I__14684 (
            .O(N__58719),
            .I(N__58627));
    CascadeMux I__14683 (
            .O(N__58718),
            .I(N__58623));
    CascadeMux I__14682 (
            .O(N__58717),
            .I(N__58619));
    CascadeMux I__14681 (
            .O(N__58716),
            .I(N__58615));
    CascadeMux I__14680 (
            .O(N__58715),
            .I(N__58611));
    Span4Mux_v I__14679 (
            .O(N__58712),
            .I(N__58608));
    LocalMux I__14678 (
            .O(N__58709),
            .I(N__58605));
    InMux I__14677 (
            .O(N__58708),
            .I(N__58598));
    InMux I__14676 (
            .O(N__58707),
            .I(N__58598));
    InMux I__14675 (
            .O(N__58706),
            .I(N__58598));
    InMux I__14674 (
            .O(N__58705),
            .I(N__58589));
    InMux I__14673 (
            .O(N__58704),
            .I(N__58589));
    InMux I__14672 (
            .O(N__58703),
            .I(N__58589));
    InMux I__14671 (
            .O(N__58702),
            .I(N__58589));
    Span4Mux_s2_v I__14670 (
            .O(N__58699),
            .I(N__58586));
    InMux I__14669 (
            .O(N__58696),
            .I(N__58571));
    InMux I__14668 (
            .O(N__58695),
            .I(N__58571));
    InMux I__14667 (
            .O(N__58692),
            .I(N__58571));
    InMux I__14666 (
            .O(N__58691),
            .I(N__58571));
    InMux I__14665 (
            .O(N__58688),
            .I(N__58571));
    InMux I__14664 (
            .O(N__58687),
            .I(N__58571));
    InMux I__14663 (
            .O(N__58684),
            .I(N__58571));
    InMux I__14662 (
            .O(N__58683),
            .I(N__58554));
    InMux I__14661 (
            .O(N__58680),
            .I(N__58554));
    InMux I__14660 (
            .O(N__58679),
            .I(N__58554));
    InMux I__14659 (
            .O(N__58676),
            .I(N__58554));
    InMux I__14658 (
            .O(N__58675),
            .I(N__58554));
    InMux I__14657 (
            .O(N__58672),
            .I(N__58554));
    InMux I__14656 (
            .O(N__58671),
            .I(N__58554));
    InMux I__14655 (
            .O(N__58668),
            .I(N__58554));
    InMux I__14654 (
            .O(N__58665),
            .I(N__58539));
    InMux I__14653 (
            .O(N__58664),
            .I(N__58539));
    InMux I__14652 (
            .O(N__58661),
            .I(N__58539));
    InMux I__14651 (
            .O(N__58660),
            .I(N__58539));
    InMux I__14650 (
            .O(N__58657),
            .I(N__58539));
    InMux I__14649 (
            .O(N__58656),
            .I(N__58539));
    InMux I__14648 (
            .O(N__58653),
            .I(N__58539));
    Span4Mux_v I__14647 (
            .O(N__58644),
            .I(N__58534));
    LocalMux I__14646 (
            .O(N__58641),
            .I(N__58534));
    Span4Mux_v I__14645 (
            .O(N__58636),
            .I(N__58525));
    LocalMux I__14644 (
            .O(N__58633),
            .I(N__58525));
    LocalMux I__14643 (
            .O(N__58630),
            .I(N__58525));
    LocalMux I__14642 (
            .O(N__58627),
            .I(N__58525));
    InMux I__14641 (
            .O(N__58626),
            .I(N__58508));
    InMux I__14640 (
            .O(N__58623),
            .I(N__58508));
    InMux I__14639 (
            .O(N__58622),
            .I(N__58508));
    InMux I__14638 (
            .O(N__58619),
            .I(N__58508));
    InMux I__14637 (
            .O(N__58618),
            .I(N__58508));
    InMux I__14636 (
            .O(N__58615),
            .I(N__58508));
    InMux I__14635 (
            .O(N__58614),
            .I(N__58508));
    InMux I__14634 (
            .O(N__58611),
            .I(N__58508));
    Span4Mux_v I__14633 (
            .O(N__58608),
            .I(N__58503));
    Span4Mux_h I__14632 (
            .O(N__58605),
            .I(N__58503));
    LocalMux I__14631 (
            .O(N__58598),
            .I(N__58498));
    LocalMux I__14630 (
            .O(N__58589),
            .I(N__58498));
    Sp12to4 I__14629 (
            .O(N__58586),
            .I(N__58495));
    LocalMux I__14628 (
            .O(N__58571),
            .I(N__58490));
    LocalMux I__14627 (
            .O(N__58554),
            .I(N__58490));
    LocalMux I__14626 (
            .O(N__58539),
            .I(N__58487));
    Span4Mux_v I__14625 (
            .O(N__58534),
            .I(N__58481));
    Span4Mux_v I__14624 (
            .O(N__58525),
            .I(N__58481));
    LocalMux I__14623 (
            .O(N__58508),
            .I(N__58478));
    Span4Mux_h I__14622 (
            .O(N__58503),
            .I(N__58475));
    Span4Mux_v I__14621 (
            .O(N__58498),
            .I(N__58472));
    Span12Mux_h I__14620 (
            .O(N__58495),
            .I(N__58469));
    Span4Mux_v I__14619 (
            .O(N__58490),
            .I(N__58466));
    Span4Mux_v I__14618 (
            .O(N__58487),
            .I(N__58463));
    SRMux I__14617 (
            .O(N__58486),
            .I(N__58460));
    Span4Mux_h I__14616 (
            .O(N__58481),
            .I(N__58455));
    Span4Mux_h I__14615 (
            .O(N__58478),
            .I(N__58455));
    Span4Mux_h I__14614 (
            .O(N__58475),
            .I(N__58450));
    Span4Mux_v I__14613 (
            .O(N__58472),
            .I(N__58450));
    Span12Mux_v I__14612 (
            .O(N__58469),
            .I(N__58441));
    Sp12to4 I__14611 (
            .O(N__58466),
            .I(N__58441));
    Sp12to4 I__14610 (
            .O(N__58463),
            .I(N__58441));
    LocalMux I__14609 (
            .O(N__58460),
            .I(N__58441));
    Span4Mux_h I__14608 (
            .O(N__58455),
            .I(N__58438));
    Odrv4 I__14607 (
            .O(N__58450),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__14606 (
            .O(N__58441),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__14605 (
            .O(N__58438),
            .I(CONSTANT_ONE_NET));
    InMux I__14604 (
            .O(N__58431),
            .I(N__58427));
    InMux I__14603 (
            .O(N__58430),
            .I(N__58424));
    LocalMux I__14602 (
            .O(N__58427),
            .I(N__58421));
    LocalMux I__14601 (
            .O(N__58424),
            .I(N__58418));
    Odrv4 I__14600 (
            .O(N__58421),
            .I(\comm_spi.n14800 ));
    Odrv4 I__14599 (
            .O(N__58418),
            .I(\comm_spi.n14800 ));
    ClkMux I__14598 (
            .O(N__58413),
            .I(N__58409));
    ClkMux I__14597 (
            .O(N__58412),
            .I(N__58403));
    LocalMux I__14596 (
            .O(N__58409),
            .I(N__58396));
    ClkMux I__14595 (
            .O(N__58408),
            .I(N__58393));
    ClkMux I__14594 (
            .O(N__58407),
            .I(N__58388));
    ClkMux I__14593 (
            .O(N__58406),
            .I(N__58385));
    LocalMux I__14592 (
            .O(N__58403),
            .I(N__58381));
    ClkMux I__14591 (
            .O(N__58402),
            .I(N__58378));
    ClkMux I__14590 (
            .O(N__58401),
            .I(N__58375));
    ClkMux I__14589 (
            .O(N__58400),
            .I(N__58372));
    ClkMux I__14588 (
            .O(N__58399),
            .I(N__58368));
    Span4Mux_v I__14587 (
            .O(N__58396),
            .I(N__58362));
    LocalMux I__14586 (
            .O(N__58393),
            .I(N__58362));
    ClkMux I__14585 (
            .O(N__58392),
            .I(N__58359));
    ClkMux I__14584 (
            .O(N__58391),
            .I(N__58353));
    LocalMux I__14583 (
            .O(N__58388),
            .I(N__58347));
    LocalMux I__14582 (
            .O(N__58385),
            .I(N__58347));
    ClkMux I__14581 (
            .O(N__58384),
            .I(N__58344));
    Span4Mux_v I__14580 (
            .O(N__58381),
            .I(N__58341));
    LocalMux I__14579 (
            .O(N__58378),
            .I(N__58338));
    LocalMux I__14578 (
            .O(N__58375),
            .I(N__58332));
    LocalMux I__14577 (
            .O(N__58372),
            .I(N__58332));
    ClkMux I__14576 (
            .O(N__58371),
            .I(N__58329));
    LocalMux I__14575 (
            .O(N__58368),
            .I(N__58325));
    ClkMux I__14574 (
            .O(N__58367),
            .I(N__58322));
    Span4Mux_v I__14573 (
            .O(N__58362),
            .I(N__58317));
    LocalMux I__14572 (
            .O(N__58359),
            .I(N__58317));
    ClkMux I__14571 (
            .O(N__58358),
            .I(N__58314));
    ClkMux I__14570 (
            .O(N__58357),
            .I(N__58311));
    ClkMux I__14569 (
            .O(N__58356),
            .I(N__58308));
    LocalMux I__14568 (
            .O(N__58353),
            .I(N__58304));
    ClkMux I__14567 (
            .O(N__58352),
            .I(N__58301));
    Span4Mux_v I__14566 (
            .O(N__58347),
            .I(N__58298));
    LocalMux I__14565 (
            .O(N__58344),
            .I(N__58295));
    Span4Mux_h I__14564 (
            .O(N__58341),
            .I(N__58290));
    Span4Mux_h I__14563 (
            .O(N__58338),
            .I(N__58290));
    ClkMux I__14562 (
            .O(N__58337),
            .I(N__58287));
    Span4Mux_v I__14561 (
            .O(N__58332),
            .I(N__58284));
    LocalMux I__14560 (
            .O(N__58329),
            .I(N__58281));
    ClkMux I__14559 (
            .O(N__58328),
            .I(N__58278));
    Span4Mux_h I__14558 (
            .O(N__58325),
            .I(N__58273));
    LocalMux I__14557 (
            .O(N__58322),
            .I(N__58273));
    Span4Mux_h I__14556 (
            .O(N__58317),
            .I(N__58270));
    LocalMux I__14555 (
            .O(N__58314),
            .I(N__58267));
    LocalMux I__14554 (
            .O(N__58311),
            .I(N__58264));
    LocalMux I__14553 (
            .O(N__58308),
            .I(N__58261));
    ClkMux I__14552 (
            .O(N__58307),
            .I(N__58258));
    Span4Mux_v I__14551 (
            .O(N__58304),
            .I(N__58252));
    LocalMux I__14550 (
            .O(N__58301),
            .I(N__58252));
    Span4Mux_h I__14549 (
            .O(N__58298),
            .I(N__58243));
    Span4Mux_h I__14548 (
            .O(N__58295),
            .I(N__58243));
    Span4Mux_v I__14547 (
            .O(N__58290),
            .I(N__58243));
    LocalMux I__14546 (
            .O(N__58287),
            .I(N__58243));
    Span4Mux_h I__14545 (
            .O(N__58284),
            .I(N__58236));
    Span4Mux_h I__14544 (
            .O(N__58281),
            .I(N__58236));
    LocalMux I__14543 (
            .O(N__58278),
            .I(N__58236));
    Span4Mux_h I__14542 (
            .O(N__58273),
            .I(N__58231));
    Span4Mux_v I__14541 (
            .O(N__58270),
            .I(N__58231));
    Span4Mux_h I__14540 (
            .O(N__58267),
            .I(N__58222));
    Span4Mux_v I__14539 (
            .O(N__58264),
            .I(N__58222));
    Span4Mux_v I__14538 (
            .O(N__58261),
            .I(N__58222));
    LocalMux I__14537 (
            .O(N__58258),
            .I(N__58222));
    ClkMux I__14536 (
            .O(N__58257),
            .I(N__58219));
    Span4Mux_v I__14535 (
            .O(N__58252),
            .I(N__58216));
    Span4Mux_v I__14534 (
            .O(N__58243),
            .I(N__58211));
    Span4Mux_h I__14533 (
            .O(N__58236),
            .I(N__58211));
    Span4Mux_v I__14532 (
            .O(N__58231),
            .I(N__58206));
    Span4Mux_h I__14531 (
            .O(N__58222),
            .I(N__58206));
    LocalMux I__14530 (
            .O(N__58219),
            .I(N__58203));
    Odrv4 I__14529 (
            .O(N__58216),
            .I(\comm_spi.iclk ));
    Odrv4 I__14528 (
            .O(N__58211),
            .I(\comm_spi.iclk ));
    Odrv4 I__14527 (
            .O(N__58206),
            .I(\comm_spi.iclk ));
    Odrv12 I__14526 (
            .O(N__58203),
            .I(\comm_spi.iclk ));
    InMux I__14525 (
            .O(N__58194),
            .I(N__58187));
    InMux I__14524 (
            .O(N__58193),
            .I(N__58187));
    InMux I__14523 (
            .O(N__58192),
            .I(N__58184));
    LocalMux I__14522 (
            .O(N__58187),
            .I(N__58181));
    LocalMux I__14521 (
            .O(N__58184),
            .I(N__58178));
    Span4Mux_v I__14520 (
            .O(N__58181),
            .I(N__58173));
    Span4Mux_v I__14519 (
            .O(N__58178),
            .I(N__58173));
    Sp12to4 I__14518 (
            .O(N__58173),
            .I(N__58170));
    Odrv12 I__14517 (
            .O(N__58170),
            .I(comm_tx_buf_0));
    CascadeMux I__14516 (
            .O(N__58167),
            .I(N__58153));
    CascadeMux I__14515 (
            .O(N__58166),
            .I(N__58150));
    SRMux I__14514 (
            .O(N__58165),
            .I(N__58146));
    InMux I__14513 (
            .O(N__58164),
            .I(N__58140));
    InMux I__14512 (
            .O(N__58163),
            .I(N__58140));
    CascadeMux I__14511 (
            .O(N__58162),
            .I(N__58136));
    CascadeMux I__14510 (
            .O(N__58161),
            .I(N__58133));
    CascadeMux I__14509 (
            .O(N__58160),
            .I(N__58128));
    InMux I__14508 (
            .O(N__58159),
            .I(N__58123));
    InMux I__14507 (
            .O(N__58158),
            .I(N__58117));
    InMux I__14506 (
            .O(N__58157),
            .I(N__58114));
    CascadeMux I__14505 (
            .O(N__58156),
            .I(N__58110));
    InMux I__14504 (
            .O(N__58153),
            .I(N__58101));
    InMux I__14503 (
            .O(N__58150),
            .I(N__58101));
    InMux I__14502 (
            .O(N__58149),
            .I(N__58101));
    LocalMux I__14501 (
            .O(N__58146),
            .I(N__58098));
    SRMux I__14500 (
            .O(N__58145),
            .I(N__58095));
    LocalMux I__14499 (
            .O(N__58140),
            .I(N__58092));
    InMux I__14498 (
            .O(N__58139),
            .I(N__58081));
    InMux I__14497 (
            .O(N__58136),
            .I(N__58081));
    InMux I__14496 (
            .O(N__58133),
            .I(N__58081));
    InMux I__14495 (
            .O(N__58132),
            .I(N__58081));
    InMux I__14494 (
            .O(N__58131),
            .I(N__58081));
    InMux I__14493 (
            .O(N__58128),
            .I(N__58074));
    InMux I__14492 (
            .O(N__58127),
            .I(N__58074));
    InMux I__14491 (
            .O(N__58126),
            .I(N__58074));
    LocalMux I__14490 (
            .O(N__58123),
            .I(N__58071));
    SRMux I__14489 (
            .O(N__58122),
            .I(N__58068));
    InMux I__14488 (
            .O(N__58121),
            .I(N__58060));
    InMux I__14487 (
            .O(N__58120),
            .I(N__58060));
    LocalMux I__14486 (
            .O(N__58117),
            .I(N__58055));
    LocalMux I__14485 (
            .O(N__58114),
            .I(N__58048));
    InMux I__14484 (
            .O(N__58113),
            .I(N__58045));
    InMux I__14483 (
            .O(N__58110),
            .I(N__58038));
    InMux I__14482 (
            .O(N__58109),
            .I(N__58038));
    InMux I__14481 (
            .O(N__58108),
            .I(N__58038));
    LocalMux I__14480 (
            .O(N__58101),
            .I(N__58035));
    Span4Mux_v I__14479 (
            .O(N__58098),
            .I(N__58030));
    LocalMux I__14478 (
            .O(N__58095),
            .I(N__58030));
    Span4Mux_h I__14477 (
            .O(N__58092),
            .I(N__58023));
    LocalMux I__14476 (
            .O(N__58081),
            .I(N__58023));
    LocalMux I__14475 (
            .O(N__58074),
            .I(N__58023));
    Span4Mux_v I__14474 (
            .O(N__58071),
            .I(N__58018));
    LocalMux I__14473 (
            .O(N__58068),
            .I(N__58018));
    InMux I__14472 (
            .O(N__58067),
            .I(N__58013));
    InMux I__14471 (
            .O(N__58066),
            .I(N__58013));
    InMux I__14470 (
            .O(N__58065),
            .I(N__58010));
    LocalMux I__14469 (
            .O(N__58060),
            .I(N__58007));
    InMux I__14468 (
            .O(N__58059),
            .I(N__58002));
    InMux I__14467 (
            .O(N__58058),
            .I(N__58002));
    Span4Mux_v I__14466 (
            .O(N__58055),
            .I(N__57999));
    InMux I__14465 (
            .O(N__58054),
            .I(N__57994));
    InMux I__14464 (
            .O(N__58053),
            .I(N__57994));
    InMux I__14463 (
            .O(N__58052),
            .I(N__57989));
    InMux I__14462 (
            .O(N__58051),
            .I(N__57989));
    Span4Mux_h I__14461 (
            .O(N__58048),
            .I(N__57982));
    LocalMux I__14460 (
            .O(N__58045),
            .I(N__57982));
    LocalMux I__14459 (
            .O(N__58038),
            .I(N__57979));
    Span4Mux_v I__14458 (
            .O(N__58035),
            .I(N__57976));
    Span4Mux_h I__14457 (
            .O(N__58030),
            .I(N__57973));
    Span4Mux_v I__14456 (
            .O(N__58023),
            .I(N__57970));
    Span4Mux_v I__14455 (
            .O(N__58018),
            .I(N__57967));
    LocalMux I__14454 (
            .O(N__58013),
            .I(N__57960));
    LocalMux I__14453 (
            .O(N__58010),
            .I(N__57960));
    Span12Mux_s10_v I__14452 (
            .O(N__58007),
            .I(N__57960));
    LocalMux I__14451 (
            .O(N__58002),
            .I(N__57957));
    Sp12to4 I__14450 (
            .O(N__57999),
            .I(N__57950));
    LocalMux I__14449 (
            .O(N__57994),
            .I(N__57950));
    LocalMux I__14448 (
            .O(N__57989),
            .I(N__57950));
    InMux I__14447 (
            .O(N__57988),
            .I(N__57945));
    InMux I__14446 (
            .O(N__57987),
            .I(N__57945));
    Span4Mux_h I__14445 (
            .O(N__57982),
            .I(N__57940));
    Span4Mux_v I__14444 (
            .O(N__57979),
            .I(N__57940));
    Span4Mux_h I__14443 (
            .O(N__57976),
            .I(N__57935));
    Span4Mux_v I__14442 (
            .O(N__57973),
            .I(N__57935));
    Span4Mux_v I__14441 (
            .O(N__57970),
            .I(N__57932));
    Span4Mux_v I__14440 (
            .O(N__57967),
            .I(N__57929));
    Span12Mux_v I__14439 (
            .O(N__57960),
            .I(N__57926));
    Span12Mux_h I__14438 (
            .O(N__57957),
            .I(N__57919));
    Span12Mux_s11_h I__14437 (
            .O(N__57950),
            .I(N__57919));
    LocalMux I__14436 (
            .O(N__57945),
            .I(N__57919));
    Span4Mux_v I__14435 (
            .O(N__57940),
            .I(N__57916));
    Odrv4 I__14434 (
            .O(N__57935),
            .I(comm_clear));
    Odrv4 I__14433 (
            .O(N__57932),
            .I(comm_clear));
    Odrv4 I__14432 (
            .O(N__57929),
            .I(comm_clear));
    Odrv12 I__14431 (
            .O(N__57926),
            .I(comm_clear));
    Odrv12 I__14430 (
            .O(N__57919),
            .I(comm_clear));
    Odrv4 I__14429 (
            .O(N__57916),
            .I(comm_clear));
    SRMux I__14428 (
            .O(N__57903),
            .I(N__57900));
    LocalMux I__14427 (
            .O(N__57900),
            .I(\comm_spi.data_tx_7__N_813 ));
    InMux I__14426 (
            .O(N__57897),
            .I(N__57893));
    InMux I__14425 (
            .O(N__57896),
            .I(N__57890));
    LocalMux I__14424 (
            .O(N__57893),
            .I(N__57887));
    LocalMux I__14423 (
            .O(N__57890),
            .I(\ADC_VDC.genclk.t0on_8 ));
    Odrv4 I__14422 (
            .O(N__57887),
            .I(\ADC_VDC.genclk.t0on_8 ));
    InMux I__14421 (
            .O(N__57882),
            .I(bfn_22_8_0_));
    CascadeMux I__14420 (
            .O(N__57879),
            .I(N__57875));
    InMux I__14419 (
            .O(N__57878),
            .I(N__57872));
    InMux I__14418 (
            .O(N__57875),
            .I(N__57869));
    LocalMux I__14417 (
            .O(N__57872),
            .I(N__57866));
    LocalMux I__14416 (
            .O(N__57869),
            .I(\ADC_VDC.genclk.t0on_9 ));
    Odrv4 I__14415 (
            .O(N__57866),
            .I(\ADC_VDC.genclk.t0on_9 ));
    InMux I__14414 (
            .O(N__57861),
            .I(\ADC_VDC.genclk.n19911 ));
    InMux I__14413 (
            .O(N__57858),
            .I(N__57855));
    LocalMux I__14412 (
            .O(N__57855),
            .I(N__57851));
    InMux I__14411 (
            .O(N__57854),
            .I(N__57848));
    Span4Mux_h I__14410 (
            .O(N__57851),
            .I(N__57845));
    LocalMux I__14409 (
            .O(N__57848),
            .I(\ADC_VDC.genclk.t0on_10 ));
    Odrv4 I__14408 (
            .O(N__57845),
            .I(\ADC_VDC.genclk.t0on_10 ));
    InMux I__14407 (
            .O(N__57840),
            .I(\ADC_VDC.genclk.n19912 ));
    CascadeMux I__14406 (
            .O(N__57837),
            .I(N__57833));
    InMux I__14405 (
            .O(N__57836),
            .I(N__57830));
    InMux I__14404 (
            .O(N__57833),
            .I(N__57827));
    LocalMux I__14403 (
            .O(N__57830),
            .I(N__57824));
    LocalMux I__14402 (
            .O(N__57827),
            .I(\ADC_VDC.genclk.t0on_11 ));
    Odrv4 I__14401 (
            .O(N__57824),
            .I(\ADC_VDC.genclk.t0on_11 ));
    InMux I__14400 (
            .O(N__57819),
            .I(\ADC_VDC.genclk.n19913 ));
    InMux I__14399 (
            .O(N__57816),
            .I(N__57813));
    LocalMux I__14398 (
            .O(N__57813),
            .I(N__57809));
    InMux I__14397 (
            .O(N__57812),
            .I(N__57806));
    Span4Mux_h I__14396 (
            .O(N__57809),
            .I(N__57803));
    LocalMux I__14395 (
            .O(N__57806),
            .I(\ADC_VDC.genclk.t0on_12 ));
    Odrv4 I__14394 (
            .O(N__57803),
            .I(\ADC_VDC.genclk.t0on_12 ));
    InMux I__14393 (
            .O(N__57798),
            .I(\ADC_VDC.genclk.n19914 ));
    CascadeMux I__14392 (
            .O(N__57795),
            .I(N__57791));
    InMux I__14391 (
            .O(N__57794),
            .I(N__57788));
    InMux I__14390 (
            .O(N__57791),
            .I(N__57785));
    LocalMux I__14389 (
            .O(N__57788),
            .I(N__57782));
    LocalMux I__14388 (
            .O(N__57785),
            .I(\ADC_VDC.genclk.t0on_13 ));
    Odrv4 I__14387 (
            .O(N__57782),
            .I(\ADC_VDC.genclk.t0on_13 ));
    InMux I__14386 (
            .O(N__57777),
            .I(\ADC_VDC.genclk.n19915 ));
    InMux I__14385 (
            .O(N__57774),
            .I(N__57770));
    InMux I__14384 (
            .O(N__57773),
            .I(N__57767));
    LocalMux I__14383 (
            .O(N__57770),
            .I(N__57764));
    LocalMux I__14382 (
            .O(N__57767),
            .I(\ADC_VDC.genclk.t0on_14 ));
    Odrv4 I__14381 (
            .O(N__57764),
            .I(\ADC_VDC.genclk.t0on_14 ));
    InMux I__14380 (
            .O(N__57759),
            .I(\ADC_VDC.genclk.n19916 ));
    InMux I__14379 (
            .O(N__57756),
            .I(\ADC_VDC.genclk.n19917 ));
    CascadeMux I__14378 (
            .O(N__57753),
            .I(N__57750));
    InMux I__14377 (
            .O(N__57750),
            .I(N__57746));
    InMux I__14376 (
            .O(N__57749),
            .I(N__57743));
    LocalMux I__14375 (
            .O(N__57746),
            .I(N__57740));
    LocalMux I__14374 (
            .O(N__57743),
            .I(\ADC_VDC.genclk.t0on_15 ));
    Odrv4 I__14373 (
            .O(N__57740),
            .I(\ADC_VDC.genclk.t0on_15 ));
    CEMux I__14372 (
            .O(N__57735),
            .I(N__57731));
    CEMux I__14371 (
            .O(N__57734),
            .I(N__57728));
    LocalMux I__14370 (
            .O(N__57731),
            .I(N__57725));
    LocalMux I__14369 (
            .O(N__57728),
            .I(N__57722));
    Span4Mux_h I__14368 (
            .O(N__57725),
            .I(N__57719));
    Odrv4 I__14367 (
            .O(N__57722),
            .I(\ADC_VDC.genclk.div_state_1__N_1432 ));
    Odrv4 I__14366 (
            .O(N__57719),
            .I(\ADC_VDC.genclk.div_state_1__N_1432 ));
    InMux I__14365 (
            .O(N__57714),
            .I(N__57710));
    InMux I__14364 (
            .O(N__57713),
            .I(N__57707));
    LocalMux I__14363 (
            .O(N__57710),
            .I(N__57704));
    LocalMux I__14362 (
            .O(N__57707),
            .I(\ADC_VDC.genclk.t0on_0 ));
    Odrv4 I__14361 (
            .O(N__57704),
            .I(\ADC_VDC.genclk.t0on_0 ));
    InMux I__14360 (
            .O(N__57699),
            .I(bfn_22_7_0_));
    InMux I__14359 (
            .O(N__57696),
            .I(N__57692));
    InMux I__14358 (
            .O(N__57695),
            .I(N__57689));
    LocalMux I__14357 (
            .O(N__57692),
            .I(N__57686));
    LocalMux I__14356 (
            .O(N__57689),
            .I(\ADC_VDC.genclk.t0on_1 ));
    Odrv4 I__14355 (
            .O(N__57686),
            .I(\ADC_VDC.genclk.t0on_1 ));
    InMux I__14354 (
            .O(N__57681),
            .I(\ADC_VDC.genclk.n19903 ));
    CascadeMux I__14353 (
            .O(N__57678),
            .I(N__57674));
    InMux I__14352 (
            .O(N__57677),
            .I(N__57671));
    InMux I__14351 (
            .O(N__57674),
            .I(N__57668));
    LocalMux I__14350 (
            .O(N__57671),
            .I(N__57665));
    LocalMux I__14349 (
            .O(N__57668),
            .I(\ADC_VDC.genclk.t0on_2 ));
    Odrv4 I__14348 (
            .O(N__57665),
            .I(\ADC_VDC.genclk.t0on_2 ));
    InMux I__14347 (
            .O(N__57660),
            .I(\ADC_VDC.genclk.n19904 ));
    InMux I__14346 (
            .O(N__57657),
            .I(N__57654));
    LocalMux I__14345 (
            .O(N__57654),
            .I(N__57650));
    InMux I__14344 (
            .O(N__57653),
            .I(N__57647));
    Span4Mux_h I__14343 (
            .O(N__57650),
            .I(N__57644));
    LocalMux I__14342 (
            .O(N__57647),
            .I(\ADC_VDC.genclk.t0on_3 ));
    Odrv4 I__14341 (
            .O(N__57644),
            .I(\ADC_VDC.genclk.t0on_3 ));
    InMux I__14340 (
            .O(N__57639),
            .I(\ADC_VDC.genclk.n19905 ));
    CascadeMux I__14339 (
            .O(N__57636),
            .I(N__57632));
    CascadeMux I__14338 (
            .O(N__57635),
            .I(N__57629));
    InMux I__14337 (
            .O(N__57632),
            .I(N__57626));
    InMux I__14336 (
            .O(N__57629),
            .I(N__57623));
    LocalMux I__14335 (
            .O(N__57626),
            .I(N__57620));
    LocalMux I__14334 (
            .O(N__57623),
            .I(\ADC_VDC.genclk.t0on_4 ));
    Odrv4 I__14333 (
            .O(N__57620),
            .I(\ADC_VDC.genclk.t0on_4 ));
    InMux I__14332 (
            .O(N__57615),
            .I(\ADC_VDC.genclk.n19906 ));
    CascadeMux I__14331 (
            .O(N__57612),
            .I(N__57609));
    InMux I__14330 (
            .O(N__57609),
            .I(N__57606));
    LocalMux I__14329 (
            .O(N__57606),
            .I(N__57602));
    InMux I__14328 (
            .O(N__57605),
            .I(N__57599));
    Span4Mux_v I__14327 (
            .O(N__57602),
            .I(N__57596));
    LocalMux I__14326 (
            .O(N__57599),
            .I(\ADC_VDC.genclk.t0on_5 ));
    Odrv4 I__14325 (
            .O(N__57596),
            .I(\ADC_VDC.genclk.t0on_5 ));
    InMux I__14324 (
            .O(N__57591),
            .I(\ADC_VDC.genclk.n19907 ));
    CascadeMux I__14323 (
            .O(N__57588),
            .I(N__57584));
    InMux I__14322 (
            .O(N__57587),
            .I(N__57581));
    InMux I__14321 (
            .O(N__57584),
            .I(N__57578));
    LocalMux I__14320 (
            .O(N__57581),
            .I(N__57575));
    LocalMux I__14319 (
            .O(N__57578),
            .I(\ADC_VDC.genclk.t0on_6 ));
    Odrv4 I__14318 (
            .O(N__57575),
            .I(\ADC_VDC.genclk.t0on_6 ));
    InMux I__14317 (
            .O(N__57570),
            .I(\ADC_VDC.genclk.n19908 ));
    CascadeMux I__14316 (
            .O(N__57567),
            .I(N__57564));
    InMux I__14315 (
            .O(N__57564),
            .I(N__57560));
    InMux I__14314 (
            .O(N__57563),
            .I(N__57557));
    LocalMux I__14313 (
            .O(N__57560),
            .I(N__57554));
    LocalMux I__14312 (
            .O(N__57557),
            .I(\ADC_VDC.genclk.t0on_7 ));
    Odrv4 I__14311 (
            .O(N__57554),
            .I(\ADC_VDC.genclk.t0on_7 ));
    InMux I__14310 (
            .O(N__57549),
            .I(\ADC_VDC.genclk.n19909 ));
    SRMux I__14309 (
            .O(N__57546),
            .I(N__57543));
    LocalMux I__14308 (
            .O(N__57543),
            .I(N__57540));
    Odrv12 I__14307 (
            .O(N__57540),
            .I(\comm_spi.data_tx_7__N_829 ));
    InMux I__14306 (
            .O(N__57537),
            .I(N__57532));
    InMux I__14305 (
            .O(N__57536),
            .I(N__57529));
    InMux I__14304 (
            .O(N__57535),
            .I(N__57526));
    LocalMux I__14303 (
            .O(N__57532),
            .I(\comm_spi.n23098 ));
    LocalMux I__14302 (
            .O(N__57529),
            .I(\comm_spi.n23098 ));
    LocalMux I__14301 (
            .O(N__57526),
            .I(\comm_spi.n23098 ));
    InMux I__14300 (
            .O(N__57519),
            .I(N__57516));
    LocalMux I__14299 (
            .O(N__57516),
            .I(N__57512));
    InMux I__14298 (
            .O(N__57515),
            .I(N__57509));
    Span4Mux_v I__14297 (
            .O(N__57512),
            .I(N__57506));
    LocalMux I__14296 (
            .O(N__57509),
            .I(N__57503));
    Span4Mux_h I__14295 (
            .O(N__57506),
            .I(N__57500));
    Span4Mux_v I__14294 (
            .O(N__57503),
            .I(N__57497));
    Odrv4 I__14293 (
            .O(N__57500),
            .I(\comm_spi.n14838 ));
    Odrv4 I__14292 (
            .O(N__57497),
            .I(\comm_spi.n14838 ));
    InMux I__14291 (
            .O(N__57492),
            .I(N__57488));
    InMux I__14290 (
            .O(N__57491),
            .I(N__57485));
    LocalMux I__14289 (
            .O(N__57488),
            .I(N__57482));
    LocalMux I__14288 (
            .O(N__57485),
            .I(N__57479));
    Odrv4 I__14287 (
            .O(N__57482),
            .I(\comm_spi.n14839 ));
    Odrv12 I__14286 (
            .O(N__57479),
            .I(\comm_spi.n14839 ));
    InMux I__14285 (
            .O(N__57474),
            .I(N__57471));
    LocalMux I__14284 (
            .O(N__57471),
            .I(N__57467));
    InMux I__14283 (
            .O(N__57470),
            .I(N__57464));
    Span4Mux_v I__14282 (
            .O(N__57467),
            .I(N__57459));
    LocalMux I__14281 (
            .O(N__57464),
            .I(N__57459));
    Span4Mux_h I__14280 (
            .O(N__57459),
            .I(N__57456));
    Span4Mux_h I__14279 (
            .O(N__57456),
            .I(N__57453));
    Odrv4 I__14278 (
            .O(N__57453),
            .I(\comm_spi.n14843 ));
    SRMux I__14277 (
            .O(N__57450),
            .I(N__57447));
    LocalMux I__14276 (
            .O(N__57447),
            .I(N__57444));
    Odrv4 I__14275 (
            .O(N__57444),
            .I(\comm_spi.data_tx_7__N_820 ));
    InMux I__14274 (
            .O(N__57441),
            .I(N__57438));
    LocalMux I__14273 (
            .O(N__57438),
            .I(N__57434));
    InMux I__14272 (
            .O(N__57437),
            .I(N__57431));
    Sp12to4 I__14271 (
            .O(N__57434),
            .I(N__57425));
    LocalMux I__14270 (
            .O(N__57431),
            .I(N__57425));
    InMux I__14269 (
            .O(N__57430),
            .I(N__57422));
    Odrv12 I__14268 (
            .O(N__57425),
            .I(\comm_spi.n23104 ));
    LocalMux I__14267 (
            .O(N__57422),
            .I(\comm_spi.n23104 ));
    InMux I__14266 (
            .O(N__57417),
            .I(N__57414));
    LocalMux I__14265 (
            .O(N__57414),
            .I(N__57410));
    InMux I__14264 (
            .O(N__57413),
            .I(N__57407));
    Sp12to4 I__14263 (
            .O(N__57410),
            .I(N__57402));
    LocalMux I__14262 (
            .O(N__57407),
            .I(N__57402));
    Odrv12 I__14261 (
            .O(N__57402),
            .I(\comm_spi.n14830 ));
    InMux I__14260 (
            .O(N__57399),
            .I(N__57396));
    LocalMux I__14259 (
            .O(N__57396),
            .I(N__57392));
    InMux I__14258 (
            .O(N__57395),
            .I(N__57389));
    Span4Mux_v I__14257 (
            .O(N__57392),
            .I(N__57386));
    LocalMux I__14256 (
            .O(N__57389),
            .I(N__57383));
    Odrv4 I__14255 (
            .O(N__57386),
            .I(\comm_spi.n14831 ));
    Odrv4 I__14254 (
            .O(N__57383),
            .I(\comm_spi.n14831 ));
    InMux I__14253 (
            .O(N__57378),
            .I(N__57375));
    LocalMux I__14252 (
            .O(N__57375),
            .I(N__57372));
    Span4Mux_h I__14251 (
            .O(N__57372),
            .I(N__57368));
    InMux I__14250 (
            .O(N__57371),
            .I(N__57365));
    Span4Mux_v I__14249 (
            .O(N__57368),
            .I(N__57362));
    LocalMux I__14248 (
            .O(N__57365),
            .I(N__57359));
    Odrv4 I__14247 (
            .O(N__57362),
            .I(\comm_spi.n14835 ));
    Odrv12 I__14246 (
            .O(N__57359),
            .I(\comm_spi.n14835 ));
    SRMux I__14245 (
            .O(N__57354),
            .I(N__57351));
    LocalMux I__14244 (
            .O(N__57351),
            .I(N__57348));
    Span4Mux_h I__14243 (
            .O(N__57348),
            .I(N__57345));
    Odrv4 I__14242 (
            .O(N__57345),
            .I(\comm_spi.data_tx_7__N_826 ));
    InMux I__14241 (
            .O(N__57342),
            .I(N__57339));
    LocalMux I__14240 (
            .O(N__57339),
            .I(buf_data_iac_13));
    InMux I__14239 (
            .O(N__57336),
            .I(N__57333));
    LocalMux I__14238 (
            .O(N__57333),
            .I(N__57330));
    Span12Mux_h I__14237 (
            .O(N__57330),
            .I(N__57327));
    Odrv12 I__14236 (
            .O(N__57327),
            .I(n21456));
    InMux I__14235 (
            .O(N__57324),
            .I(N__57321));
    LocalMux I__14234 (
            .O(N__57321),
            .I(buf_data_iac_12));
    InMux I__14233 (
            .O(N__57318),
            .I(N__57315));
    LocalMux I__14232 (
            .O(N__57315),
            .I(N__57312));
    Span4Mux_h I__14231 (
            .O(N__57312),
            .I(N__57309));
    Span4Mux_h I__14230 (
            .O(N__57309),
            .I(N__57306));
    Span4Mux_h I__14229 (
            .O(N__57306),
            .I(N__57303));
    Odrv4 I__14228 (
            .O(N__57303),
            .I(n21447));
    InMux I__14227 (
            .O(N__57300),
            .I(N__57297));
    LocalMux I__14226 (
            .O(N__57297),
            .I(N__57294));
    Odrv4 I__14225 (
            .O(N__57294),
            .I(buf_data_iac_9));
    InMux I__14224 (
            .O(N__57291),
            .I(N__57288));
    LocalMux I__14223 (
            .O(N__57288),
            .I(N__57285));
    Span4Mux_h I__14222 (
            .O(N__57285),
            .I(N__57282));
    Odrv4 I__14221 (
            .O(N__57282),
            .I(n21512));
    InMux I__14220 (
            .O(N__57279),
            .I(N__57276));
    LocalMux I__14219 (
            .O(N__57276),
            .I(buf_data_iac_11));
    CascadeMux I__14218 (
            .O(N__57273),
            .I(N__57254));
    InMux I__14217 (
            .O(N__57272),
            .I(N__57246));
    InMux I__14216 (
            .O(N__57271),
            .I(N__57243));
    InMux I__14215 (
            .O(N__57270),
            .I(N__57240));
    InMux I__14214 (
            .O(N__57269),
            .I(N__57233));
    InMux I__14213 (
            .O(N__57268),
            .I(N__57233));
    InMux I__14212 (
            .O(N__57267),
            .I(N__57230));
    InMux I__14211 (
            .O(N__57266),
            .I(N__57227));
    InMux I__14210 (
            .O(N__57265),
            .I(N__57224));
    InMux I__14209 (
            .O(N__57264),
            .I(N__57221));
    InMux I__14208 (
            .O(N__57263),
            .I(N__57218));
    CascadeMux I__14207 (
            .O(N__57262),
            .I(N__57214));
    CascadeMux I__14206 (
            .O(N__57261),
            .I(N__57199));
    InMux I__14205 (
            .O(N__57260),
            .I(N__57191));
    CascadeMux I__14204 (
            .O(N__57259),
            .I(N__57188));
    CascadeMux I__14203 (
            .O(N__57258),
            .I(N__57181));
    InMux I__14202 (
            .O(N__57257),
            .I(N__57170));
    InMux I__14201 (
            .O(N__57254),
            .I(N__57170));
    InMux I__14200 (
            .O(N__57253),
            .I(N__57170));
    InMux I__14199 (
            .O(N__57252),
            .I(N__57170));
    InMux I__14198 (
            .O(N__57251),
            .I(N__57167));
    InMux I__14197 (
            .O(N__57250),
            .I(N__57164));
    CascadeMux I__14196 (
            .O(N__57249),
            .I(N__57159));
    LocalMux I__14195 (
            .O(N__57246),
            .I(N__57152));
    LocalMux I__14194 (
            .O(N__57243),
            .I(N__57152));
    LocalMux I__14193 (
            .O(N__57240),
            .I(N__57152));
    InMux I__14192 (
            .O(N__57239),
            .I(N__57143));
    InMux I__14191 (
            .O(N__57238),
            .I(N__57140));
    LocalMux I__14190 (
            .O(N__57233),
            .I(N__57137));
    LocalMux I__14189 (
            .O(N__57230),
            .I(N__57122));
    LocalMux I__14188 (
            .O(N__57227),
            .I(N__57122));
    LocalMux I__14187 (
            .O(N__57224),
            .I(N__57115));
    LocalMux I__14186 (
            .O(N__57221),
            .I(N__57115));
    LocalMux I__14185 (
            .O(N__57218),
            .I(N__57115));
    CascadeMux I__14184 (
            .O(N__57217),
            .I(N__57106));
    InMux I__14183 (
            .O(N__57214),
            .I(N__57102));
    InMux I__14182 (
            .O(N__57213),
            .I(N__57094));
    InMux I__14181 (
            .O(N__57212),
            .I(N__57088));
    InMux I__14180 (
            .O(N__57211),
            .I(N__57083));
    InMux I__14179 (
            .O(N__57210),
            .I(N__57083));
    CascadeMux I__14178 (
            .O(N__57209),
            .I(N__57080));
    InMux I__14177 (
            .O(N__57208),
            .I(N__57077));
    InMux I__14176 (
            .O(N__57207),
            .I(N__57072));
    InMux I__14175 (
            .O(N__57206),
            .I(N__57072));
    InMux I__14174 (
            .O(N__57205),
            .I(N__57067));
    InMux I__14173 (
            .O(N__57204),
            .I(N__57067));
    InMux I__14172 (
            .O(N__57203),
            .I(N__57062));
    InMux I__14171 (
            .O(N__57202),
            .I(N__57062));
    InMux I__14170 (
            .O(N__57199),
            .I(N__57059));
    InMux I__14169 (
            .O(N__57198),
            .I(N__57052));
    InMux I__14168 (
            .O(N__57197),
            .I(N__57052));
    InMux I__14167 (
            .O(N__57196),
            .I(N__57052));
    InMux I__14166 (
            .O(N__57195),
            .I(N__57049));
    InMux I__14165 (
            .O(N__57194),
            .I(N__57046));
    LocalMux I__14164 (
            .O(N__57191),
            .I(N__57043));
    InMux I__14163 (
            .O(N__57188),
            .I(N__57038));
    InMux I__14162 (
            .O(N__57187),
            .I(N__57038));
    InMux I__14161 (
            .O(N__57186),
            .I(N__57035));
    InMux I__14160 (
            .O(N__57185),
            .I(N__57032));
    InMux I__14159 (
            .O(N__57184),
            .I(N__57029));
    InMux I__14158 (
            .O(N__57181),
            .I(N__57018));
    InMux I__14157 (
            .O(N__57180),
            .I(N__57018));
    InMux I__14156 (
            .O(N__57179),
            .I(N__57015));
    LocalMux I__14155 (
            .O(N__57170),
            .I(N__57012));
    LocalMux I__14154 (
            .O(N__57167),
            .I(N__57007));
    LocalMux I__14153 (
            .O(N__57164),
            .I(N__57007));
    InMux I__14152 (
            .O(N__57163),
            .I(N__57004));
    InMux I__14151 (
            .O(N__57162),
            .I(N__56999));
    InMux I__14150 (
            .O(N__57159),
            .I(N__56999));
    Span4Mux_v I__14149 (
            .O(N__57152),
            .I(N__56996));
    InMux I__14148 (
            .O(N__57151),
            .I(N__56993));
    InMux I__14147 (
            .O(N__57150),
            .I(N__56986));
    InMux I__14146 (
            .O(N__57149),
            .I(N__56986));
    InMux I__14145 (
            .O(N__57148),
            .I(N__56986));
    InMux I__14144 (
            .O(N__57147),
            .I(N__56983));
    InMux I__14143 (
            .O(N__57146),
            .I(N__56980));
    LocalMux I__14142 (
            .O(N__57143),
            .I(N__56975));
    LocalMux I__14141 (
            .O(N__57140),
            .I(N__56975));
    Span4Mux_h I__14140 (
            .O(N__57137),
            .I(N__56972));
    InMux I__14139 (
            .O(N__57136),
            .I(N__56961));
    InMux I__14138 (
            .O(N__57135),
            .I(N__56961));
    InMux I__14137 (
            .O(N__57134),
            .I(N__56961));
    InMux I__14136 (
            .O(N__57133),
            .I(N__56961));
    InMux I__14135 (
            .O(N__57132),
            .I(N__56961));
    InMux I__14134 (
            .O(N__57131),
            .I(N__56954));
    InMux I__14133 (
            .O(N__57130),
            .I(N__56949));
    InMux I__14132 (
            .O(N__57129),
            .I(N__56949));
    InMux I__14131 (
            .O(N__57128),
            .I(N__56946));
    InMux I__14130 (
            .O(N__57127),
            .I(N__56943));
    Span4Mux_v I__14129 (
            .O(N__57122),
            .I(N__56938));
    Span4Mux_v I__14128 (
            .O(N__57115),
            .I(N__56938));
    InMux I__14127 (
            .O(N__57114),
            .I(N__56934));
    InMux I__14126 (
            .O(N__57113),
            .I(N__56931));
    InMux I__14125 (
            .O(N__57112),
            .I(N__56928));
    InMux I__14124 (
            .O(N__57111),
            .I(N__56925));
    InMux I__14123 (
            .O(N__57110),
            .I(N__56918));
    InMux I__14122 (
            .O(N__57109),
            .I(N__56918));
    InMux I__14121 (
            .O(N__57106),
            .I(N__56918));
    InMux I__14120 (
            .O(N__57105),
            .I(N__56915));
    LocalMux I__14119 (
            .O(N__57102),
            .I(N__56910));
    InMux I__14118 (
            .O(N__57101),
            .I(N__56901));
    InMux I__14117 (
            .O(N__57100),
            .I(N__56901));
    InMux I__14116 (
            .O(N__57099),
            .I(N__56901));
    InMux I__14115 (
            .O(N__57098),
            .I(N__56901));
    InMux I__14114 (
            .O(N__57097),
            .I(N__56895));
    LocalMux I__14113 (
            .O(N__57094),
            .I(N__56892));
    InMux I__14112 (
            .O(N__57093),
            .I(N__56889));
    InMux I__14111 (
            .O(N__57092),
            .I(N__56884));
    InMux I__14110 (
            .O(N__57091),
            .I(N__56884));
    LocalMux I__14109 (
            .O(N__57088),
            .I(N__56881));
    LocalMux I__14108 (
            .O(N__57083),
            .I(N__56878));
    InMux I__14107 (
            .O(N__57080),
            .I(N__56875));
    LocalMux I__14106 (
            .O(N__57077),
            .I(N__56870));
    LocalMux I__14105 (
            .O(N__57072),
            .I(N__56856));
    LocalMux I__14104 (
            .O(N__57067),
            .I(N__56856));
    LocalMux I__14103 (
            .O(N__57062),
            .I(N__56856));
    LocalMux I__14102 (
            .O(N__57059),
            .I(N__56856));
    LocalMux I__14101 (
            .O(N__57052),
            .I(N__56853));
    LocalMux I__14100 (
            .O(N__57049),
            .I(N__56848));
    LocalMux I__14099 (
            .O(N__57046),
            .I(N__56848));
    Span4Mux_h I__14098 (
            .O(N__57043),
            .I(N__56843));
    LocalMux I__14097 (
            .O(N__57038),
            .I(N__56843));
    LocalMux I__14096 (
            .O(N__57035),
            .I(N__56836));
    LocalMux I__14095 (
            .O(N__57032),
            .I(N__56836));
    LocalMux I__14094 (
            .O(N__57029),
            .I(N__56836));
    InMux I__14093 (
            .O(N__57028),
            .I(N__56827));
    InMux I__14092 (
            .O(N__57027),
            .I(N__56827));
    InMux I__14091 (
            .O(N__57026),
            .I(N__56827));
    InMux I__14090 (
            .O(N__57025),
            .I(N__56827));
    InMux I__14089 (
            .O(N__57024),
            .I(N__56822));
    InMux I__14088 (
            .O(N__57023),
            .I(N__56822));
    LocalMux I__14087 (
            .O(N__57018),
            .I(N__56807));
    LocalMux I__14086 (
            .O(N__57015),
            .I(N__56807));
    Span4Mux_v I__14085 (
            .O(N__57012),
            .I(N__56807));
    Span4Mux_v I__14084 (
            .O(N__57007),
            .I(N__56807));
    LocalMux I__14083 (
            .O(N__57004),
            .I(N__56807));
    LocalMux I__14082 (
            .O(N__56999),
            .I(N__56807));
    Span4Mux_v I__14081 (
            .O(N__56996),
            .I(N__56807));
    LocalMux I__14080 (
            .O(N__56993),
            .I(N__56802));
    LocalMux I__14079 (
            .O(N__56986),
            .I(N__56802));
    LocalMux I__14078 (
            .O(N__56983),
            .I(N__56791));
    LocalMux I__14077 (
            .O(N__56980),
            .I(N__56791));
    Span4Mux_v I__14076 (
            .O(N__56975),
            .I(N__56791));
    Span4Mux_h I__14075 (
            .O(N__56972),
            .I(N__56791));
    LocalMux I__14074 (
            .O(N__56961),
            .I(N__56791));
    CascadeMux I__14073 (
            .O(N__56960),
            .I(N__56788));
    CascadeMux I__14072 (
            .O(N__56959),
            .I(N__56784));
    InMux I__14071 (
            .O(N__56958),
            .I(N__56778));
    InMux I__14070 (
            .O(N__56957),
            .I(N__56778));
    LocalMux I__14069 (
            .O(N__56954),
            .I(N__56767));
    LocalMux I__14068 (
            .O(N__56949),
            .I(N__56767));
    LocalMux I__14067 (
            .O(N__56946),
            .I(N__56767));
    LocalMux I__14066 (
            .O(N__56943),
            .I(N__56767));
    Sp12to4 I__14065 (
            .O(N__56938),
            .I(N__56767));
    InMux I__14064 (
            .O(N__56937),
            .I(N__56764));
    LocalMux I__14063 (
            .O(N__56934),
            .I(N__56753));
    LocalMux I__14062 (
            .O(N__56931),
            .I(N__56753));
    LocalMux I__14061 (
            .O(N__56928),
            .I(N__56753));
    LocalMux I__14060 (
            .O(N__56925),
            .I(N__56753));
    LocalMux I__14059 (
            .O(N__56918),
            .I(N__56753));
    LocalMux I__14058 (
            .O(N__56915),
            .I(N__56748));
    InMux I__14057 (
            .O(N__56914),
            .I(N__56743));
    InMux I__14056 (
            .O(N__56913),
            .I(N__56743));
    Span4Mux_v I__14055 (
            .O(N__56910),
            .I(N__56738));
    LocalMux I__14054 (
            .O(N__56901),
            .I(N__56738));
    InMux I__14053 (
            .O(N__56900),
            .I(N__56731));
    InMux I__14052 (
            .O(N__56899),
            .I(N__56731));
    InMux I__14051 (
            .O(N__56898),
            .I(N__56731));
    LocalMux I__14050 (
            .O(N__56895),
            .I(N__56728));
    Span4Mux_v I__14049 (
            .O(N__56892),
            .I(N__56723));
    LocalMux I__14048 (
            .O(N__56889),
            .I(N__56723));
    LocalMux I__14047 (
            .O(N__56884),
            .I(N__56720));
    Span4Mux_v I__14046 (
            .O(N__56881),
            .I(N__56713));
    Span4Mux_h I__14045 (
            .O(N__56878),
            .I(N__56713));
    LocalMux I__14044 (
            .O(N__56875),
            .I(N__56713));
    InMux I__14043 (
            .O(N__56874),
            .I(N__56710));
    InMux I__14042 (
            .O(N__56873),
            .I(N__56707));
    Span4Mux_v I__14041 (
            .O(N__56870),
            .I(N__56704));
    InMux I__14040 (
            .O(N__56869),
            .I(N__56697));
    InMux I__14039 (
            .O(N__56868),
            .I(N__56697));
    InMux I__14038 (
            .O(N__56867),
            .I(N__56697));
    InMux I__14037 (
            .O(N__56866),
            .I(N__56692));
    InMux I__14036 (
            .O(N__56865),
            .I(N__56692));
    Span4Mux_v I__14035 (
            .O(N__56856),
            .I(N__56687));
    Span4Mux_v I__14034 (
            .O(N__56853),
            .I(N__56687));
    Span4Mux_h I__14033 (
            .O(N__56848),
            .I(N__56680));
    Span4Mux_h I__14032 (
            .O(N__56843),
            .I(N__56680));
    Span4Mux_h I__14031 (
            .O(N__56836),
            .I(N__56680));
    LocalMux I__14030 (
            .O(N__56827),
            .I(N__56669));
    LocalMux I__14029 (
            .O(N__56822),
            .I(N__56669));
    Span4Mux_h I__14028 (
            .O(N__56807),
            .I(N__56669));
    Span4Mux_h I__14027 (
            .O(N__56802),
            .I(N__56669));
    Span4Mux_v I__14026 (
            .O(N__56791),
            .I(N__56669));
    InMux I__14025 (
            .O(N__56788),
            .I(N__56660));
    InMux I__14024 (
            .O(N__56787),
            .I(N__56660));
    InMux I__14023 (
            .O(N__56784),
            .I(N__56660));
    InMux I__14022 (
            .O(N__56783),
            .I(N__56660));
    LocalMux I__14021 (
            .O(N__56778),
            .I(N__56655));
    Span12Mux_h I__14020 (
            .O(N__56767),
            .I(N__56655));
    LocalMux I__14019 (
            .O(N__56764),
            .I(N__56650));
    Span12Mux_v I__14018 (
            .O(N__56753),
            .I(N__56650));
    InMux I__14017 (
            .O(N__56752),
            .I(N__56645));
    InMux I__14016 (
            .O(N__56751),
            .I(N__56645));
    Span4Mux_v I__14015 (
            .O(N__56748),
            .I(N__56628));
    LocalMux I__14014 (
            .O(N__56743),
            .I(N__56628));
    Span4Mux_h I__14013 (
            .O(N__56738),
            .I(N__56628));
    LocalMux I__14012 (
            .O(N__56731),
            .I(N__56628));
    Span4Mux_v I__14011 (
            .O(N__56728),
            .I(N__56628));
    Span4Mux_h I__14010 (
            .O(N__56723),
            .I(N__56628));
    Span4Mux_h I__14009 (
            .O(N__56720),
            .I(N__56628));
    Span4Mux_h I__14008 (
            .O(N__56713),
            .I(N__56628));
    LocalMux I__14007 (
            .O(N__56710),
            .I(comm_cmd_0));
    LocalMux I__14006 (
            .O(N__56707),
            .I(comm_cmd_0));
    Odrv4 I__14005 (
            .O(N__56704),
            .I(comm_cmd_0));
    LocalMux I__14004 (
            .O(N__56697),
            .I(comm_cmd_0));
    LocalMux I__14003 (
            .O(N__56692),
            .I(comm_cmd_0));
    Odrv4 I__14002 (
            .O(N__56687),
            .I(comm_cmd_0));
    Odrv4 I__14001 (
            .O(N__56680),
            .I(comm_cmd_0));
    Odrv4 I__14000 (
            .O(N__56669),
            .I(comm_cmd_0));
    LocalMux I__13999 (
            .O(N__56660),
            .I(comm_cmd_0));
    Odrv12 I__13998 (
            .O(N__56655),
            .I(comm_cmd_0));
    Odrv12 I__13997 (
            .O(N__56650),
            .I(comm_cmd_0));
    LocalMux I__13996 (
            .O(N__56645),
            .I(comm_cmd_0));
    Odrv4 I__13995 (
            .O(N__56628),
            .I(comm_cmd_0));
    InMux I__13994 (
            .O(N__56601),
            .I(N__56598));
    LocalMux I__13993 (
            .O(N__56598),
            .I(N__56595));
    Span4Mux_v I__13992 (
            .O(N__56595),
            .I(N__56592));
    Span4Mux_h I__13991 (
            .O(N__56592),
            .I(N__56589));
    Odrv4 I__13990 (
            .O(N__56589),
            .I(n21434));
    InMux I__13989 (
            .O(N__56586),
            .I(N__56583));
    LocalMux I__13988 (
            .O(N__56583),
            .I(N__56579));
    InMux I__13987 (
            .O(N__56582),
            .I(N__56575));
    Span12Mux_s11_v I__13986 (
            .O(N__56579),
            .I(N__56568));
    InMux I__13985 (
            .O(N__56578),
            .I(N__56565));
    LocalMux I__13984 (
            .O(N__56575),
            .I(N__56562));
    InMux I__13983 (
            .O(N__56574),
            .I(N__56557));
    InMux I__13982 (
            .O(N__56573),
            .I(N__56557));
    InMux I__13981 (
            .O(N__56572),
            .I(N__56552));
    InMux I__13980 (
            .O(N__56571),
            .I(N__56552));
    Odrv12 I__13979 (
            .O(N__56568),
            .I(\ADC_VDC.genclk.div_state_1 ));
    LocalMux I__13978 (
            .O(N__56565),
            .I(\ADC_VDC.genclk.div_state_1 ));
    Odrv4 I__13977 (
            .O(N__56562),
            .I(\ADC_VDC.genclk.div_state_1 ));
    LocalMux I__13976 (
            .O(N__56557),
            .I(\ADC_VDC.genclk.div_state_1 ));
    LocalMux I__13975 (
            .O(N__56552),
            .I(\ADC_VDC.genclk.div_state_1 ));
    CascadeMux I__13974 (
            .O(N__56541),
            .I(N__56538));
    InMux I__13973 (
            .O(N__56538),
            .I(N__56534));
    InMux I__13972 (
            .O(N__56537),
            .I(N__56531));
    LocalMux I__13971 (
            .O(N__56534),
            .I(\ADC_VDC.genclk.t0off_11 ));
    LocalMux I__13970 (
            .O(N__56531),
            .I(\ADC_VDC.genclk.t0off_11 ));
    InMux I__13969 (
            .O(N__56526),
            .I(N__56523));
    LocalMux I__13968 (
            .O(N__56523),
            .I(N__56520));
    Odrv4 I__13967 (
            .O(N__56520),
            .I(\ADC_VDC.genclk.n28 ));
    InMux I__13966 (
            .O(N__56517),
            .I(N__56514));
    LocalMux I__13965 (
            .O(N__56514),
            .I(\ADC_VDC.genclk.n26_adj_1448 ));
    InMux I__13964 (
            .O(N__56511),
            .I(N__56508));
    LocalMux I__13963 (
            .O(N__56508),
            .I(N__56505));
    Span4Mux_v I__13962 (
            .O(N__56505),
            .I(N__56500));
    InMux I__13961 (
            .O(N__56504),
            .I(N__56497));
    InMux I__13960 (
            .O(N__56503),
            .I(N__56494));
    Odrv4 I__13959 (
            .O(N__56500),
            .I(\comm_spi.n23101 ));
    LocalMux I__13958 (
            .O(N__56497),
            .I(\comm_spi.n23101 ));
    LocalMux I__13957 (
            .O(N__56494),
            .I(\comm_spi.n23101 ));
    InMux I__13956 (
            .O(N__56487),
            .I(N__56483));
    InMux I__13955 (
            .O(N__56486),
            .I(N__56480));
    LocalMux I__13954 (
            .O(N__56483),
            .I(N__56477));
    LocalMux I__13953 (
            .O(N__56480),
            .I(N__56474));
    Span4Mux_h I__13952 (
            .O(N__56477),
            .I(N__56469));
    Span4Mux_v I__13951 (
            .O(N__56474),
            .I(N__56469));
    Odrv4 I__13950 (
            .O(N__56469),
            .I(\comm_spi.n14834 ));
    SRMux I__13949 (
            .O(N__56466),
            .I(N__56463));
    LocalMux I__13948 (
            .O(N__56463),
            .I(N__56460));
    Odrv12 I__13947 (
            .O(N__56460),
            .I(\comm_spi.data_tx_7__N_823 ));
    SRMux I__13946 (
            .O(N__56457),
            .I(N__56454));
    LocalMux I__13945 (
            .O(N__56454),
            .I(N__56451));
    Odrv12 I__13944 (
            .O(N__56451),
            .I(\comm_spi.data_tx_7__N_811 ));
    InMux I__13943 (
            .O(N__56448),
            .I(N__56443));
    InMux I__13942 (
            .O(N__56447),
            .I(N__56438));
    InMux I__13941 (
            .O(N__56446),
            .I(N__56438));
    LocalMux I__13940 (
            .O(N__56443),
            .I(N__56435));
    LocalMux I__13939 (
            .O(N__56438),
            .I(N__56432));
    Span4Mux_h I__13938 (
            .O(N__56435),
            .I(N__56429));
    Span4Mux_h I__13937 (
            .O(N__56432),
            .I(N__56426));
    Odrv4 I__13936 (
            .O(N__56429),
            .I(comm_tx_buf_4));
    Odrv4 I__13935 (
            .O(N__56426),
            .I(comm_tx_buf_4));
    SRMux I__13934 (
            .O(N__56421),
            .I(N__56418));
    LocalMux I__13933 (
            .O(N__56418),
            .I(N__56415));
    Span4Mux_v I__13932 (
            .O(N__56415),
            .I(N__56412));
    Span4Mux_h I__13931 (
            .O(N__56412),
            .I(N__56409));
    Span4Mux_h I__13930 (
            .O(N__56409),
            .I(N__56406));
    Odrv4 I__13929 (
            .O(N__56406),
            .I(\comm_spi.data_tx_7__N_809 ));
    InMux I__13928 (
            .O(N__56403),
            .I(N__56394));
    InMux I__13927 (
            .O(N__56402),
            .I(N__56394));
    InMux I__13926 (
            .O(N__56401),
            .I(N__56394));
    LocalMux I__13925 (
            .O(N__56394),
            .I(N__56391));
    Span4Mux_v I__13924 (
            .O(N__56391),
            .I(N__56388));
    Odrv4 I__13923 (
            .O(N__56388),
            .I(comm_tx_buf_2));
    CascadeMux I__13922 (
            .O(N__56385),
            .I(N__56382));
    InMux I__13921 (
            .O(N__56382),
            .I(N__56378));
    InMux I__13920 (
            .O(N__56381),
            .I(N__56375));
    LocalMux I__13919 (
            .O(N__56378),
            .I(\ADC_VDC.genclk.t0off_6 ));
    LocalMux I__13918 (
            .O(N__56375),
            .I(\ADC_VDC.genclk.t0off_6 ));
    InMux I__13917 (
            .O(N__56370),
            .I(N__56366));
    InMux I__13916 (
            .O(N__56369),
            .I(N__56363));
    LocalMux I__13915 (
            .O(N__56366),
            .I(\ADC_VDC.genclk.t0off_1 ));
    LocalMux I__13914 (
            .O(N__56363),
            .I(\ADC_VDC.genclk.t0off_1 ));
    CascadeMux I__13913 (
            .O(N__56358),
            .I(N__56354));
    CascadeMux I__13912 (
            .O(N__56357),
            .I(N__56351));
    InMux I__13911 (
            .O(N__56354),
            .I(N__56348));
    InMux I__13910 (
            .O(N__56351),
            .I(N__56345));
    LocalMux I__13909 (
            .O(N__56348),
            .I(\ADC_VDC.genclk.t0off_4 ));
    LocalMux I__13908 (
            .O(N__56345),
            .I(\ADC_VDC.genclk.t0off_4 ));
    InMux I__13907 (
            .O(N__56340),
            .I(N__56336));
    InMux I__13906 (
            .O(N__56339),
            .I(N__56333));
    LocalMux I__13905 (
            .O(N__56336),
            .I(\ADC_VDC.genclk.t0off_0 ));
    LocalMux I__13904 (
            .O(N__56333),
            .I(\ADC_VDC.genclk.t0off_0 ));
    InMux I__13903 (
            .O(N__56328),
            .I(N__56325));
    LocalMux I__13902 (
            .O(N__56325),
            .I(\ADC_VDC.genclk.n21600 ));
    CascadeMux I__13901 (
            .O(N__56322),
            .I(\ADC_VDC.genclk.n27_adj_1449_cascade_ ));
    InMux I__13900 (
            .O(N__56319),
            .I(N__56316));
    LocalMux I__13899 (
            .O(N__56316),
            .I(\ADC_VDC.genclk.n21597 ));
    InMux I__13898 (
            .O(N__56313),
            .I(N__56310));
    LocalMux I__13897 (
            .O(N__56310),
            .I(\ADC_VDC.genclk.n21598 ));
    CascadeMux I__13896 (
            .O(N__56307),
            .I(\ADC_VDC.genclk.n21597_cascade_ ));
    InMux I__13895 (
            .O(N__56304),
            .I(N__56301));
    LocalMux I__13894 (
            .O(N__56301),
            .I(\ADC_VDC.genclk.n21603 ));
    CascadeMux I__13893 (
            .O(N__56298),
            .I(N__56294));
    InMux I__13892 (
            .O(N__56297),
            .I(N__56291));
    InMux I__13891 (
            .O(N__56294),
            .I(N__56288));
    LocalMux I__13890 (
            .O(N__56291),
            .I(N__56285));
    LocalMux I__13889 (
            .O(N__56288),
            .I(\ADC_VDC.genclk.t0off_13 ));
    Odrv4 I__13888 (
            .O(N__56285),
            .I(\ADC_VDC.genclk.t0off_13 ));
    InMux I__13887 (
            .O(N__56280),
            .I(N__56276));
    InMux I__13886 (
            .O(N__56279),
            .I(N__56273));
    LocalMux I__13885 (
            .O(N__56276),
            .I(N__56270));
    LocalMux I__13884 (
            .O(N__56273),
            .I(\ADC_VDC.genclk.t0off_3 ));
    Odrv4 I__13883 (
            .O(N__56270),
            .I(\ADC_VDC.genclk.t0off_3 ));
    CascadeMux I__13882 (
            .O(N__56265),
            .I(N__56261));
    InMux I__13881 (
            .O(N__56264),
            .I(N__56258));
    InMux I__13880 (
            .O(N__56261),
            .I(N__56255));
    LocalMux I__13879 (
            .O(N__56258),
            .I(\ADC_VDC.genclk.t0off_5 ));
    LocalMux I__13878 (
            .O(N__56255),
            .I(\ADC_VDC.genclk.t0off_5 ));
    InMux I__13877 (
            .O(N__56250),
            .I(N__56246));
    InMux I__13876 (
            .O(N__56249),
            .I(N__56243));
    LocalMux I__13875 (
            .O(N__56246),
            .I(\ADC_VDC.genclk.t0off_8 ));
    LocalMux I__13874 (
            .O(N__56243),
            .I(\ADC_VDC.genclk.t0off_8 ));
    InMux I__13873 (
            .O(N__56238),
            .I(N__56235));
    LocalMux I__13872 (
            .O(N__56235),
            .I(\ADC_VDC.genclk.n26 ));
    InMux I__13871 (
            .O(N__56232),
            .I(N__56225));
    InMux I__13870 (
            .O(N__56231),
            .I(N__56222));
    InMux I__13869 (
            .O(N__56230),
            .I(N__56217));
    InMux I__13868 (
            .O(N__56229),
            .I(N__56217));
    InMux I__13867 (
            .O(N__56228),
            .I(N__56214));
    LocalMux I__13866 (
            .O(N__56225),
            .I(\ADC_VDC.genclk.div_state_0 ));
    LocalMux I__13865 (
            .O(N__56222),
            .I(\ADC_VDC.genclk.div_state_0 ));
    LocalMux I__13864 (
            .O(N__56217),
            .I(\ADC_VDC.genclk.div_state_0 ));
    LocalMux I__13863 (
            .O(N__56214),
            .I(\ADC_VDC.genclk.div_state_0 ));
    InMux I__13862 (
            .O(N__56205),
            .I(N__56202));
    LocalMux I__13861 (
            .O(N__56202),
            .I(\ADC_VDC.genclk.n28_adj_1447 ));
    InMux I__13860 (
            .O(N__56199),
            .I(N__56195));
    InMux I__13859 (
            .O(N__56198),
            .I(N__56192));
    LocalMux I__13858 (
            .O(N__56195),
            .I(N__56187));
    LocalMux I__13857 (
            .O(N__56192),
            .I(N__56187));
    Odrv4 I__13856 (
            .O(N__56187),
            .I(\ADC_VDC.genclk.t0off_14 ));
    CascadeMux I__13855 (
            .O(N__56184),
            .I(N__56181));
    InMux I__13854 (
            .O(N__56181),
            .I(N__56177));
    InMux I__13853 (
            .O(N__56180),
            .I(N__56174));
    LocalMux I__13852 (
            .O(N__56177),
            .I(\ADC_VDC.genclk.t0off_9 ));
    LocalMux I__13851 (
            .O(N__56174),
            .I(\ADC_VDC.genclk.t0off_9 ));
    CascadeMux I__13850 (
            .O(N__56169),
            .I(N__56165));
    InMux I__13849 (
            .O(N__56168),
            .I(N__56162));
    InMux I__13848 (
            .O(N__56165),
            .I(N__56159));
    LocalMux I__13847 (
            .O(N__56162),
            .I(\ADC_VDC.genclk.t0off_15 ));
    LocalMux I__13846 (
            .O(N__56159),
            .I(\ADC_VDC.genclk.t0off_15 ));
    InMux I__13845 (
            .O(N__56154),
            .I(N__56151));
    LocalMux I__13844 (
            .O(N__56151),
            .I(N__56148));
    Span4Mux_v I__13843 (
            .O(N__56148),
            .I(N__56144));
    InMux I__13842 (
            .O(N__56147),
            .I(N__56141));
    Span4Mux_v I__13841 (
            .O(N__56144),
            .I(N__56135));
    LocalMux I__13840 (
            .O(N__56141),
            .I(N__56135));
    InMux I__13839 (
            .O(N__56140),
            .I(N__56132));
    Span4Mux_v I__13838 (
            .O(N__56135),
            .I(N__56129));
    LocalMux I__13837 (
            .O(N__56132),
            .I(N__56126));
    Sp12to4 I__13836 (
            .O(N__56129),
            .I(N__56121));
    Span12Mux_v I__13835 (
            .O(N__56126),
            .I(N__56121));
    Odrv12 I__13834 (
            .O(N__56121),
            .I(comm_tx_buf_3));
    IoInMux I__13833 (
            .O(N__56118),
            .I(N__56115));
    LocalMux I__13832 (
            .O(N__56115),
            .I(N__56112));
    Span12Mux_s9_h I__13831 (
            .O(N__56112),
            .I(N__56109));
    Span12Mux_v I__13830 (
            .O(N__56109),
            .I(N__56106));
    Odrv12 I__13829 (
            .O(N__56106),
            .I(ICE_GPMI_0));
    ClkMux I__13828 (
            .O(N__56103),
            .I(N__55602));
    ClkMux I__13827 (
            .O(N__56102),
            .I(N__55602));
    ClkMux I__13826 (
            .O(N__56101),
            .I(N__55602));
    ClkMux I__13825 (
            .O(N__56100),
            .I(N__55602));
    ClkMux I__13824 (
            .O(N__56099),
            .I(N__55602));
    ClkMux I__13823 (
            .O(N__56098),
            .I(N__55602));
    ClkMux I__13822 (
            .O(N__56097),
            .I(N__55602));
    ClkMux I__13821 (
            .O(N__56096),
            .I(N__55602));
    ClkMux I__13820 (
            .O(N__56095),
            .I(N__55602));
    ClkMux I__13819 (
            .O(N__56094),
            .I(N__55602));
    ClkMux I__13818 (
            .O(N__56093),
            .I(N__55602));
    ClkMux I__13817 (
            .O(N__56092),
            .I(N__55602));
    ClkMux I__13816 (
            .O(N__56091),
            .I(N__55602));
    ClkMux I__13815 (
            .O(N__56090),
            .I(N__55602));
    ClkMux I__13814 (
            .O(N__56089),
            .I(N__55602));
    ClkMux I__13813 (
            .O(N__56088),
            .I(N__55602));
    ClkMux I__13812 (
            .O(N__56087),
            .I(N__55602));
    ClkMux I__13811 (
            .O(N__56086),
            .I(N__55602));
    ClkMux I__13810 (
            .O(N__56085),
            .I(N__55602));
    ClkMux I__13809 (
            .O(N__56084),
            .I(N__55602));
    ClkMux I__13808 (
            .O(N__56083),
            .I(N__55602));
    ClkMux I__13807 (
            .O(N__56082),
            .I(N__55602));
    ClkMux I__13806 (
            .O(N__56081),
            .I(N__55602));
    ClkMux I__13805 (
            .O(N__56080),
            .I(N__55602));
    ClkMux I__13804 (
            .O(N__56079),
            .I(N__55602));
    ClkMux I__13803 (
            .O(N__56078),
            .I(N__55602));
    ClkMux I__13802 (
            .O(N__56077),
            .I(N__55602));
    ClkMux I__13801 (
            .O(N__56076),
            .I(N__55602));
    ClkMux I__13800 (
            .O(N__56075),
            .I(N__55602));
    ClkMux I__13799 (
            .O(N__56074),
            .I(N__55602));
    ClkMux I__13798 (
            .O(N__56073),
            .I(N__55602));
    ClkMux I__13797 (
            .O(N__56072),
            .I(N__55602));
    ClkMux I__13796 (
            .O(N__56071),
            .I(N__55602));
    ClkMux I__13795 (
            .O(N__56070),
            .I(N__55602));
    ClkMux I__13794 (
            .O(N__56069),
            .I(N__55602));
    ClkMux I__13793 (
            .O(N__56068),
            .I(N__55602));
    ClkMux I__13792 (
            .O(N__56067),
            .I(N__55602));
    ClkMux I__13791 (
            .O(N__56066),
            .I(N__55602));
    ClkMux I__13790 (
            .O(N__56065),
            .I(N__55602));
    ClkMux I__13789 (
            .O(N__56064),
            .I(N__55602));
    ClkMux I__13788 (
            .O(N__56063),
            .I(N__55602));
    ClkMux I__13787 (
            .O(N__56062),
            .I(N__55602));
    ClkMux I__13786 (
            .O(N__56061),
            .I(N__55602));
    ClkMux I__13785 (
            .O(N__56060),
            .I(N__55602));
    ClkMux I__13784 (
            .O(N__56059),
            .I(N__55602));
    ClkMux I__13783 (
            .O(N__56058),
            .I(N__55602));
    ClkMux I__13782 (
            .O(N__56057),
            .I(N__55602));
    ClkMux I__13781 (
            .O(N__56056),
            .I(N__55602));
    ClkMux I__13780 (
            .O(N__56055),
            .I(N__55602));
    ClkMux I__13779 (
            .O(N__56054),
            .I(N__55602));
    ClkMux I__13778 (
            .O(N__56053),
            .I(N__55602));
    ClkMux I__13777 (
            .O(N__56052),
            .I(N__55602));
    ClkMux I__13776 (
            .O(N__56051),
            .I(N__55602));
    ClkMux I__13775 (
            .O(N__56050),
            .I(N__55602));
    ClkMux I__13774 (
            .O(N__56049),
            .I(N__55602));
    ClkMux I__13773 (
            .O(N__56048),
            .I(N__55602));
    ClkMux I__13772 (
            .O(N__56047),
            .I(N__55602));
    ClkMux I__13771 (
            .O(N__56046),
            .I(N__55602));
    ClkMux I__13770 (
            .O(N__56045),
            .I(N__55602));
    ClkMux I__13769 (
            .O(N__56044),
            .I(N__55602));
    ClkMux I__13768 (
            .O(N__56043),
            .I(N__55602));
    ClkMux I__13767 (
            .O(N__56042),
            .I(N__55602));
    ClkMux I__13766 (
            .O(N__56041),
            .I(N__55602));
    ClkMux I__13765 (
            .O(N__56040),
            .I(N__55602));
    ClkMux I__13764 (
            .O(N__56039),
            .I(N__55602));
    ClkMux I__13763 (
            .O(N__56038),
            .I(N__55602));
    ClkMux I__13762 (
            .O(N__56037),
            .I(N__55602));
    ClkMux I__13761 (
            .O(N__56036),
            .I(N__55602));
    ClkMux I__13760 (
            .O(N__56035),
            .I(N__55602));
    ClkMux I__13759 (
            .O(N__56034),
            .I(N__55602));
    ClkMux I__13758 (
            .O(N__56033),
            .I(N__55602));
    ClkMux I__13757 (
            .O(N__56032),
            .I(N__55602));
    ClkMux I__13756 (
            .O(N__56031),
            .I(N__55602));
    ClkMux I__13755 (
            .O(N__56030),
            .I(N__55602));
    ClkMux I__13754 (
            .O(N__56029),
            .I(N__55602));
    ClkMux I__13753 (
            .O(N__56028),
            .I(N__55602));
    ClkMux I__13752 (
            .O(N__56027),
            .I(N__55602));
    ClkMux I__13751 (
            .O(N__56026),
            .I(N__55602));
    ClkMux I__13750 (
            .O(N__56025),
            .I(N__55602));
    ClkMux I__13749 (
            .O(N__56024),
            .I(N__55602));
    ClkMux I__13748 (
            .O(N__56023),
            .I(N__55602));
    ClkMux I__13747 (
            .O(N__56022),
            .I(N__55602));
    ClkMux I__13746 (
            .O(N__56021),
            .I(N__55602));
    ClkMux I__13745 (
            .O(N__56020),
            .I(N__55602));
    ClkMux I__13744 (
            .O(N__56019),
            .I(N__55602));
    ClkMux I__13743 (
            .O(N__56018),
            .I(N__55602));
    ClkMux I__13742 (
            .O(N__56017),
            .I(N__55602));
    ClkMux I__13741 (
            .O(N__56016),
            .I(N__55602));
    ClkMux I__13740 (
            .O(N__56015),
            .I(N__55602));
    ClkMux I__13739 (
            .O(N__56014),
            .I(N__55602));
    ClkMux I__13738 (
            .O(N__56013),
            .I(N__55602));
    ClkMux I__13737 (
            .O(N__56012),
            .I(N__55602));
    ClkMux I__13736 (
            .O(N__56011),
            .I(N__55602));
    ClkMux I__13735 (
            .O(N__56010),
            .I(N__55602));
    ClkMux I__13734 (
            .O(N__56009),
            .I(N__55602));
    ClkMux I__13733 (
            .O(N__56008),
            .I(N__55602));
    ClkMux I__13732 (
            .O(N__56007),
            .I(N__55602));
    ClkMux I__13731 (
            .O(N__56006),
            .I(N__55602));
    ClkMux I__13730 (
            .O(N__56005),
            .I(N__55602));
    ClkMux I__13729 (
            .O(N__56004),
            .I(N__55602));
    ClkMux I__13728 (
            .O(N__56003),
            .I(N__55602));
    ClkMux I__13727 (
            .O(N__56002),
            .I(N__55602));
    ClkMux I__13726 (
            .O(N__56001),
            .I(N__55602));
    ClkMux I__13725 (
            .O(N__56000),
            .I(N__55602));
    ClkMux I__13724 (
            .O(N__55999),
            .I(N__55602));
    ClkMux I__13723 (
            .O(N__55998),
            .I(N__55602));
    ClkMux I__13722 (
            .O(N__55997),
            .I(N__55602));
    ClkMux I__13721 (
            .O(N__55996),
            .I(N__55602));
    ClkMux I__13720 (
            .O(N__55995),
            .I(N__55602));
    ClkMux I__13719 (
            .O(N__55994),
            .I(N__55602));
    ClkMux I__13718 (
            .O(N__55993),
            .I(N__55602));
    ClkMux I__13717 (
            .O(N__55992),
            .I(N__55602));
    ClkMux I__13716 (
            .O(N__55991),
            .I(N__55602));
    ClkMux I__13715 (
            .O(N__55990),
            .I(N__55602));
    ClkMux I__13714 (
            .O(N__55989),
            .I(N__55602));
    ClkMux I__13713 (
            .O(N__55988),
            .I(N__55602));
    ClkMux I__13712 (
            .O(N__55987),
            .I(N__55602));
    ClkMux I__13711 (
            .O(N__55986),
            .I(N__55602));
    ClkMux I__13710 (
            .O(N__55985),
            .I(N__55602));
    ClkMux I__13709 (
            .O(N__55984),
            .I(N__55602));
    ClkMux I__13708 (
            .O(N__55983),
            .I(N__55602));
    ClkMux I__13707 (
            .O(N__55982),
            .I(N__55602));
    ClkMux I__13706 (
            .O(N__55981),
            .I(N__55602));
    ClkMux I__13705 (
            .O(N__55980),
            .I(N__55602));
    ClkMux I__13704 (
            .O(N__55979),
            .I(N__55602));
    ClkMux I__13703 (
            .O(N__55978),
            .I(N__55602));
    ClkMux I__13702 (
            .O(N__55977),
            .I(N__55602));
    ClkMux I__13701 (
            .O(N__55976),
            .I(N__55602));
    ClkMux I__13700 (
            .O(N__55975),
            .I(N__55602));
    ClkMux I__13699 (
            .O(N__55974),
            .I(N__55602));
    ClkMux I__13698 (
            .O(N__55973),
            .I(N__55602));
    ClkMux I__13697 (
            .O(N__55972),
            .I(N__55602));
    ClkMux I__13696 (
            .O(N__55971),
            .I(N__55602));
    ClkMux I__13695 (
            .O(N__55970),
            .I(N__55602));
    ClkMux I__13694 (
            .O(N__55969),
            .I(N__55602));
    ClkMux I__13693 (
            .O(N__55968),
            .I(N__55602));
    ClkMux I__13692 (
            .O(N__55967),
            .I(N__55602));
    ClkMux I__13691 (
            .O(N__55966),
            .I(N__55602));
    ClkMux I__13690 (
            .O(N__55965),
            .I(N__55602));
    ClkMux I__13689 (
            .O(N__55964),
            .I(N__55602));
    ClkMux I__13688 (
            .O(N__55963),
            .I(N__55602));
    ClkMux I__13687 (
            .O(N__55962),
            .I(N__55602));
    ClkMux I__13686 (
            .O(N__55961),
            .I(N__55602));
    ClkMux I__13685 (
            .O(N__55960),
            .I(N__55602));
    ClkMux I__13684 (
            .O(N__55959),
            .I(N__55602));
    ClkMux I__13683 (
            .O(N__55958),
            .I(N__55602));
    ClkMux I__13682 (
            .O(N__55957),
            .I(N__55602));
    ClkMux I__13681 (
            .O(N__55956),
            .I(N__55602));
    ClkMux I__13680 (
            .O(N__55955),
            .I(N__55602));
    ClkMux I__13679 (
            .O(N__55954),
            .I(N__55602));
    ClkMux I__13678 (
            .O(N__55953),
            .I(N__55602));
    ClkMux I__13677 (
            .O(N__55952),
            .I(N__55602));
    ClkMux I__13676 (
            .O(N__55951),
            .I(N__55602));
    ClkMux I__13675 (
            .O(N__55950),
            .I(N__55602));
    ClkMux I__13674 (
            .O(N__55949),
            .I(N__55602));
    ClkMux I__13673 (
            .O(N__55948),
            .I(N__55602));
    ClkMux I__13672 (
            .O(N__55947),
            .I(N__55602));
    ClkMux I__13671 (
            .O(N__55946),
            .I(N__55602));
    ClkMux I__13670 (
            .O(N__55945),
            .I(N__55602));
    ClkMux I__13669 (
            .O(N__55944),
            .I(N__55602));
    ClkMux I__13668 (
            .O(N__55943),
            .I(N__55602));
    ClkMux I__13667 (
            .O(N__55942),
            .I(N__55602));
    ClkMux I__13666 (
            .O(N__55941),
            .I(N__55602));
    ClkMux I__13665 (
            .O(N__55940),
            .I(N__55602));
    ClkMux I__13664 (
            .O(N__55939),
            .I(N__55602));
    ClkMux I__13663 (
            .O(N__55938),
            .I(N__55602));
    ClkMux I__13662 (
            .O(N__55937),
            .I(N__55602));
    GlobalMux I__13661 (
            .O(N__55602),
            .I(clk_32MHz));
    CEMux I__13660 (
            .O(N__55599),
            .I(N__55596));
    LocalMux I__13659 (
            .O(N__55596),
            .I(N__55593));
    Span4Mux_v I__13658 (
            .O(N__55593),
            .I(N__55590));
    Span4Mux_h I__13657 (
            .O(N__55590),
            .I(N__55587));
    Sp12to4 I__13656 (
            .O(N__55587),
            .I(N__55584));
    Span12Mux_s10_h I__13655 (
            .O(N__55584),
            .I(N__55581));
    Odrv12 I__13654 (
            .O(N__55581),
            .I(n11600));
    InMux I__13653 (
            .O(N__55578),
            .I(N__55575));
    LocalMux I__13652 (
            .O(N__55575),
            .I(N__55568));
    InMux I__13651 (
            .O(N__55574),
            .I(N__55565));
    InMux I__13650 (
            .O(N__55573),
            .I(N__55559));
    InMux I__13649 (
            .O(N__55572),
            .I(N__55554));
    InMux I__13648 (
            .O(N__55571),
            .I(N__55554));
    Span4Mux_v I__13647 (
            .O(N__55568),
            .I(N__55548));
    LocalMux I__13646 (
            .O(N__55565),
            .I(N__55548));
    InMux I__13645 (
            .O(N__55564),
            .I(N__55545));
    InMux I__13644 (
            .O(N__55563),
            .I(N__55541));
    InMux I__13643 (
            .O(N__55562),
            .I(N__55538));
    LocalMux I__13642 (
            .O(N__55559),
            .I(N__55533));
    LocalMux I__13641 (
            .O(N__55554),
            .I(N__55530));
    InMux I__13640 (
            .O(N__55553),
            .I(N__55527));
    Span4Mux_h I__13639 (
            .O(N__55548),
            .I(N__55524));
    LocalMux I__13638 (
            .O(N__55545),
            .I(N__55521));
    InMux I__13637 (
            .O(N__55544),
            .I(N__55518));
    LocalMux I__13636 (
            .O(N__55541),
            .I(N__55513));
    LocalMux I__13635 (
            .O(N__55538),
            .I(N__55513));
    InMux I__13634 (
            .O(N__55537),
            .I(N__55508));
    InMux I__13633 (
            .O(N__55536),
            .I(N__55508));
    Span4Mux_h I__13632 (
            .O(N__55533),
            .I(N__55503));
    Span4Mux_v I__13631 (
            .O(N__55530),
            .I(N__55503));
    LocalMux I__13630 (
            .O(N__55527),
            .I(N__55496));
    Span4Mux_v I__13629 (
            .O(N__55524),
            .I(N__55496));
    Span4Mux_h I__13628 (
            .O(N__55521),
            .I(N__55496));
    LocalMux I__13627 (
            .O(N__55518),
            .I(N__55489));
    Span12Mux_v I__13626 (
            .O(N__55513),
            .I(N__55489));
    LocalMux I__13625 (
            .O(N__55508),
            .I(N__55489));
    Odrv4 I__13624 (
            .O(N__55503),
            .I(n12433));
    Odrv4 I__13623 (
            .O(N__55496),
            .I(n12433));
    Odrv12 I__13622 (
            .O(N__55489),
            .I(n12433));
    CascadeMux I__13621 (
            .O(N__55482),
            .I(n10_adj_1619_cascade_));
    CascadeMux I__13620 (
            .O(N__55479),
            .I(N__55475));
    SRMux I__13619 (
            .O(N__55478),
            .I(N__55456));
    InMux I__13618 (
            .O(N__55475),
            .I(N__55452));
    InMux I__13617 (
            .O(N__55474),
            .I(N__55441));
    InMux I__13616 (
            .O(N__55473),
            .I(N__55441));
    InMux I__13615 (
            .O(N__55472),
            .I(N__55441));
    InMux I__13614 (
            .O(N__55471),
            .I(N__55441));
    InMux I__13613 (
            .O(N__55470),
            .I(N__55441));
    CascadeMux I__13612 (
            .O(N__55469),
            .I(N__55424));
    CascadeMux I__13611 (
            .O(N__55468),
            .I(N__55415));
    CascadeMux I__13610 (
            .O(N__55467),
            .I(N__55411));
    CascadeMux I__13609 (
            .O(N__55466),
            .I(N__55407));
    CascadeMux I__13608 (
            .O(N__55465),
            .I(N__55403));
    InMux I__13607 (
            .O(N__55464),
            .I(N__55399));
    CascadeMux I__13606 (
            .O(N__55463),
            .I(N__55396));
    InMux I__13605 (
            .O(N__55462),
            .I(N__55389));
    InMux I__13604 (
            .O(N__55461),
            .I(N__55389));
    InMux I__13603 (
            .O(N__55460),
            .I(N__55389));
    InMux I__13602 (
            .O(N__55459),
            .I(N__55384));
    LocalMux I__13601 (
            .O(N__55456),
            .I(N__55381));
    InMux I__13600 (
            .O(N__55455),
            .I(N__55378));
    LocalMux I__13599 (
            .O(N__55452),
            .I(N__55373));
    LocalMux I__13598 (
            .O(N__55441),
            .I(N__55373));
    InMux I__13597 (
            .O(N__55440),
            .I(N__55368));
    InMux I__13596 (
            .O(N__55439),
            .I(N__55368));
    InMux I__13595 (
            .O(N__55438),
            .I(N__55359));
    InMux I__13594 (
            .O(N__55437),
            .I(N__55359));
    InMux I__13593 (
            .O(N__55436),
            .I(N__55359));
    InMux I__13592 (
            .O(N__55435),
            .I(N__55359));
    CascadeMux I__13591 (
            .O(N__55434),
            .I(N__55355));
    InMux I__13590 (
            .O(N__55433),
            .I(N__55352));
    InMux I__13589 (
            .O(N__55432),
            .I(N__55347));
    InMux I__13588 (
            .O(N__55431),
            .I(N__55347));
    InMux I__13587 (
            .O(N__55430),
            .I(N__55343));
    InMux I__13586 (
            .O(N__55429),
            .I(N__55336));
    InMux I__13585 (
            .O(N__55428),
            .I(N__55336));
    InMux I__13584 (
            .O(N__55427),
            .I(N__55336));
    InMux I__13583 (
            .O(N__55424),
            .I(N__55325));
    InMux I__13582 (
            .O(N__55423),
            .I(N__55325));
    InMux I__13581 (
            .O(N__55422),
            .I(N__55325));
    InMux I__13580 (
            .O(N__55421),
            .I(N__55325));
    InMux I__13579 (
            .O(N__55420),
            .I(N__55325));
    InMux I__13578 (
            .O(N__55419),
            .I(N__55322));
    InMux I__13577 (
            .O(N__55418),
            .I(N__55319));
    InMux I__13576 (
            .O(N__55415),
            .I(N__55302));
    InMux I__13575 (
            .O(N__55414),
            .I(N__55302));
    InMux I__13574 (
            .O(N__55411),
            .I(N__55302));
    InMux I__13573 (
            .O(N__55410),
            .I(N__55302));
    InMux I__13572 (
            .O(N__55407),
            .I(N__55302));
    InMux I__13571 (
            .O(N__55406),
            .I(N__55302));
    InMux I__13570 (
            .O(N__55403),
            .I(N__55302));
    InMux I__13569 (
            .O(N__55402),
            .I(N__55302));
    LocalMux I__13568 (
            .O(N__55399),
            .I(N__55299));
    InMux I__13567 (
            .O(N__55396),
            .I(N__55289));
    LocalMux I__13566 (
            .O(N__55389),
            .I(N__55282));
    CascadeMux I__13565 (
            .O(N__55388),
            .I(N__55276));
    InMux I__13564 (
            .O(N__55387),
            .I(N__55273));
    LocalMux I__13563 (
            .O(N__55384),
            .I(N__55255));
    Span4Mux_v I__13562 (
            .O(N__55381),
            .I(N__55255));
    LocalMux I__13561 (
            .O(N__55378),
            .I(N__55255));
    Span4Mux_v I__13560 (
            .O(N__55373),
            .I(N__55255));
    LocalMux I__13559 (
            .O(N__55368),
            .I(N__55255));
    LocalMux I__13558 (
            .O(N__55359),
            .I(N__55255));
    CascadeMux I__13557 (
            .O(N__55358),
            .I(N__55252));
    InMux I__13556 (
            .O(N__55355),
            .I(N__55244));
    LocalMux I__13555 (
            .O(N__55352),
            .I(N__55239));
    LocalMux I__13554 (
            .O(N__55347),
            .I(N__55239));
    InMux I__13553 (
            .O(N__55346),
            .I(N__55230));
    LocalMux I__13552 (
            .O(N__55343),
            .I(N__55227));
    LocalMux I__13551 (
            .O(N__55336),
            .I(N__55216));
    LocalMux I__13550 (
            .O(N__55325),
            .I(N__55216));
    LocalMux I__13549 (
            .O(N__55322),
            .I(N__55216));
    LocalMux I__13548 (
            .O(N__55319),
            .I(N__55216));
    LocalMux I__13547 (
            .O(N__55302),
            .I(N__55216));
    Span4Mux_v I__13546 (
            .O(N__55299),
            .I(N__55213));
    InMux I__13545 (
            .O(N__55298),
            .I(N__55208));
    InMux I__13544 (
            .O(N__55297),
            .I(N__55208));
    InMux I__13543 (
            .O(N__55296),
            .I(N__55204));
    InMux I__13542 (
            .O(N__55295),
            .I(N__55195));
    InMux I__13541 (
            .O(N__55294),
            .I(N__55195));
    InMux I__13540 (
            .O(N__55293),
            .I(N__55195));
    InMux I__13539 (
            .O(N__55292),
            .I(N__55195));
    LocalMux I__13538 (
            .O(N__55289),
            .I(N__55192));
    InMux I__13537 (
            .O(N__55288),
            .I(N__55187));
    InMux I__13536 (
            .O(N__55287),
            .I(N__55187));
    InMux I__13535 (
            .O(N__55286),
            .I(N__55184));
    CascadeMux I__13534 (
            .O(N__55285),
            .I(N__55177));
    Span4Mux_h I__13533 (
            .O(N__55282),
            .I(N__55174));
    InMux I__13532 (
            .O(N__55281),
            .I(N__55171));
    InMux I__13531 (
            .O(N__55280),
            .I(N__55166));
    InMux I__13530 (
            .O(N__55279),
            .I(N__55166));
    InMux I__13529 (
            .O(N__55276),
            .I(N__55160));
    LocalMux I__13528 (
            .O(N__55273),
            .I(N__55157));
    InMux I__13527 (
            .O(N__55272),
            .I(N__55154));
    InMux I__13526 (
            .O(N__55271),
            .I(N__55149));
    InMux I__13525 (
            .O(N__55270),
            .I(N__55149));
    InMux I__13524 (
            .O(N__55269),
            .I(N__55144));
    InMux I__13523 (
            .O(N__55268),
            .I(N__55144));
    Span4Mux_v I__13522 (
            .O(N__55255),
            .I(N__55141));
    InMux I__13521 (
            .O(N__55252),
            .I(N__55136));
    InMux I__13520 (
            .O(N__55251),
            .I(N__55136));
    InMux I__13519 (
            .O(N__55250),
            .I(N__55131));
    InMux I__13518 (
            .O(N__55249),
            .I(N__55131));
    InMux I__13517 (
            .O(N__55248),
            .I(N__55126));
    InMux I__13516 (
            .O(N__55247),
            .I(N__55126));
    LocalMux I__13515 (
            .O(N__55244),
            .I(N__55121));
    Span4Mux_v I__13514 (
            .O(N__55239),
            .I(N__55121));
    InMux I__13513 (
            .O(N__55238),
            .I(N__55109));
    InMux I__13512 (
            .O(N__55237),
            .I(N__55109));
    InMux I__13511 (
            .O(N__55236),
            .I(N__55109));
    InMux I__13510 (
            .O(N__55235),
            .I(N__55109));
    InMux I__13509 (
            .O(N__55234),
            .I(N__55109));
    InMux I__13508 (
            .O(N__55233),
            .I(N__55105));
    LocalMux I__13507 (
            .O(N__55230),
            .I(N__55101));
    Span4Mux_h I__13506 (
            .O(N__55227),
            .I(N__55096));
    Span4Mux_v I__13505 (
            .O(N__55216),
            .I(N__55096));
    Span4Mux_h I__13504 (
            .O(N__55213),
            .I(N__55091));
    LocalMux I__13503 (
            .O(N__55208),
            .I(N__55091));
    InMux I__13502 (
            .O(N__55207),
            .I(N__55088));
    LocalMux I__13501 (
            .O(N__55204),
            .I(N__55085));
    LocalMux I__13500 (
            .O(N__55195),
            .I(N__55076));
    Span4Mux_v I__13499 (
            .O(N__55192),
            .I(N__55076));
    LocalMux I__13498 (
            .O(N__55187),
            .I(N__55076));
    LocalMux I__13497 (
            .O(N__55184),
            .I(N__55076));
    InMux I__13496 (
            .O(N__55183),
            .I(N__55069));
    InMux I__13495 (
            .O(N__55182),
            .I(N__55069));
    InMux I__13494 (
            .O(N__55181),
            .I(N__55069));
    InMux I__13493 (
            .O(N__55180),
            .I(N__55062));
    InMux I__13492 (
            .O(N__55177),
            .I(N__55059));
    Span4Mux_h I__13491 (
            .O(N__55174),
            .I(N__55056));
    LocalMux I__13490 (
            .O(N__55171),
            .I(N__55051));
    LocalMux I__13489 (
            .O(N__55166),
            .I(N__55051));
    InMux I__13488 (
            .O(N__55165),
            .I(N__55044));
    InMux I__13487 (
            .O(N__55164),
            .I(N__55044));
    InMux I__13486 (
            .O(N__55163),
            .I(N__55044));
    LocalMux I__13485 (
            .O(N__55160),
            .I(N__55033));
    Span4Mux_v I__13484 (
            .O(N__55157),
            .I(N__55033));
    LocalMux I__13483 (
            .O(N__55154),
            .I(N__55033));
    LocalMux I__13482 (
            .O(N__55149),
            .I(N__55033));
    LocalMux I__13481 (
            .O(N__55144),
            .I(N__55033));
    Span4Mux_h I__13480 (
            .O(N__55141),
            .I(N__55030));
    LocalMux I__13479 (
            .O(N__55136),
            .I(N__55024));
    LocalMux I__13478 (
            .O(N__55131),
            .I(N__55017));
    LocalMux I__13477 (
            .O(N__55126),
            .I(N__55017));
    Span4Mux_h I__13476 (
            .O(N__55121),
            .I(N__55017));
    InMux I__13475 (
            .O(N__55120),
            .I(N__55014));
    LocalMux I__13474 (
            .O(N__55109),
            .I(N__55011));
    InMux I__13473 (
            .O(N__55108),
            .I(N__55008));
    LocalMux I__13472 (
            .O(N__55105),
            .I(N__55005));
    InMux I__13471 (
            .O(N__55104),
            .I(N__55002));
    Span4Mux_v I__13470 (
            .O(N__55101),
            .I(N__54995));
    Span4Mux_h I__13469 (
            .O(N__55096),
            .I(N__54995));
    Span4Mux_v I__13468 (
            .O(N__55091),
            .I(N__54995));
    LocalMux I__13467 (
            .O(N__55088),
            .I(N__54990));
    Span4Mux_v I__13466 (
            .O(N__55085),
            .I(N__54990));
    Span4Mux_v I__13465 (
            .O(N__55076),
            .I(N__54985));
    LocalMux I__13464 (
            .O(N__55069),
            .I(N__54985));
    InMux I__13463 (
            .O(N__55068),
            .I(N__54980));
    InMux I__13462 (
            .O(N__55067),
            .I(N__54980));
    InMux I__13461 (
            .O(N__55066),
            .I(N__54977));
    InMux I__13460 (
            .O(N__55065),
            .I(N__54974));
    LocalMux I__13459 (
            .O(N__55062),
            .I(N__54965));
    LocalMux I__13458 (
            .O(N__55059),
            .I(N__54965));
    Span4Mux_h I__13457 (
            .O(N__55056),
            .I(N__54965));
    Span4Mux_v I__13456 (
            .O(N__55051),
            .I(N__54965));
    LocalMux I__13455 (
            .O(N__55044),
            .I(N__54958));
    Span4Mux_v I__13454 (
            .O(N__55033),
            .I(N__54958));
    Span4Mux_h I__13453 (
            .O(N__55030),
            .I(N__54958));
    InMux I__13452 (
            .O(N__55029),
            .I(N__54951));
    InMux I__13451 (
            .O(N__55028),
            .I(N__54951));
    InMux I__13450 (
            .O(N__55027),
            .I(N__54951));
    Span4Mux_v I__13449 (
            .O(N__55024),
            .I(N__54946));
    Span4Mux_v I__13448 (
            .O(N__55017),
            .I(N__54946));
    LocalMux I__13447 (
            .O(N__55014),
            .I(N__54941));
    Span4Mux_h I__13446 (
            .O(N__55011),
            .I(N__54941));
    LocalMux I__13445 (
            .O(N__55008),
            .I(N__54934));
    Span12Mux_v I__13444 (
            .O(N__55005),
            .I(N__54934));
    LocalMux I__13443 (
            .O(N__55002),
            .I(N__54934));
    Span4Mux_h I__13442 (
            .O(N__54995),
            .I(N__54931));
    Span4Mux_h I__13441 (
            .O(N__54990),
            .I(N__54924));
    Span4Mux_v I__13440 (
            .O(N__54985),
            .I(N__54924));
    LocalMux I__13439 (
            .O(N__54980),
            .I(N__54924));
    LocalMux I__13438 (
            .O(N__54977),
            .I(comm_state_3));
    LocalMux I__13437 (
            .O(N__54974),
            .I(comm_state_3));
    Odrv4 I__13436 (
            .O(N__54965),
            .I(comm_state_3));
    Odrv4 I__13435 (
            .O(N__54958),
            .I(comm_state_3));
    LocalMux I__13434 (
            .O(N__54951),
            .I(comm_state_3));
    Odrv4 I__13433 (
            .O(N__54946),
            .I(comm_state_3));
    Odrv4 I__13432 (
            .O(N__54941),
            .I(comm_state_3));
    Odrv12 I__13431 (
            .O(N__54934),
            .I(comm_state_3));
    Odrv4 I__13430 (
            .O(N__54931),
            .I(comm_state_3));
    Odrv4 I__13429 (
            .O(N__54924),
            .I(comm_state_3));
    CEMux I__13428 (
            .O(N__54903),
            .I(N__54900));
    LocalMux I__13427 (
            .O(N__54900),
            .I(N__54897));
    Odrv12 I__13426 (
            .O(N__54897),
            .I(n12079));
    CascadeMux I__13425 (
            .O(N__54894),
            .I(N__54888));
    InMux I__13424 (
            .O(N__54893),
            .I(N__54881));
    InMux I__13423 (
            .O(N__54892),
            .I(N__54876));
    InMux I__13422 (
            .O(N__54891),
            .I(N__54876));
    InMux I__13421 (
            .O(N__54888),
            .I(N__54871));
    InMux I__13420 (
            .O(N__54887),
            .I(N__54864));
    InMux I__13419 (
            .O(N__54886),
            .I(N__54864));
    InMux I__13418 (
            .O(N__54885),
            .I(N__54864));
    InMux I__13417 (
            .O(N__54884),
            .I(N__54854));
    LocalMux I__13416 (
            .O(N__54881),
            .I(N__54848));
    LocalMux I__13415 (
            .O(N__54876),
            .I(N__54844));
    InMux I__13414 (
            .O(N__54875),
            .I(N__54836));
    InMux I__13413 (
            .O(N__54874),
            .I(N__54833));
    LocalMux I__13412 (
            .O(N__54871),
            .I(N__54828));
    LocalMux I__13411 (
            .O(N__54864),
            .I(N__54828));
    InMux I__13410 (
            .O(N__54863),
            .I(N__54822));
    InMux I__13409 (
            .O(N__54862),
            .I(N__54811));
    InMux I__13408 (
            .O(N__54861),
            .I(N__54811));
    InMux I__13407 (
            .O(N__54860),
            .I(N__54811));
    InMux I__13406 (
            .O(N__54859),
            .I(N__54811));
    InMux I__13405 (
            .O(N__54858),
            .I(N__54811));
    InMux I__13404 (
            .O(N__54857),
            .I(N__54807));
    LocalMux I__13403 (
            .O(N__54854),
            .I(N__54804));
    CascadeMux I__13402 (
            .O(N__54853),
            .I(N__54800));
    CascadeMux I__13401 (
            .O(N__54852),
            .I(N__54797));
    InMux I__13400 (
            .O(N__54851),
            .I(N__54792));
    Span4Mux_h I__13399 (
            .O(N__54848),
            .I(N__54789));
    InMux I__13398 (
            .O(N__54847),
            .I(N__54784));
    Span4Mux_h I__13397 (
            .O(N__54844),
            .I(N__54781));
    InMux I__13396 (
            .O(N__54843),
            .I(N__54778));
    CascadeMux I__13395 (
            .O(N__54842),
            .I(N__54774));
    InMux I__13394 (
            .O(N__54841),
            .I(N__54771));
    InMux I__13393 (
            .O(N__54840),
            .I(N__54766));
    InMux I__13392 (
            .O(N__54839),
            .I(N__54766));
    LocalMux I__13391 (
            .O(N__54836),
            .I(N__54761));
    LocalMux I__13390 (
            .O(N__54833),
            .I(N__54761));
    Span4Mux_v I__13389 (
            .O(N__54828),
            .I(N__54758));
    InMux I__13388 (
            .O(N__54827),
            .I(N__54755));
    InMux I__13387 (
            .O(N__54826),
            .I(N__54750));
    InMux I__13386 (
            .O(N__54825),
            .I(N__54747));
    LocalMux I__13385 (
            .O(N__54822),
            .I(N__54744));
    LocalMux I__13384 (
            .O(N__54811),
            .I(N__54741));
    CascadeMux I__13383 (
            .O(N__54810),
            .I(N__54734));
    LocalMux I__13382 (
            .O(N__54807),
            .I(N__54731));
    Span4Mux_v I__13381 (
            .O(N__54804),
            .I(N__54728));
    InMux I__13380 (
            .O(N__54803),
            .I(N__54725));
    InMux I__13379 (
            .O(N__54800),
            .I(N__54716));
    InMux I__13378 (
            .O(N__54797),
            .I(N__54716));
    InMux I__13377 (
            .O(N__54796),
            .I(N__54716));
    InMux I__13376 (
            .O(N__54795),
            .I(N__54716));
    LocalMux I__13375 (
            .O(N__54792),
            .I(N__54711));
    Span4Mux_h I__13374 (
            .O(N__54789),
            .I(N__54711));
    CascadeMux I__13373 (
            .O(N__54788),
            .I(N__54707));
    InMux I__13372 (
            .O(N__54787),
            .I(N__54703));
    LocalMux I__13371 (
            .O(N__54784),
            .I(N__54696));
    Span4Mux_v I__13370 (
            .O(N__54781),
            .I(N__54696));
    LocalMux I__13369 (
            .O(N__54778),
            .I(N__54696));
    InMux I__13368 (
            .O(N__54777),
            .I(N__54691));
    InMux I__13367 (
            .O(N__54774),
            .I(N__54691));
    LocalMux I__13366 (
            .O(N__54771),
            .I(N__54686));
    LocalMux I__13365 (
            .O(N__54766),
            .I(N__54686));
    Span4Mux_v I__13364 (
            .O(N__54761),
            .I(N__54680));
    Span4Mux_h I__13363 (
            .O(N__54758),
            .I(N__54675));
    LocalMux I__13362 (
            .O(N__54755),
            .I(N__54675));
    InMux I__13361 (
            .O(N__54754),
            .I(N__54670));
    InMux I__13360 (
            .O(N__54753),
            .I(N__54670));
    LocalMux I__13359 (
            .O(N__54750),
            .I(N__54667));
    LocalMux I__13358 (
            .O(N__54747),
            .I(N__54662));
    Span4Mux_v I__13357 (
            .O(N__54744),
            .I(N__54662));
    Span4Mux_h I__13356 (
            .O(N__54741),
            .I(N__54659));
    InMux I__13355 (
            .O(N__54740),
            .I(N__54652));
    InMux I__13354 (
            .O(N__54739),
            .I(N__54652));
    InMux I__13353 (
            .O(N__54738),
            .I(N__54652));
    InMux I__13352 (
            .O(N__54737),
            .I(N__54649));
    InMux I__13351 (
            .O(N__54734),
            .I(N__54646));
    Span12Mux_h I__13350 (
            .O(N__54731),
            .I(N__54643));
    Span4Mux_h I__13349 (
            .O(N__54728),
            .I(N__54640));
    LocalMux I__13348 (
            .O(N__54725),
            .I(N__54633));
    LocalMux I__13347 (
            .O(N__54716),
            .I(N__54633));
    Span4Mux_h I__13346 (
            .O(N__54711),
            .I(N__54633));
    InMux I__13345 (
            .O(N__54710),
            .I(N__54626));
    InMux I__13344 (
            .O(N__54707),
            .I(N__54626));
    InMux I__13343 (
            .O(N__54706),
            .I(N__54626));
    LocalMux I__13342 (
            .O(N__54703),
            .I(N__54617));
    Span4Mux_v I__13341 (
            .O(N__54696),
            .I(N__54617));
    LocalMux I__13340 (
            .O(N__54691),
            .I(N__54617));
    Span4Mux_v I__13339 (
            .O(N__54686),
            .I(N__54617));
    InMux I__13338 (
            .O(N__54685),
            .I(N__54610));
    InMux I__13337 (
            .O(N__54684),
            .I(N__54610));
    InMux I__13336 (
            .O(N__54683),
            .I(N__54610));
    Span4Mux_h I__13335 (
            .O(N__54680),
            .I(N__54603));
    Span4Mux_v I__13334 (
            .O(N__54675),
            .I(N__54603));
    LocalMux I__13333 (
            .O(N__54670),
            .I(N__54603));
    Span4Mux_v I__13332 (
            .O(N__54667),
            .I(N__54594));
    Span4Mux_h I__13331 (
            .O(N__54662),
            .I(N__54594));
    Span4Mux_v I__13330 (
            .O(N__54659),
            .I(N__54594));
    LocalMux I__13329 (
            .O(N__54652),
            .I(N__54594));
    LocalMux I__13328 (
            .O(N__54649),
            .I(comm_state_2));
    LocalMux I__13327 (
            .O(N__54646),
            .I(comm_state_2));
    Odrv12 I__13326 (
            .O(N__54643),
            .I(comm_state_2));
    Odrv4 I__13325 (
            .O(N__54640),
            .I(comm_state_2));
    Odrv4 I__13324 (
            .O(N__54633),
            .I(comm_state_2));
    LocalMux I__13323 (
            .O(N__54626),
            .I(comm_state_2));
    Odrv4 I__13322 (
            .O(N__54617),
            .I(comm_state_2));
    LocalMux I__13321 (
            .O(N__54610),
            .I(comm_state_2));
    Odrv4 I__13320 (
            .O(N__54603),
            .I(comm_state_2));
    Odrv4 I__13319 (
            .O(N__54594),
            .I(comm_state_2));
    InMux I__13318 (
            .O(N__54573),
            .I(N__54568));
    InMux I__13317 (
            .O(N__54572),
            .I(N__54563));
    InMux I__13316 (
            .O(N__54571),
            .I(N__54560));
    LocalMux I__13315 (
            .O(N__54568),
            .I(N__54557));
    InMux I__13314 (
            .O(N__54567),
            .I(N__54538));
    InMux I__13313 (
            .O(N__54566),
            .I(N__54535));
    LocalMux I__13312 (
            .O(N__54563),
            .I(N__54531));
    LocalMux I__13311 (
            .O(N__54560),
            .I(N__54526));
    Span4Mux_v I__13310 (
            .O(N__54557),
            .I(N__54526));
    InMux I__13309 (
            .O(N__54556),
            .I(N__54522));
    InMux I__13308 (
            .O(N__54555),
            .I(N__54519));
    InMux I__13307 (
            .O(N__54554),
            .I(N__54511));
    InMux I__13306 (
            .O(N__54553),
            .I(N__54495));
    CascadeMux I__13305 (
            .O(N__54552),
            .I(N__54491));
    InMux I__13304 (
            .O(N__54551),
            .I(N__54467));
    InMux I__13303 (
            .O(N__54550),
            .I(N__54467));
    InMux I__13302 (
            .O(N__54549),
            .I(N__54467));
    InMux I__13301 (
            .O(N__54548),
            .I(N__54467));
    InMux I__13300 (
            .O(N__54547),
            .I(N__54467));
    InMux I__13299 (
            .O(N__54546),
            .I(N__54467));
    InMux I__13298 (
            .O(N__54545),
            .I(N__54467));
    InMux I__13297 (
            .O(N__54544),
            .I(N__54467));
    InMux I__13296 (
            .O(N__54543),
            .I(N__54464));
    InMux I__13295 (
            .O(N__54542),
            .I(N__54461));
    InMux I__13294 (
            .O(N__54541),
            .I(N__54458));
    LocalMux I__13293 (
            .O(N__54538),
            .I(N__54455));
    LocalMux I__13292 (
            .O(N__54535),
            .I(N__54452));
    InMux I__13291 (
            .O(N__54534),
            .I(N__54449));
    Span4Mux_h I__13290 (
            .O(N__54531),
            .I(N__54444));
    Span4Mux_h I__13289 (
            .O(N__54526),
            .I(N__54444));
    InMux I__13288 (
            .O(N__54525),
            .I(N__54441));
    LocalMux I__13287 (
            .O(N__54522),
            .I(N__54426));
    LocalMux I__13286 (
            .O(N__54519),
            .I(N__54423));
    InMux I__13285 (
            .O(N__54518),
            .I(N__54418));
    InMux I__13284 (
            .O(N__54517),
            .I(N__54418));
    InMux I__13283 (
            .O(N__54516),
            .I(N__54414));
    CascadeMux I__13282 (
            .O(N__54515),
            .I(N__54411));
    InMux I__13281 (
            .O(N__54514),
            .I(N__54406));
    LocalMux I__13280 (
            .O(N__54511),
            .I(N__54403));
    InMux I__13279 (
            .O(N__54510),
            .I(N__54397));
    InMux I__13278 (
            .O(N__54509),
            .I(N__54390));
    InMux I__13277 (
            .O(N__54508),
            .I(N__54390));
    InMux I__13276 (
            .O(N__54507),
            .I(N__54390));
    InMux I__13275 (
            .O(N__54506),
            .I(N__54381));
    InMux I__13274 (
            .O(N__54505),
            .I(N__54381));
    InMux I__13273 (
            .O(N__54504),
            .I(N__54381));
    InMux I__13272 (
            .O(N__54503),
            .I(N__54381));
    CascadeMux I__13271 (
            .O(N__54502),
            .I(N__54376));
    InMux I__13270 (
            .O(N__54501),
            .I(N__54371));
    InMux I__13269 (
            .O(N__54500),
            .I(N__54368));
    InMux I__13268 (
            .O(N__54499),
            .I(N__54363));
    InMux I__13267 (
            .O(N__54498),
            .I(N__54360));
    LocalMux I__13266 (
            .O(N__54495),
            .I(N__54357));
    InMux I__13265 (
            .O(N__54494),
            .I(N__54350));
    InMux I__13264 (
            .O(N__54491),
            .I(N__54350));
    InMux I__13263 (
            .O(N__54490),
            .I(N__54350));
    InMux I__13262 (
            .O(N__54489),
            .I(N__54343));
    InMux I__13261 (
            .O(N__54488),
            .I(N__54343));
    InMux I__13260 (
            .O(N__54487),
            .I(N__54343));
    InMux I__13259 (
            .O(N__54486),
            .I(N__54326));
    InMux I__13258 (
            .O(N__54485),
            .I(N__54326));
    InMux I__13257 (
            .O(N__54484),
            .I(N__54323));
    LocalMux I__13256 (
            .O(N__54467),
            .I(N__54308));
    LocalMux I__13255 (
            .O(N__54464),
            .I(N__54308));
    LocalMux I__13254 (
            .O(N__54461),
            .I(N__54308));
    LocalMux I__13253 (
            .O(N__54458),
            .I(N__54308));
    Span4Mux_h I__13252 (
            .O(N__54455),
            .I(N__54308));
    Span4Mux_v I__13251 (
            .O(N__54452),
            .I(N__54308));
    LocalMux I__13250 (
            .O(N__54449),
            .I(N__54308));
    Span4Mux_h I__13249 (
            .O(N__54444),
            .I(N__54303));
    LocalMux I__13248 (
            .O(N__54441),
            .I(N__54303));
    InMux I__13247 (
            .O(N__54440),
            .I(N__54300));
    InMux I__13246 (
            .O(N__54439),
            .I(N__54293));
    InMux I__13245 (
            .O(N__54438),
            .I(N__54293));
    InMux I__13244 (
            .O(N__54437),
            .I(N__54293));
    InMux I__13243 (
            .O(N__54436),
            .I(N__54276));
    InMux I__13242 (
            .O(N__54435),
            .I(N__54276));
    InMux I__13241 (
            .O(N__54434),
            .I(N__54276));
    InMux I__13240 (
            .O(N__54433),
            .I(N__54276));
    InMux I__13239 (
            .O(N__54432),
            .I(N__54276));
    InMux I__13238 (
            .O(N__54431),
            .I(N__54276));
    InMux I__13237 (
            .O(N__54430),
            .I(N__54276));
    InMux I__13236 (
            .O(N__54429),
            .I(N__54276));
    Span4Mux_v I__13235 (
            .O(N__54426),
            .I(N__54269));
    Span4Mux_h I__13234 (
            .O(N__54423),
            .I(N__54269));
    LocalMux I__13233 (
            .O(N__54418),
            .I(N__54269));
    InMux I__13232 (
            .O(N__54417),
            .I(N__54266));
    LocalMux I__13231 (
            .O(N__54414),
            .I(N__54263));
    InMux I__13230 (
            .O(N__54411),
            .I(N__54256));
    InMux I__13229 (
            .O(N__54410),
            .I(N__54256));
    InMux I__13228 (
            .O(N__54409),
            .I(N__54256));
    LocalMux I__13227 (
            .O(N__54406),
            .I(N__54251));
    Span4Mux_v I__13226 (
            .O(N__54403),
            .I(N__54251));
    InMux I__13225 (
            .O(N__54402),
            .I(N__54248));
    InMux I__13224 (
            .O(N__54401),
            .I(N__54245));
    InMux I__13223 (
            .O(N__54400),
            .I(N__54242));
    LocalMux I__13222 (
            .O(N__54397),
            .I(N__54235));
    LocalMux I__13221 (
            .O(N__54390),
            .I(N__54235));
    LocalMux I__13220 (
            .O(N__54381),
            .I(N__54235));
    InMux I__13219 (
            .O(N__54380),
            .I(N__54232));
    InMux I__13218 (
            .O(N__54379),
            .I(N__54225));
    InMux I__13217 (
            .O(N__54376),
            .I(N__54225));
    InMux I__13216 (
            .O(N__54375),
            .I(N__54225));
    InMux I__13215 (
            .O(N__54374),
            .I(N__54222));
    LocalMux I__13214 (
            .O(N__54371),
            .I(N__54217));
    LocalMux I__13213 (
            .O(N__54368),
            .I(N__54217));
    InMux I__13212 (
            .O(N__54367),
            .I(N__54212));
    InMux I__13211 (
            .O(N__54366),
            .I(N__54212));
    LocalMux I__13210 (
            .O(N__54363),
            .I(N__54201));
    LocalMux I__13209 (
            .O(N__54360),
            .I(N__54201));
    Span4Mux_v I__13208 (
            .O(N__54357),
            .I(N__54201));
    LocalMux I__13207 (
            .O(N__54350),
            .I(N__54201));
    LocalMux I__13206 (
            .O(N__54343),
            .I(N__54201));
    InMux I__13205 (
            .O(N__54342),
            .I(N__54188));
    InMux I__13204 (
            .O(N__54341),
            .I(N__54185));
    CascadeMux I__13203 (
            .O(N__54340),
            .I(N__54180));
    CascadeMux I__13202 (
            .O(N__54339),
            .I(N__54174));
    InMux I__13201 (
            .O(N__54338),
            .I(N__54155));
    InMux I__13200 (
            .O(N__54337),
            .I(N__54155));
    InMux I__13199 (
            .O(N__54336),
            .I(N__54155));
    InMux I__13198 (
            .O(N__54335),
            .I(N__54155));
    InMux I__13197 (
            .O(N__54334),
            .I(N__54155));
    InMux I__13196 (
            .O(N__54333),
            .I(N__54155));
    InMux I__13195 (
            .O(N__54332),
            .I(N__54155));
    InMux I__13194 (
            .O(N__54331),
            .I(N__54155));
    LocalMux I__13193 (
            .O(N__54326),
            .I(N__54152));
    LocalMux I__13192 (
            .O(N__54323),
            .I(N__54141));
    Span4Mux_v I__13191 (
            .O(N__54308),
            .I(N__54141));
    Span4Mux_h I__13190 (
            .O(N__54303),
            .I(N__54141));
    LocalMux I__13189 (
            .O(N__54300),
            .I(N__54141));
    LocalMux I__13188 (
            .O(N__54293),
            .I(N__54141));
    LocalMux I__13187 (
            .O(N__54276),
            .I(N__54136));
    Span4Mux_h I__13186 (
            .O(N__54269),
            .I(N__54136));
    LocalMux I__13185 (
            .O(N__54266),
            .I(N__54129));
    Span4Mux_v I__13184 (
            .O(N__54263),
            .I(N__54129));
    LocalMux I__13183 (
            .O(N__54256),
            .I(N__54129));
    Sp12to4 I__13182 (
            .O(N__54251),
            .I(N__54126));
    LocalMux I__13181 (
            .O(N__54248),
            .I(N__54115));
    LocalMux I__13180 (
            .O(N__54245),
            .I(N__54115));
    LocalMux I__13179 (
            .O(N__54242),
            .I(N__54115));
    Sp12to4 I__13178 (
            .O(N__54235),
            .I(N__54115));
    LocalMux I__13177 (
            .O(N__54232),
            .I(N__54115));
    LocalMux I__13176 (
            .O(N__54225),
            .I(N__54112));
    LocalMux I__13175 (
            .O(N__54222),
            .I(N__54103));
    Span4Mux_h I__13174 (
            .O(N__54217),
            .I(N__54103));
    LocalMux I__13173 (
            .O(N__54212),
            .I(N__54103));
    Span4Mux_v I__13172 (
            .O(N__54201),
            .I(N__54103));
    InMux I__13171 (
            .O(N__54200),
            .I(N__54086));
    InMux I__13170 (
            .O(N__54199),
            .I(N__54086));
    InMux I__13169 (
            .O(N__54198),
            .I(N__54086));
    InMux I__13168 (
            .O(N__54197),
            .I(N__54086));
    InMux I__13167 (
            .O(N__54196),
            .I(N__54086));
    InMux I__13166 (
            .O(N__54195),
            .I(N__54086));
    InMux I__13165 (
            .O(N__54194),
            .I(N__54086));
    InMux I__13164 (
            .O(N__54193),
            .I(N__54086));
    InMux I__13163 (
            .O(N__54192),
            .I(N__54081));
    InMux I__13162 (
            .O(N__54191),
            .I(N__54081));
    LocalMux I__13161 (
            .O(N__54188),
            .I(N__54078));
    LocalMux I__13160 (
            .O(N__54185),
            .I(N__54075));
    InMux I__13159 (
            .O(N__54184),
            .I(N__54068));
    InMux I__13158 (
            .O(N__54183),
            .I(N__54068));
    InMux I__13157 (
            .O(N__54180),
            .I(N__54068));
    InMux I__13156 (
            .O(N__54179),
            .I(N__54063));
    InMux I__13155 (
            .O(N__54178),
            .I(N__54063));
    InMux I__13154 (
            .O(N__54177),
            .I(N__54054));
    InMux I__13153 (
            .O(N__54174),
            .I(N__54054));
    InMux I__13152 (
            .O(N__54173),
            .I(N__54054));
    InMux I__13151 (
            .O(N__54172),
            .I(N__54054));
    LocalMux I__13150 (
            .O(N__54155),
            .I(N__54047));
    Span4Mux_v I__13149 (
            .O(N__54152),
            .I(N__54047));
    Span4Mux_v I__13148 (
            .O(N__54141),
            .I(N__54047));
    Span4Mux_h I__13147 (
            .O(N__54136),
            .I(N__54042));
    Span4Mux_v I__13146 (
            .O(N__54129),
            .I(N__54042));
    Span12Mux_h I__13145 (
            .O(N__54126),
            .I(N__54037));
    Span12Mux_v I__13144 (
            .O(N__54115),
            .I(N__54037));
    Span4Mux_h I__13143 (
            .O(N__54112),
            .I(N__54032));
    Span4Mux_h I__13142 (
            .O(N__54103),
            .I(N__54032));
    LocalMux I__13141 (
            .O(N__54086),
            .I(comm_state_1));
    LocalMux I__13140 (
            .O(N__54081),
            .I(comm_state_1));
    Odrv12 I__13139 (
            .O(N__54078),
            .I(comm_state_1));
    Odrv12 I__13138 (
            .O(N__54075),
            .I(comm_state_1));
    LocalMux I__13137 (
            .O(N__54068),
            .I(comm_state_1));
    LocalMux I__13136 (
            .O(N__54063),
            .I(comm_state_1));
    LocalMux I__13135 (
            .O(N__54054),
            .I(comm_state_1));
    Odrv4 I__13134 (
            .O(N__54047),
            .I(comm_state_1));
    Odrv4 I__13133 (
            .O(N__54042),
            .I(comm_state_1));
    Odrv12 I__13132 (
            .O(N__54037),
            .I(comm_state_1));
    Odrv4 I__13131 (
            .O(N__54032),
            .I(comm_state_1));
    InMux I__13130 (
            .O(N__54009),
            .I(N__53998));
    InMux I__13129 (
            .O(N__54008),
            .I(N__53994));
    InMux I__13128 (
            .O(N__54007),
            .I(N__53989));
    InMux I__13127 (
            .O(N__54006),
            .I(N__53989));
    CascadeMux I__13126 (
            .O(N__54005),
            .I(N__53983));
    InMux I__13125 (
            .O(N__54004),
            .I(N__53970));
    InMux I__13124 (
            .O(N__54003),
            .I(N__53970));
    InMux I__13123 (
            .O(N__54002),
            .I(N__53970));
    InMux I__13122 (
            .O(N__54001),
            .I(N__53966));
    LocalMux I__13121 (
            .O(N__53998),
            .I(N__53959));
    InMux I__13120 (
            .O(N__53997),
            .I(N__53956));
    LocalMux I__13119 (
            .O(N__53994),
            .I(N__53951));
    LocalMux I__13118 (
            .O(N__53989),
            .I(N__53951));
    InMux I__13117 (
            .O(N__53988),
            .I(N__53948));
    InMux I__13116 (
            .O(N__53987),
            .I(N__53943));
    CascadeMux I__13115 (
            .O(N__53986),
            .I(N__53940));
    InMux I__13114 (
            .O(N__53983),
            .I(N__53931));
    InMux I__13113 (
            .O(N__53982),
            .I(N__53931));
    InMux I__13112 (
            .O(N__53981),
            .I(N__53931));
    InMux I__13111 (
            .O(N__53980),
            .I(N__53931));
    InMux I__13110 (
            .O(N__53979),
            .I(N__53924));
    InMux I__13109 (
            .O(N__53978),
            .I(N__53924));
    InMux I__13108 (
            .O(N__53977),
            .I(N__53924));
    LocalMux I__13107 (
            .O(N__53970),
            .I(N__53916));
    InMux I__13106 (
            .O(N__53969),
            .I(N__53913));
    LocalMux I__13105 (
            .O(N__53966),
            .I(N__53910));
    InMux I__13104 (
            .O(N__53965),
            .I(N__53905));
    InMux I__13103 (
            .O(N__53964),
            .I(N__53905));
    InMux I__13102 (
            .O(N__53963),
            .I(N__53900));
    InMux I__13101 (
            .O(N__53962),
            .I(N__53900));
    Span4Mux_v I__13100 (
            .O(N__53959),
            .I(N__53897));
    LocalMux I__13099 (
            .O(N__53956),
            .I(N__53894));
    Span4Mux_h I__13098 (
            .O(N__53951),
            .I(N__53889));
    LocalMux I__13097 (
            .O(N__53948),
            .I(N__53889));
    InMux I__13096 (
            .O(N__53947),
            .I(N__53886));
    InMux I__13095 (
            .O(N__53946),
            .I(N__53883));
    LocalMux I__13094 (
            .O(N__53943),
            .I(N__53880));
    InMux I__13093 (
            .O(N__53940),
            .I(N__53877));
    LocalMux I__13092 (
            .O(N__53931),
            .I(N__53874));
    LocalMux I__13091 (
            .O(N__53924),
            .I(N__53865));
    InMux I__13090 (
            .O(N__53923),
            .I(N__53860));
    InMux I__13089 (
            .O(N__53922),
            .I(N__53860));
    InMux I__13088 (
            .O(N__53921),
            .I(N__53853));
    InMux I__13087 (
            .O(N__53920),
            .I(N__53853));
    InMux I__13086 (
            .O(N__53919),
            .I(N__53853));
    Span4Mux_v I__13085 (
            .O(N__53916),
            .I(N__53850));
    LocalMux I__13084 (
            .O(N__53913),
            .I(N__53845));
    Span4Mux_v I__13083 (
            .O(N__53910),
            .I(N__53845));
    LocalMux I__13082 (
            .O(N__53905),
            .I(N__53838));
    LocalMux I__13081 (
            .O(N__53900),
            .I(N__53838));
    Span4Mux_h I__13080 (
            .O(N__53897),
            .I(N__53838));
    Span4Mux_v I__13079 (
            .O(N__53894),
            .I(N__53833));
    Span4Mux_v I__13078 (
            .O(N__53889),
            .I(N__53833));
    LocalMux I__13077 (
            .O(N__53886),
            .I(N__53830));
    LocalMux I__13076 (
            .O(N__53883),
            .I(N__53823));
    Span4Mux_v I__13075 (
            .O(N__53880),
            .I(N__53823));
    LocalMux I__13074 (
            .O(N__53877),
            .I(N__53823));
    Span4Mux_v I__13073 (
            .O(N__53874),
            .I(N__53820));
    InMux I__13072 (
            .O(N__53873),
            .I(N__53811));
    InMux I__13071 (
            .O(N__53872),
            .I(N__53811));
    InMux I__13070 (
            .O(N__53871),
            .I(N__53811));
    InMux I__13069 (
            .O(N__53870),
            .I(N__53811));
    InMux I__13068 (
            .O(N__53869),
            .I(N__53806));
    InMux I__13067 (
            .O(N__53868),
            .I(N__53806));
    Span4Mux_v I__13066 (
            .O(N__53865),
            .I(N__53793));
    LocalMux I__13065 (
            .O(N__53860),
            .I(N__53793));
    LocalMux I__13064 (
            .O(N__53853),
            .I(N__53793));
    Span4Mux_v I__13063 (
            .O(N__53850),
            .I(N__53793));
    Span4Mux_h I__13062 (
            .O(N__53845),
            .I(N__53793));
    Span4Mux_v I__13061 (
            .O(N__53838),
            .I(N__53793));
    Span4Mux_h I__13060 (
            .O(N__53833),
            .I(N__53790));
    Odrv12 I__13059 (
            .O(N__53830),
            .I(comm_state_0));
    Odrv4 I__13058 (
            .O(N__53823),
            .I(comm_state_0));
    Odrv4 I__13057 (
            .O(N__53820),
            .I(comm_state_0));
    LocalMux I__13056 (
            .O(N__53811),
            .I(comm_state_0));
    LocalMux I__13055 (
            .O(N__53806),
            .I(comm_state_0));
    Odrv4 I__13054 (
            .O(N__53793),
            .I(comm_state_0));
    Odrv4 I__13053 (
            .O(N__53790),
            .I(comm_state_0));
    InMux I__13052 (
            .O(N__53775),
            .I(N__53772));
    LocalMux I__13051 (
            .O(N__53772),
            .I(N__53769));
    Span4Mux_v I__13050 (
            .O(N__53769),
            .I(N__53766));
    Span4Mux_h I__13049 (
            .O(N__53766),
            .I(N__53763));
    Odrv4 I__13048 (
            .O(N__53763),
            .I(n10804));
    InMux I__13047 (
            .O(N__53760),
            .I(N__53757));
    LocalMux I__13046 (
            .O(N__53757),
            .I(N__53753));
    InMux I__13045 (
            .O(N__53756),
            .I(N__53750));
    Span4Mux_h I__13044 (
            .O(N__53753),
            .I(N__53747));
    LocalMux I__13043 (
            .O(N__53750),
            .I(\ADC_VDC.genclk.t0off_12 ));
    Odrv4 I__13042 (
            .O(N__53747),
            .I(\ADC_VDC.genclk.t0off_12 ));
    CascadeMux I__13041 (
            .O(N__53742),
            .I(N__53738));
    InMux I__13040 (
            .O(N__53741),
            .I(N__53735));
    InMux I__13039 (
            .O(N__53738),
            .I(N__53732));
    LocalMux I__13038 (
            .O(N__53735),
            .I(\ADC_VDC.genclk.t0off_2 ));
    LocalMux I__13037 (
            .O(N__53732),
            .I(\ADC_VDC.genclk.t0off_2 ));
    CascadeMux I__13036 (
            .O(N__53727),
            .I(N__53723));
    InMux I__13035 (
            .O(N__53726),
            .I(N__53720));
    InMux I__13034 (
            .O(N__53723),
            .I(N__53717));
    LocalMux I__13033 (
            .O(N__53720),
            .I(\ADC_VDC.genclk.t0off_7 ));
    LocalMux I__13032 (
            .O(N__53717),
            .I(\ADC_VDC.genclk.t0off_7 ));
    InMux I__13031 (
            .O(N__53712),
            .I(N__53708));
    InMux I__13030 (
            .O(N__53711),
            .I(N__53705));
    LocalMux I__13029 (
            .O(N__53708),
            .I(N__53702));
    LocalMux I__13028 (
            .O(N__53705),
            .I(\ADC_VDC.genclk.t0off_10 ));
    Odrv4 I__13027 (
            .O(N__53702),
            .I(\ADC_VDC.genclk.t0off_10 ));
    CascadeMux I__13026 (
            .O(N__53697),
            .I(\ADC_VDC.genclk.n27_cascade_ ));
    CascadeMux I__13025 (
            .O(N__53694),
            .I(\ADC_VDC.genclk.n21598_cascade_ ));
    CEMux I__13024 (
            .O(N__53691),
            .I(N__53688));
    LocalMux I__13023 (
            .O(N__53688),
            .I(\ADC_VDC.genclk.n6 ));
    InMux I__13022 (
            .O(N__53685),
            .I(N__53682));
    LocalMux I__13021 (
            .O(N__53682),
            .I(N__53679));
    Span4Mux_h I__13020 (
            .O(N__53679),
            .I(N__53676));
    Span4Mux_h I__13019 (
            .O(N__53676),
            .I(N__53671));
    InMux I__13018 (
            .O(N__53675),
            .I(N__53666));
    InMux I__13017 (
            .O(N__53674),
            .I(N__53666));
    Span4Mux_v I__13016 (
            .O(N__53671),
            .I(N__53663));
    LocalMux I__13015 (
            .O(N__53666),
            .I(N__53660));
    Odrv4 I__13014 (
            .O(N__53663),
            .I(comm_tx_buf_5));
    Odrv4 I__13013 (
            .O(N__53660),
            .I(comm_tx_buf_5));
    SRMux I__13012 (
            .O(N__53655),
            .I(N__53652));
    LocalMux I__13011 (
            .O(N__53652),
            .I(\comm_spi.data_tx_7__N_808 ));
    InMux I__13010 (
            .O(N__53649),
            .I(N__53646));
    LocalMux I__13009 (
            .O(N__53646),
            .I(N__53641));
    InMux I__13008 (
            .O(N__53645),
            .I(N__53637));
    InMux I__13007 (
            .O(N__53644),
            .I(N__53633));
    Span4Mux_h I__13006 (
            .O(N__53641),
            .I(N__53630));
    InMux I__13005 (
            .O(N__53640),
            .I(N__53627));
    LocalMux I__13004 (
            .O(N__53637),
            .I(N__53624));
    InMux I__13003 (
            .O(N__53636),
            .I(N__53621));
    LocalMux I__13002 (
            .O(N__53633),
            .I(N__53612));
    Span4Mux_h I__13001 (
            .O(N__53630),
            .I(N__53612));
    LocalMux I__13000 (
            .O(N__53627),
            .I(N__53612));
    Span4Mux_v I__12999 (
            .O(N__53624),
            .I(N__53607));
    LocalMux I__12998 (
            .O(N__53621),
            .I(N__53607));
    InMux I__12997 (
            .O(N__53620),
            .I(N__53604));
    InMux I__12996 (
            .O(N__53619),
            .I(N__53601));
    Span4Mux_v I__12995 (
            .O(N__53612),
            .I(N__53597));
    Span4Mux_v I__12994 (
            .O(N__53607),
            .I(N__53594));
    LocalMux I__12993 (
            .O(N__53604),
            .I(N__53591));
    LocalMux I__12992 (
            .O(N__53601),
            .I(N__53588));
    InMux I__12991 (
            .O(N__53600),
            .I(N__53585));
    Sp12to4 I__12990 (
            .O(N__53597),
            .I(N__53581));
    Span4Mux_h I__12989 (
            .O(N__53594),
            .I(N__53578));
    Span4Mux_h I__12988 (
            .O(N__53591),
            .I(N__53573));
    Span4Mux_h I__12987 (
            .O(N__53588),
            .I(N__53573));
    LocalMux I__12986 (
            .O(N__53585),
            .I(N__53570));
    InMux I__12985 (
            .O(N__53584),
            .I(N__53567));
    Odrv12 I__12984 (
            .O(N__53581),
            .I(comm_rx_buf_4));
    Odrv4 I__12983 (
            .O(N__53578),
            .I(comm_rx_buf_4));
    Odrv4 I__12982 (
            .O(N__53573),
            .I(comm_rx_buf_4));
    Odrv4 I__12981 (
            .O(N__53570),
            .I(comm_rx_buf_4));
    LocalMux I__12980 (
            .O(N__53567),
            .I(comm_rx_buf_4));
    InMux I__12979 (
            .O(N__53556),
            .I(N__53553));
    LocalMux I__12978 (
            .O(N__53553),
            .I(N__53549));
    InMux I__12977 (
            .O(N__53552),
            .I(N__53546));
    Span4Mux_h I__12976 (
            .O(N__53549),
            .I(N__53543));
    LocalMux I__12975 (
            .O(N__53546),
            .I(comm_buf_6_4));
    Odrv4 I__12974 (
            .O(N__53543),
            .I(comm_buf_6_4));
    InMux I__12973 (
            .O(N__53538),
            .I(N__53535));
    LocalMux I__12972 (
            .O(N__53535),
            .I(N__53532));
    Odrv4 I__12971 (
            .O(N__53532),
            .I(comm_buf_3_1));
    InMux I__12970 (
            .O(N__53529),
            .I(N__53526));
    LocalMux I__12969 (
            .O(N__53526),
            .I(N__53523));
    Span4Mux_h I__12968 (
            .O(N__53523),
            .I(N__53520));
    Odrv4 I__12967 (
            .O(N__53520),
            .I(comm_buf_2_1));
    InMux I__12966 (
            .O(N__53517),
            .I(N__53514));
    LocalMux I__12965 (
            .O(N__53514),
            .I(n2_adj_1587));
    InMux I__12964 (
            .O(N__53511),
            .I(N__53507));
    InMux I__12963 (
            .O(N__53510),
            .I(N__53504));
    LocalMux I__12962 (
            .O(N__53507),
            .I(N__53500));
    LocalMux I__12961 (
            .O(N__53504),
            .I(N__53496));
    InMux I__12960 (
            .O(N__53503),
            .I(N__53493));
    Span4Mux_v I__12959 (
            .O(N__53500),
            .I(N__53490));
    InMux I__12958 (
            .O(N__53499),
            .I(N__53487));
    Span4Mux_h I__12957 (
            .O(N__53496),
            .I(N__53482));
    LocalMux I__12956 (
            .O(N__53493),
            .I(N__53482));
    Sp12to4 I__12955 (
            .O(N__53490),
            .I(N__53477));
    LocalMux I__12954 (
            .O(N__53487),
            .I(N__53477));
    Span4Mux_h I__12953 (
            .O(N__53482),
            .I(N__53474));
    Span12Mux_s11_v I__12952 (
            .O(N__53477),
            .I(N__53471));
    Odrv4 I__12951 (
            .O(N__53474),
            .I(comm_buf_1_1));
    Odrv12 I__12950 (
            .O(N__53471),
            .I(comm_buf_1_1));
    CascadeMux I__12949 (
            .O(N__53466),
            .I(N__53463));
    InMux I__12948 (
            .O(N__53463),
            .I(N__53459));
    CascadeMux I__12947 (
            .O(N__53462),
            .I(N__53455));
    LocalMux I__12946 (
            .O(N__53459),
            .I(N__53452));
    CascadeMux I__12945 (
            .O(N__53458),
            .I(N__53449));
    InMux I__12944 (
            .O(N__53455),
            .I(N__53445));
    Span4Mux_h I__12943 (
            .O(N__53452),
            .I(N__53442));
    InMux I__12942 (
            .O(N__53449),
            .I(N__53439));
    InMux I__12941 (
            .O(N__53448),
            .I(N__53432));
    LocalMux I__12940 (
            .O(N__53445),
            .I(N__53425));
    Span4Mux_h I__12939 (
            .O(N__53442),
            .I(N__53425));
    LocalMux I__12938 (
            .O(N__53439),
            .I(N__53425));
    InMux I__12937 (
            .O(N__53438),
            .I(N__53418));
    InMux I__12936 (
            .O(N__53437),
            .I(N__53418));
    InMux I__12935 (
            .O(N__53436),
            .I(N__53415));
    InMux I__12934 (
            .O(N__53435),
            .I(N__53412));
    LocalMux I__12933 (
            .O(N__53432),
            .I(N__53407));
    Span4Mux_v I__12932 (
            .O(N__53425),
            .I(N__53407));
    InMux I__12931 (
            .O(N__53424),
            .I(N__53404));
    InMux I__12930 (
            .O(N__53423),
            .I(N__53401));
    LocalMux I__12929 (
            .O(N__53418),
            .I(N__53398));
    LocalMux I__12928 (
            .O(N__53415),
            .I(N__53393));
    LocalMux I__12927 (
            .O(N__53412),
            .I(N__53393));
    Span4Mux_h I__12926 (
            .O(N__53407),
            .I(N__53390));
    LocalMux I__12925 (
            .O(N__53404),
            .I(N__53387));
    LocalMux I__12924 (
            .O(N__53401),
            .I(N__53384));
    Span4Mux_h I__12923 (
            .O(N__53398),
            .I(N__53381));
    Span4Mux_v I__12922 (
            .O(N__53393),
            .I(N__53378));
    Span4Mux_h I__12921 (
            .O(N__53390),
            .I(N__53375));
    Span4Mux_v I__12920 (
            .O(N__53387),
            .I(N__53370));
    Span4Mux_v I__12919 (
            .O(N__53384),
            .I(N__53370));
    Span4Mux_v I__12918 (
            .O(N__53381),
            .I(N__53367));
    Odrv4 I__12917 (
            .O(N__53378),
            .I(comm_buf_0_1));
    Odrv4 I__12916 (
            .O(N__53375),
            .I(comm_buf_0_1));
    Odrv4 I__12915 (
            .O(N__53370),
            .I(comm_buf_0_1));
    Odrv4 I__12914 (
            .O(N__53367),
            .I(comm_buf_0_1));
    InMux I__12913 (
            .O(N__53358),
            .I(N__53355));
    LocalMux I__12912 (
            .O(N__53355),
            .I(N__53352));
    Odrv4 I__12911 (
            .O(N__53352),
            .I(n1_adj_1586));
    CascadeMux I__12910 (
            .O(N__53349),
            .I(N__53346));
    InMux I__12909 (
            .O(N__53346),
            .I(N__53339));
    CascadeMux I__12908 (
            .O(N__53345),
            .I(N__53336));
    CascadeMux I__12907 (
            .O(N__53344),
            .I(N__53333));
    InMux I__12906 (
            .O(N__53343),
            .I(N__53328));
    InMux I__12905 (
            .O(N__53342),
            .I(N__53325));
    LocalMux I__12904 (
            .O(N__53339),
            .I(N__53322));
    InMux I__12903 (
            .O(N__53336),
            .I(N__53319));
    InMux I__12902 (
            .O(N__53333),
            .I(N__53316));
    InMux I__12901 (
            .O(N__53332),
            .I(N__53313));
    InMux I__12900 (
            .O(N__53331),
            .I(N__53310));
    LocalMux I__12899 (
            .O(N__53328),
            .I(N__53305));
    LocalMux I__12898 (
            .O(N__53325),
            .I(N__53305));
    Span4Mux_h I__12897 (
            .O(N__53322),
            .I(N__53298));
    LocalMux I__12896 (
            .O(N__53319),
            .I(N__53298));
    LocalMux I__12895 (
            .O(N__53316),
            .I(N__53298));
    LocalMux I__12894 (
            .O(N__53313),
            .I(N__53293));
    LocalMux I__12893 (
            .O(N__53310),
            .I(N__53293));
    Span4Mux_v I__12892 (
            .O(N__53305),
            .I(N__53288));
    Span4Mux_v I__12891 (
            .O(N__53298),
            .I(N__53283));
    Span4Mux_v I__12890 (
            .O(N__53293),
            .I(N__53283));
    InMux I__12889 (
            .O(N__53292),
            .I(N__53280));
    InMux I__12888 (
            .O(N__53291),
            .I(N__53277));
    Odrv4 I__12887 (
            .O(N__53288),
            .I(comm_rx_buf_5));
    Odrv4 I__12886 (
            .O(N__53283),
            .I(comm_rx_buf_5));
    LocalMux I__12885 (
            .O(N__53280),
            .I(comm_rx_buf_5));
    LocalMux I__12884 (
            .O(N__53277),
            .I(comm_rx_buf_5));
    InMux I__12883 (
            .O(N__53268),
            .I(N__53264));
    InMux I__12882 (
            .O(N__53267),
            .I(N__53261));
    LocalMux I__12881 (
            .O(N__53264),
            .I(comm_buf_6_5));
    LocalMux I__12880 (
            .O(N__53261),
            .I(comm_buf_6_5));
    InMux I__12879 (
            .O(N__53256),
            .I(N__53253));
    LocalMux I__12878 (
            .O(N__53253),
            .I(N__53250));
    Span4Mux_h I__12877 (
            .O(N__53250),
            .I(N__53247));
    Odrv4 I__12876 (
            .O(N__53247),
            .I(buf_data_iac_14));
    InMux I__12875 (
            .O(N__53244),
            .I(N__53241));
    LocalMux I__12874 (
            .O(N__53241),
            .I(N__53238));
    Odrv4 I__12873 (
            .O(N__53238),
            .I(n21547));
    CascadeMux I__12872 (
            .O(N__53235),
            .I(N__53231));
    CascadeMux I__12871 (
            .O(N__53234),
            .I(N__53228));
    InMux I__12870 (
            .O(N__53231),
            .I(N__53222));
    InMux I__12869 (
            .O(N__53228),
            .I(N__53219));
    InMux I__12868 (
            .O(N__53227),
            .I(N__53214));
    InMux I__12867 (
            .O(N__53226),
            .I(N__53211));
    InMux I__12866 (
            .O(N__53225),
            .I(N__53208));
    LocalMux I__12865 (
            .O(N__53222),
            .I(N__53205));
    LocalMux I__12864 (
            .O(N__53219),
            .I(N__53202));
    InMux I__12863 (
            .O(N__53218),
            .I(N__53199));
    InMux I__12862 (
            .O(N__53217),
            .I(N__53196));
    LocalMux I__12861 (
            .O(N__53214),
            .I(N__53192));
    LocalMux I__12860 (
            .O(N__53211),
            .I(N__53189));
    LocalMux I__12859 (
            .O(N__53208),
            .I(N__53184));
    Span4Mux_h I__12858 (
            .O(N__53205),
            .I(N__53184));
    Span4Mux_v I__12857 (
            .O(N__53202),
            .I(N__53177));
    LocalMux I__12856 (
            .O(N__53199),
            .I(N__53177));
    LocalMux I__12855 (
            .O(N__53196),
            .I(N__53177));
    InMux I__12854 (
            .O(N__53195),
            .I(N__53174));
    Span4Mux_v I__12853 (
            .O(N__53192),
            .I(N__53171));
    Span4Mux_h I__12852 (
            .O(N__53189),
            .I(N__53166));
    Span4Mux_h I__12851 (
            .O(N__53184),
            .I(N__53166));
    Span4Mux_h I__12850 (
            .O(N__53177),
            .I(N__53161));
    LocalMux I__12849 (
            .O(N__53174),
            .I(N__53161));
    Sp12to4 I__12848 (
            .O(N__53171),
            .I(N__53157));
    Sp12to4 I__12847 (
            .O(N__53166),
            .I(N__53152));
    Sp12to4 I__12846 (
            .O(N__53161),
            .I(N__53152));
    InMux I__12845 (
            .O(N__53160),
            .I(N__53149));
    Odrv12 I__12844 (
            .O(N__53157),
            .I(comm_rx_buf_6));
    Odrv12 I__12843 (
            .O(N__53152),
            .I(comm_rx_buf_6));
    LocalMux I__12842 (
            .O(N__53149),
            .I(comm_rx_buf_6));
    InMux I__12841 (
            .O(N__53142),
            .I(N__53138));
    InMux I__12840 (
            .O(N__53141),
            .I(N__53135));
    LocalMux I__12839 (
            .O(N__53138),
            .I(N__53132));
    LocalMux I__12838 (
            .O(N__53135),
            .I(N__53123));
    Span4Mux_h I__12837 (
            .O(N__53132),
            .I(N__53120));
    InMux I__12836 (
            .O(N__53131),
            .I(N__53117));
    InMux I__12835 (
            .O(N__53130),
            .I(N__53114));
    InMux I__12834 (
            .O(N__53129),
            .I(N__53109));
    InMux I__12833 (
            .O(N__53128),
            .I(N__53109));
    InMux I__12832 (
            .O(N__53127),
            .I(N__53106));
    InMux I__12831 (
            .O(N__53126),
            .I(N__53103));
    Odrv12 I__12830 (
            .O(N__53123),
            .I(n12477));
    Odrv4 I__12829 (
            .O(N__53120),
            .I(n12477));
    LocalMux I__12828 (
            .O(N__53117),
            .I(n12477));
    LocalMux I__12827 (
            .O(N__53114),
            .I(n12477));
    LocalMux I__12826 (
            .O(N__53109),
            .I(n12477));
    LocalMux I__12825 (
            .O(N__53106),
            .I(n12477));
    LocalMux I__12824 (
            .O(N__53103),
            .I(n12477));
    CascadeMux I__12823 (
            .O(N__53088),
            .I(N__53084));
    InMux I__12822 (
            .O(N__53087),
            .I(N__53081));
    InMux I__12821 (
            .O(N__53084),
            .I(N__53078));
    LocalMux I__12820 (
            .O(N__53081),
            .I(comm_buf_6_6));
    LocalMux I__12819 (
            .O(N__53078),
            .I(comm_buf_6_6));
    InMux I__12818 (
            .O(N__53073),
            .I(N__53058));
    InMux I__12817 (
            .O(N__53072),
            .I(N__53053));
    InMux I__12816 (
            .O(N__53071),
            .I(N__53053));
    CascadeMux I__12815 (
            .O(N__53070),
            .I(N__53043));
    InMux I__12814 (
            .O(N__53069),
            .I(N__53037));
    InMux I__12813 (
            .O(N__53068),
            .I(N__53037));
    InMux I__12812 (
            .O(N__53067),
            .I(N__53034));
    InMux I__12811 (
            .O(N__53066),
            .I(N__53025));
    InMux I__12810 (
            .O(N__53065),
            .I(N__53014));
    InMux I__12809 (
            .O(N__53064),
            .I(N__53014));
    InMux I__12808 (
            .O(N__53063),
            .I(N__53014));
    InMux I__12807 (
            .O(N__53062),
            .I(N__53014));
    InMux I__12806 (
            .O(N__53061),
            .I(N__53014));
    LocalMux I__12805 (
            .O(N__53058),
            .I(N__53009));
    LocalMux I__12804 (
            .O(N__53053),
            .I(N__53009));
    InMux I__12803 (
            .O(N__53052),
            .I(N__53002));
    InMux I__12802 (
            .O(N__53051),
            .I(N__53002));
    InMux I__12801 (
            .O(N__53050),
            .I(N__53002));
    InMux I__12800 (
            .O(N__53049),
            .I(N__52993));
    InMux I__12799 (
            .O(N__53048),
            .I(N__52993));
    InMux I__12798 (
            .O(N__53047),
            .I(N__52993));
    InMux I__12797 (
            .O(N__53046),
            .I(N__52993));
    InMux I__12796 (
            .O(N__53043),
            .I(N__52983));
    InMux I__12795 (
            .O(N__53042),
            .I(N__52980));
    LocalMux I__12794 (
            .O(N__53037),
            .I(N__52975));
    LocalMux I__12793 (
            .O(N__53034),
            .I(N__52975));
    InMux I__12792 (
            .O(N__53033),
            .I(N__52966));
    InMux I__12791 (
            .O(N__53032),
            .I(N__52966));
    InMux I__12790 (
            .O(N__53031),
            .I(N__52966));
    InMux I__12789 (
            .O(N__53030),
            .I(N__52966));
    InMux I__12788 (
            .O(N__53029),
            .I(N__52963));
    InMux I__12787 (
            .O(N__53028),
            .I(N__52960));
    LocalMux I__12786 (
            .O(N__53025),
            .I(N__52951));
    LocalMux I__12785 (
            .O(N__53014),
            .I(N__52951));
    Span4Mux_v I__12784 (
            .O(N__53009),
            .I(N__52951));
    LocalMux I__12783 (
            .O(N__53002),
            .I(N__52951));
    LocalMux I__12782 (
            .O(N__52993),
            .I(N__52948));
    InMux I__12781 (
            .O(N__52992),
            .I(N__52939));
    InMux I__12780 (
            .O(N__52991),
            .I(N__52939));
    InMux I__12779 (
            .O(N__52990),
            .I(N__52939));
    InMux I__12778 (
            .O(N__52989),
            .I(N__52939));
    InMux I__12777 (
            .O(N__52988),
            .I(N__52933));
    InMux I__12776 (
            .O(N__52987),
            .I(N__52933));
    InMux I__12775 (
            .O(N__52986),
            .I(N__52930));
    LocalMux I__12774 (
            .O(N__52983),
            .I(N__52927));
    LocalMux I__12773 (
            .O(N__52980),
            .I(N__52920));
    Span4Mux_v I__12772 (
            .O(N__52975),
            .I(N__52920));
    LocalMux I__12771 (
            .O(N__52966),
            .I(N__52920));
    LocalMux I__12770 (
            .O(N__52963),
            .I(N__52915));
    LocalMux I__12769 (
            .O(N__52960),
            .I(N__52915));
    Span4Mux_v I__12768 (
            .O(N__52951),
            .I(N__52908));
    Span4Mux_h I__12767 (
            .O(N__52948),
            .I(N__52908));
    LocalMux I__12766 (
            .O(N__52939),
            .I(N__52908));
    InMux I__12765 (
            .O(N__52938),
            .I(N__52905));
    LocalMux I__12764 (
            .O(N__52933),
            .I(comm_index_0));
    LocalMux I__12763 (
            .O(N__52930),
            .I(comm_index_0));
    Odrv12 I__12762 (
            .O(N__52927),
            .I(comm_index_0));
    Odrv4 I__12761 (
            .O(N__52920),
            .I(comm_index_0));
    Odrv12 I__12760 (
            .O(N__52915),
            .I(comm_index_0));
    Odrv4 I__12759 (
            .O(N__52908),
            .I(comm_index_0));
    LocalMux I__12758 (
            .O(N__52905),
            .I(comm_index_0));
    InMux I__12757 (
            .O(N__52890),
            .I(N__52887));
    LocalMux I__12756 (
            .O(N__52887),
            .I(n8_adj_1456));
    InMux I__12755 (
            .O(N__52884),
            .I(N__52872));
    InMux I__12754 (
            .O(N__52883),
            .I(N__52872));
    InMux I__12753 (
            .O(N__52882),
            .I(N__52872));
    InMux I__12752 (
            .O(N__52881),
            .I(N__52869));
    InMux I__12751 (
            .O(N__52880),
            .I(N__52864));
    InMux I__12750 (
            .O(N__52879),
            .I(N__52864));
    LocalMux I__12749 (
            .O(N__52872),
            .I(N__52852));
    LocalMux I__12748 (
            .O(N__52869),
            .I(N__52849));
    LocalMux I__12747 (
            .O(N__52864),
            .I(N__52846));
    InMux I__12746 (
            .O(N__52863),
            .I(N__52839));
    InMux I__12745 (
            .O(N__52862),
            .I(N__52839));
    InMux I__12744 (
            .O(N__52861),
            .I(N__52839));
    InMux I__12743 (
            .O(N__52860),
            .I(N__52828));
    InMux I__12742 (
            .O(N__52859),
            .I(N__52828));
    InMux I__12741 (
            .O(N__52858),
            .I(N__52828));
    InMux I__12740 (
            .O(N__52857),
            .I(N__52828));
    InMux I__12739 (
            .O(N__52856),
            .I(N__52828));
    CascadeMux I__12738 (
            .O(N__52855),
            .I(N__52825));
    Span4Mux_v I__12737 (
            .O(N__52852),
            .I(N__52820));
    Span4Mux_v I__12736 (
            .O(N__52849),
            .I(N__52820));
    Span4Mux_v I__12735 (
            .O(N__52846),
            .I(N__52813));
    LocalMux I__12734 (
            .O(N__52839),
            .I(N__52813));
    LocalMux I__12733 (
            .O(N__52828),
            .I(N__52813));
    InMux I__12732 (
            .O(N__52825),
            .I(N__52810));
    Odrv4 I__12731 (
            .O(N__52820),
            .I(comm_data_vld));
    Odrv4 I__12730 (
            .O(N__52813),
            .I(comm_data_vld));
    LocalMux I__12729 (
            .O(N__52810),
            .I(comm_data_vld));
    CascadeMux I__12728 (
            .O(N__52803),
            .I(N__52800));
    InMux I__12727 (
            .O(N__52800),
            .I(N__52784));
    InMux I__12726 (
            .O(N__52799),
            .I(N__52784));
    InMux I__12725 (
            .O(N__52798),
            .I(N__52784));
    InMux I__12724 (
            .O(N__52797),
            .I(N__52784));
    CascadeMux I__12723 (
            .O(N__52796),
            .I(N__52778));
    CascadeMux I__12722 (
            .O(N__52795),
            .I(N__52775));
    CascadeMux I__12721 (
            .O(N__52794),
            .I(N__52772));
    CascadeMux I__12720 (
            .O(N__52793),
            .I(N__52764));
    LocalMux I__12719 (
            .O(N__52784),
            .I(N__52759));
    InMux I__12718 (
            .O(N__52783),
            .I(N__52756));
    InMux I__12717 (
            .O(N__52782),
            .I(N__52753));
    InMux I__12716 (
            .O(N__52781),
            .I(N__52750));
    InMux I__12715 (
            .O(N__52778),
            .I(N__52745));
    InMux I__12714 (
            .O(N__52775),
            .I(N__52745));
    InMux I__12713 (
            .O(N__52772),
            .I(N__52740));
    InMux I__12712 (
            .O(N__52771),
            .I(N__52740));
    InMux I__12711 (
            .O(N__52770),
            .I(N__52727));
    InMux I__12710 (
            .O(N__52769),
            .I(N__52727));
    InMux I__12709 (
            .O(N__52768),
            .I(N__52727));
    InMux I__12708 (
            .O(N__52767),
            .I(N__52727));
    InMux I__12707 (
            .O(N__52764),
            .I(N__52727));
    InMux I__12706 (
            .O(N__52763),
            .I(N__52727));
    InMux I__12705 (
            .O(N__52762),
            .I(N__52724));
    Span4Mux_h I__12704 (
            .O(N__52759),
            .I(N__52719));
    LocalMux I__12703 (
            .O(N__52756),
            .I(N__52719));
    LocalMux I__12702 (
            .O(N__52753),
            .I(N__52712));
    LocalMux I__12701 (
            .O(N__52750),
            .I(N__52712));
    LocalMux I__12700 (
            .O(N__52745),
            .I(N__52712));
    LocalMux I__12699 (
            .O(N__52740),
            .I(N__52707));
    LocalMux I__12698 (
            .O(N__52727),
            .I(N__52707));
    LocalMux I__12697 (
            .O(N__52724),
            .I(N__52704));
    Span4Mux_v I__12696 (
            .O(N__52719),
            .I(N__52701));
    Span4Mux_v I__12695 (
            .O(N__52712),
            .I(N__52698));
    Span4Mux_v I__12694 (
            .O(N__52707),
            .I(N__52695));
    Span4Mux_h I__12693 (
            .O(N__52704),
            .I(N__52692));
    Span4Mux_h I__12692 (
            .O(N__52701),
            .I(N__52685));
    Span4Mux_h I__12691 (
            .O(N__52698),
            .I(N__52685));
    Sp12to4 I__12690 (
            .O(N__52695),
            .I(N__52682));
    Span4Mux_v I__12689 (
            .O(N__52692),
            .I(N__52679));
    InMux I__12688 (
            .O(N__52691),
            .I(N__52674));
    InMux I__12687 (
            .O(N__52690),
            .I(N__52674));
    Sp12to4 I__12686 (
            .O(N__52685),
            .I(N__52669));
    Span12Mux_h I__12685 (
            .O(N__52682),
            .I(N__52669));
    Sp12to4 I__12684 (
            .O(N__52679),
            .I(N__52664));
    LocalMux I__12683 (
            .O(N__52674),
            .I(N__52664));
    Span12Mux_v I__12682 (
            .O(N__52669),
            .I(N__52661));
    Span12Mux_v I__12681 (
            .O(N__52664),
            .I(N__52658));
    Odrv12 I__12680 (
            .O(N__52661),
            .I(ICE_SPI_CE0));
    Odrv12 I__12679 (
            .O(N__52658),
            .I(ICE_SPI_CE0));
    InMux I__12678 (
            .O(N__52653),
            .I(N__52650));
    LocalMux I__12677 (
            .O(N__52650),
            .I(n6401));
    SRMux I__12676 (
            .O(N__52647),
            .I(N__52644));
    LocalMux I__12675 (
            .O(N__52644),
            .I(N__52641));
    Span4Mux_h I__12674 (
            .O(N__52641),
            .I(N__52638));
    Span4Mux_h I__12673 (
            .O(N__52638),
            .I(N__52635));
    Odrv4 I__12672 (
            .O(N__52635),
            .I(n16821));
    InMux I__12671 (
            .O(N__52632),
            .I(N__52628));
    InMux I__12670 (
            .O(N__52631),
            .I(N__52625));
    LocalMux I__12669 (
            .O(N__52628),
            .I(N__52622));
    LocalMux I__12668 (
            .O(N__52625),
            .I(N__52619));
    Span4Mux_h I__12667 (
            .O(N__52622),
            .I(N__52616));
    Span4Mux_h I__12666 (
            .O(N__52619),
            .I(N__52613));
    Span4Mux_h I__12665 (
            .O(N__52616),
            .I(N__52610));
    Span4Mux_h I__12664 (
            .O(N__52613),
            .I(N__52607));
    Odrv4 I__12663 (
            .O(N__52610),
            .I(\comm_spi.n14842 ));
    Odrv4 I__12662 (
            .O(N__52607),
            .I(\comm_spi.n14842 ));
    InMux I__12661 (
            .O(N__52602),
            .I(N__52599));
    LocalMux I__12660 (
            .O(N__52599),
            .I(N__52596));
    Span4Mux_h I__12659 (
            .O(N__52596),
            .I(N__52593));
    Odrv4 I__12658 (
            .O(N__52593),
            .I(buf_data_iac_18));
    InMux I__12657 (
            .O(N__52590),
            .I(N__52587));
    LocalMux I__12656 (
            .O(N__52587),
            .I(N__52584));
    Span4Mux_h I__12655 (
            .O(N__52584),
            .I(N__52581));
    Odrv4 I__12654 (
            .O(N__52581),
            .I(n21460));
    InMux I__12653 (
            .O(N__52578),
            .I(N__52575));
    LocalMux I__12652 (
            .O(N__52575),
            .I(N__52572));
    Span12Mux_s11_h I__12651 (
            .O(N__52572),
            .I(N__52569));
    Odrv12 I__12650 (
            .O(N__52569),
            .I(comm_buf_2_5));
    InMux I__12649 (
            .O(N__52566),
            .I(N__52546));
    InMux I__12648 (
            .O(N__52565),
            .I(N__52546));
    InMux I__12647 (
            .O(N__52564),
            .I(N__52546));
    InMux I__12646 (
            .O(N__52563),
            .I(N__52539));
    InMux I__12645 (
            .O(N__52562),
            .I(N__52539));
    InMux I__12644 (
            .O(N__52561),
            .I(N__52539));
    InMux I__12643 (
            .O(N__52560),
            .I(N__52532));
    InMux I__12642 (
            .O(N__52559),
            .I(N__52532));
    InMux I__12641 (
            .O(N__52558),
            .I(N__52532));
    InMux I__12640 (
            .O(N__52557),
            .I(N__52527));
    InMux I__12639 (
            .O(N__52556),
            .I(N__52527));
    InMux I__12638 (
            .O(N__52555),
            .I(N__52524));
    CascadeMux I__12637 (
            .O(N__52554),
            .I(N__52517));
    InMux I__12636 (
            .O(N__52553),
            .I(N__52514));
    LocalMux I__12635 (
            .O(N__52546),
            .I(N__52503));
    LocalMux I__12634 (
            .O(N__52539),
            .I(N__52503));
    LocalMux I__12633 (
            .O(N__52532),
            .I(N__52503));
    LocalMux I__12632 (
            .O(N__52527),
            .I(N__52503));
    LocalMux I__12631 (
            .O(N__52524),
            .I(N__52500));
    InMux I__12630 (
            .O(N__52523),
            .I(N__52495));
    InMux I__12629 (
            .O(N__52522),
            .I(N__52495));
    InMux I__12628 (
            .O(N__52521),
            .I(N__52490));
    InMux I__12627 (
            .O(N__52520),
            .I(N__52490));
    InMux I__12626 (
            .O(N__52517),
            .I(N__52487));
    LocalMux I__12625 (
            .O(N__52514),
            .I(N__52484));
    InMux I__12624 (
            .O(N__52513),
            .I(N__52481));
    InMux I__12623 (
            .O(N__52512),
            .I(N__52478));
    Span4Mux_v I__12622 (
            .O(N__52503),
            .I(N__52475));
    Span4Mux_v I__12621 (
            .O(N__52500),
            .I(N__52468));
    LocalMux I__12620 (
            .O(N__52495),
            .I(N__52468));
    LocalMux I__12619 (
            .O(N__52490),
            .I(N__52468));
    LocalMux I__12618 (
            .O(N__52487),
            .I(N__52463));
    Span4Mux_h I__12617 (
            .O(N__52484),
            .I(N__52463));
    LocalMux I__12616 (
            .O(N__52481),
            .I(N__52460));
    LocalMux I__12615 (
            .O(N__52478),
            .I(comm_index_2));
    Odrv4 I__12614 (
            .O(N__52475),
            .I(comm_index_2));
    Odrv4 I__12613 (
            .O(N__52468),
            .I(comm_index_2));
    Odrv4 I__12612 (
            .O(N__52463),
            .I(comm_index_2));
    Odrv4 I__12611 (
            .O(N__52460),
            .I(comm_index_2));
    InMux I__12610 (
            .O(N__52449),
            .I(N__52440));
    CascadeMux I__12609 (
            .O(N__52448),
            .I(N__52429));
    InMux I__12608 (
            .O(N__52447),
            .I(N__52426));
    InMux I__12607 (
            .O(N__52446),
            .I(N__52423));
    InMux I__12606 (
            .O(N__52445),
            .I(N__52420));
    InMux I__12605 (
            .O(N__52444),
            .I(N__52415));
    InMux I__12604 (
            .O(N__52443),
            .I(N__52415));
    LocalMux I__12603 (
            .O(N__52440),
            .I(N__52412));
    CascadeMux I__12602 (
            .O(N__52439),
            .I(N__52406));
    InMux I__12601 (
            .O(N__52438),
            .I(N__52401));
    InMux I__12600 (
            .O(N__52437),
            .I(N__52401));
    InMux I__12599 (
            .O(N__52436),
            .I(N__52396));
    InMux I__12598 (
            .O(N__52435),
            .I(N__52396));
    InMux I__12597 (
            .O(N__52434),
            .I(N__52383));
    InMux I__12596 (
            .O(N__52433),
            .I(N__52383));
    InMux I__12595 (
            .O(N__52432),
            .I(N__52383));
    InMux I__12594 (
            .O(N__52429),
            .I(N__52383));
    LocalMux I__12593 (
            .O(N__52426),
            .I(N__52371));
    LocalMux I__12592 (
            .O(N__52423),
            .I(N__52371));
    LocalMux I__12591 (
            .O(N__52420),
            .I(N__52364));
    LocalMux I__12590 (
            .O(N__52415),
            .I(N__52364));
    Span4Mux_v I__12589 (
            .O(N__52412),
            .I(N__52364));
    InMux I__12588 (
            .O(N__52411),
            .I(N__52355));
    InMux I__12587 (
            .O(N__52410),
            .I(N__52355));
    InMux I__12586 (
            .O(N__52409),
            .I(N__52355));
    InMux I__12585 (
            .O(N__52406),
            .I(N__52355));
    LocalMux I__12584 (
            .O(N__52401),
            .I(N__52350));
    LocalMux I__12583 (
            .O(N__52396),
            .I(N__52350));
    InMux I__12582 (
            .O(N__52395),
            .I(N__52345));
    InMux I__12581 (
            .O(N__52394),
            .I(N__52345));
    InMux I__12580 (
            .O(N__52393),
            .I(N__52340));
    InMux I__12579 (
            .O(N__52392),
            .I(N__52340));
    LocalMux I__12578 (
            .O(N__52383),
            .I(N__52337));
    InMux I__12577 (
            .O(N__52382),
            .I(N__52334));
    InMux I__12576 (
            .O(N__52381),
            .I(N__52325));
    InMux I__12575 (
            .O(N__52380),
            .I(N__52325));
    InMux I__12574 (
            .O(N__52379),
            .I(N__52325));
    InMux I__12573 (
            .O(N__52378),
            .I(N__52325));
    InMux I__12572 (
            .O(N__52377),
            .I(N__52320));
    InMux I__12571 (
            .O(N__52376),
            .I(N__52320));
    Span4Mux_v I__12570 (
            .O(N__52371),
            .I(N__52313));
    Span4Mux_v I__12569 (
            .O(N__52364),
            .I(N__52313));
    LocalMux I__12568 (
            .O(N__52355),
            .I(N__52313));
    Span4Mux_v I__12567 (
            .O(N__52350),
            .I(N__52304));
    LocalMux I__12566 (
            .O(N__52345),
            .I(N__52304));
    LocalMux I__12565 (
            .O(N__52340),
            .I(N__52304));
    Span4Mux_h I__12564 (
            .O(N__52337),
            .I(N__52304));
    LocalMux I__12563 (
            .O(N__52334),
            .I(N__52299));
    LocalMux I__12562 (
            .O(N__52325),
            .I(N__52299));
    LocalMux I__12561 (
            .O(N__52320),
            .I(comm_index_1));
    Odrv4 I__12560 (
            .O(N__52313),
            .I(comm_index_1));
    Odrv4 I__12559 (
            .O(N__52304),
            .I(comm_index_1));
    Odrv12 I__12558 (
            .O(N__52299),
            .I(comm_index_1));
    CascadeMux I__12557 (
            .O(N__52290),
            .I(N__52287));
    InMux I__12556 (
            .O(N__52287),
            .I(N__52282));
    CascadeMux I__12555 (
            .O(N__52286),
            .I(N__52279));
    InMux I__12554 (
            .O(N__52285),
            .I(N__52272));
    LocalMux I__12553 (
            .O(N__52282),
            .I(N__52269));
    InMux I__12552 (
            .O(N__52279),
            .I(N__52266));
    InMux I__12551 (
            .O(N__52278),
            .I(N__52263));
    InMux I__12550 (
            .O(N__52277),
            .I(N__52260));
    CascadeMux I__12549 (
            .O(N__52276),
            .I(N__52257));
    CascadeMux I__12548 (
            .O(N__52275),
            .I(N__52254));
    LocalMux I__12547 (
            .O(N__52272),
            .I(N__52251));
    Span4Mux_h I__12546 (
            .O(N__52269),
            .I(N__52246));
    LocalMux I__12545 (
            .O(N__52266),
            .I(N__52246));
    LocalMux I__12544 (
            .O(N__52263),
            .I(N__52243));
    LocalMux I__12543 (
            .O(N__52260),
            .I(N__52240));
    InMux I__12542 (
            .O(N__52257),
            .I(N__52237));
    InMux I__12541 (
            .O(N__52254),
            .I(N__52234));
    Span12Mux_v I__12540 (
            .O(N__52251),
            .I(N__52231));
    Span4Mux_h I__12539 (
            .O(N__52246),
            .I(N__52228));
    Span4Mux_h I__12538 (
            .O(N__52243),
            .I(N__52225));
    Span4Mux_v I__12537 (
            .O(N__52240),
            .I(N__52220));
    LocalMux I__12536 (
            .O(N__52237),
            .I(N__52220));
    LocalMux I__12535 (
            .O(N__52234),
            .I(N__52217));
    Span12Mux_h I__12534 (
            .O(N__52231),
            .I(N__52214));
    Span4Mux_v I__12533 (
            .O(N__52228),
            .I(N__52209));
    Span4Mux_h I__12532 (
            .O(N__52225),
            .I(N__52209));
    Odrv4 I__12531 (
            .O(N__52220),
            .I(comm_buf_0_5));
    Odrv12 I__12530 (
            .O(N__52217),
            .I(comm_buf_0_5));
    Odrv12 I__12529 (
            .O(N__52214),
            .I(comm_buf_0_5));
    Odrv4 I__12528 (
            .O(N__52209),
            .I(comm_buf_0_5));
    CascadeMux I__12527 (
            .O(N__52200),
            .I(n22503_cascade_));
    InMux I__12526 (
            .O(N__52197),
            .I(N__52194));
    LocalMux I__12525 (
            .O(N__52194),
            .I(N__52191));
    Span4Mux_h I__12524 (
            .O(N__52191),
            .I(N__52188));
    Span4Mux_v I__12523 (
            .O(N__52188),
            .I(N__52185));
    Odrv4 I__12522 (
            .O(N__52185),
            .I(comm_buf_4_5));
    InMux I__12521 (
            .O(N__52182),
            .I(N__52179));
    LocalMux I__12520 (
            .O(N__52179),
            .I(N__52176));
    Odrv4 I__12519 (
            .O(N__52176),
            .I(n22506));
    InMux I__12518 (
            .O(N__52173),
            .I(\ADC_VDC.genclk.n19902 ));
    CEMux I__12517 (
            .O(N__52170),
            .I(N__52166));
    CEMux I__12516 (
            .O(N__52169),
            .I(N__52163));
    LocalMux I__12515 (
            .O(N__52166),
            .I(N__52160));
    LocalMux I__12514 (
            .O(N__52163),
            .I(N__52157));
    Odrv12 I__12513 (
            .O(N__52160),
            .I(\ADC_VDC.genclk.n11900 ));
    Odrv4 I__12512 (
            .O(N__52157),
            .I(\ADC_VDC.genclk.n11900 ));
    CascadeMux I__12511 (
            .O(N__52152),
            .I(N__52147));
    InMux I__12510 (
            .O(N__52151),
            .I(N__52144));
    InMux I__12509 (
            .O(N__52150),
            .I(N__52141));
    InMux I__12508 (
            .O(N__52147),
            .I(N__52138));
    LocalMux I__12507 (
            .O(N__52144),
            .I(N__52135));
    LocalMux I__12506 (
            .O(N__52141),
            .I(N__52132));
    LocalMux I__12505 (
            .O(N__52138),
            .I(N__52129));
    Odrv4 I__12504 (
            .O(N__52135),
            .I(n14350));
    Odrv4 I__12503 (
            .O(N__52132),
            .I(n14350));
    Odrv4 I__12502 (
            .O(N__52129),
            .I(n14350));
    InMux I__12501 (
            .O(N__52122),
            .I(N__52119));
    LocalMux I__12500 (
            .O(N__52119),
            .I(n21453));
    CascadeMux I__12499 (
            .O(N__52116),
            .I(n21454_cascade_));
    CEMux I__12498 (
            .O(N__52113),
            .I(N__52110));
    LocalMux I__12497 (
            .O(N__52110),
            .I(n14_adj_1638));
    InMux I__12496 (
            .O(N__52107),
            .I(N__52104));
    LocalMux I__12495 (
            .O(N__52104),
            .I(N__52101));
    Span4Mux_h I__12494 (
            .O(N__52101),
            .I(N__52098));
    Odrv4 I__12493 (
            .O(N__52098),
            .I(n21481));
    CEMux I__12492 (
            .O(N__52095),
            .I(N__52091));
    InMux I__12491 (
            .O(N__52094),
            .I(N__52087));
    LocalMux I__12490 (
            .O(N__52091),
            .I(N__52084));
    InMux I__12489 (
            .O(N__52090),
            .I(N__52081));
    LocalMux I__12488 (
            .O(N__52087),
            .I(N__52078));
    Span4Mux_v I__12487 (
            .O(N__52084),
            .I(N__52075));
    LocalMux I__12486 (
            .O(N__52081),
            .I(N__52072));
    Span4Mux_h I__12485 (
            .O(N__52078),
            .I(N__52069));
    Span4Mux_h I__12484 (
            .O(N__52075),
            .I(N__52064));
    Span4Mux_v I__12483 (
            .O(N__52072),
            .I(N__52064));
    Span4Mux_h I__12482 (
            .O(N__52069),
            .I(N__52059));
    Span4Mux_h I__12481 (
            .O(N__52064),
            .I(N__52059));
    Odrv4 I__12480 (
            .O(N__52059),
            .I(n12089));
    InMux I__12479 (
            .O(N__52056),
            .I(N__52052));
    InMux I__12478 (
            .O(N__52055),
            .I(N__52049));
    LocalMux I__12477 (
            .O(N__52052),
            .I(comm_length_2));
    LocalMux I__12476 (
            .O(N__52049),
            .I(comm_length_2));
    InMux I__12475 (
            .O(N__52044),
            .I(N__52041));
    LocalMux I__12474 (
            .O(N__52041),
            .I(n6541));
    InMux I__12473 (
            .O(N__52038),
            .I(N__52035));
    LocalMux I__12472 (
            .O(N__52035),
            .I(n21154));
    InMux I__12471 (
            .O(N__52032),
            .I(\ADC_VDC.genclk.n19893 ));
    InMux I__12470 (
            .O(N__52029),
            .I(\ADC_VDC.genclk.n19894 ));
    InMux I__12469 (
            .O(N__52026),
            .I(bfn_19_8_0_));
    InMux I__12468 (
            .O(N__52023),
            .I(\ADC_VDC.genclk.n19896 ));
    InMux I__12467 (
            .O(N__52020),
            .I(\ADC_VDC.genclk.n19897 ));
    InMux I__12466 (
            .O(N__52017),
            .I(\ADC_VDC.genclk.n19898 ));
    InMux I__12465 (
            .O(N__52014),
            .I(\ADC_VDC.genclk.n19899 ));
    InMux I__12464 (
            .O(N__52011),
            .I(\ADC_VDC.genclk.n19900 ));
    InMux I__12463 (
            .O(N__52008),
            .I(\ADC_VDC.genclk.n19901 ));
    InMux I__12462 (
            .O(N__52005),
            .I(N__52001));
    CascadeMux I__12461 (
            .O(N__52004),
            .I(N__51997));
    LocalMux I__12460 (
            .O(N__52001),
            .I(N__51994));
    CascadeMux I__12459 (
            .O(N__52000),
            .I(N__51990));
    InMux I__12458 (
            .O(N__51997),
            .I(N__51987));
    Span4Mux_v I__12457 (
            .O(N__51994),
            .I(N__51982));
    InMux I__12456 (
            .O(N__51993),
            .I(N__51979));
    InMux I__12455 (
            .O(N__51990),
            .I(N__51976));
    LocalMux I__12454 (
            .O(N__51987),
            .I(N__51971));
    InMux I__12453 (
            .O(N__51986),
            .I(N__51966));
    InMux I__12452 (
            .O(N__51985),
            .I(N__51966));
    Span4Mux_h I__12451 (
            .O(N__51982),
            .I(N__51959));
    LocalMux I__12450 (
            .O(N__51979),
            .I(N__51959));
    LocalMux I__12449 (
            .O(N__51976),
            .I(N__51959));
    InMux I__12448 (
            .O(N__51975),
            .I(N__51954));
    InMux I__12447 (
            .O(N__51974),
            .I(N__51954));
    Span4Mux_v I__12446 (
            .O(N__51971),
            .I(N__51951));
    LocalMux I__12445 (
            .O(N__51966),
            .I(N__51948));
    Span4Mux_h I__12444 (
            .O(N__51959),
            .I(N__51943));
    LocalMux I__12443 (
            .O(N__51954),
            .I(N__51943));
    Span4Mux_h I__12442 (
            .O(N__51951),
            .I(N__51939));
    Span4Mux_h I__12441 (
            .O(N__51948),
            .I(N__51934));
    Span4Mux_h I__12440 (
            .O(N__51943),
            .I(N__51934));
    InMux I__12439 (
            .O(N__51942),
            .I(N__51931));
    Span4Mux_v I__12438 (
            .O(N__51939),
            .I(N__51928));
    Sp12to4 I__12437 (
            .O(N__51934),
            .I(N__51923));
    LocalMux I__12436 (
            .O(N__51931),
            .I(N__51923));
    Sp12to4 I__12435 (
            .O(N__51928),
            .I(N__51918));
    Span12Mux_v I__12434 (
            .O(N__51923),
            .I(N__51918));
    Odrv12 I__12433 (
            .O(N__51918),
            .I(VDC_SDO));
    CascadeMux I__12432 (
            .O(N__51915),
            .I(N__51912));
    InMux I__12431 (
            .O(N__51912),
            .I(N__51905));
    InMux I__12430 (
            .O(N__51911),
            .I(N__51900));
    CascadeMux I__12429 (
            .O(N__51910),
            .I(N__51897));
    CascadeMux I__12428 (
            .O(N__51909),
            .I(N__51889));
    InMux I__12427 (
            .O(N__51908),
            .I(N__51886));
    LocalMux I__12426 (
            .O(N__51905),
            .I(N__51883));
    InMux I__12425 (
            .O(N__51904),
            .I(N__51877));
    InMux I__12424 (
            .O(N__51903),
            .I(N__51874));
    LocalMux I__12423 (
            .O(N__51900),
            .I(N__51871));
    InMux I__12422 (
            .O(N__51897),
            .I(N__51868));
    InMux I__12421 (
            .O(N__51896),
            .I(N__51864));
    InMux I__12420 (
            .O(N__51895),
            .I(N__51861));
    InMux I__12419 (
            .O(N__51894),
            .I(N__51853));
    InMux I__12418 (
            .O(N__51893),
            .I(N__51846));
    InMux I__12417 (
            .O(N__51892),
            .I(N__51846));
    InMux I__12416 (
            .O(N__51889),
            .I(N__51846));
    LocalMux I__12415 (
            .O(N__51886),
            .I(N__51843));
    Span4Mux_h I__12414 (
            .O(N__51883),
            .I(N__51840));
    InMux I__12413 (
            .O(N__51882),
            .I(N__51833));
    InMux I__12412 (
            .O(N__51881),
            .I(N__51833));
    InMux I__12411 (
            .O(N__51880),
            .I(N__51833));
    LocalMux I__12410 (
            .O(N__51877),
            .I(N__51828));
    LocalMux I__12409 (
            .O(N__51874),
            .I(N__51828));
    Span4Mux_v I__12408 (
            .O(N__51871),
            .I(N__51823));
    LocalMux I__12407 (
            .O(N__51868),
            .I(N__51823));
    InMux I__12406 (
            .O(N__51867),
            .I(N__51820));
    LocalMux I__12405 (
            .O(N__51864),
            .I(N__51817));
    LocalMux I__12404 (
            .O(N__51861),
            .I(N__51814));
    InMux I__12403 (
            .O(N__51860),
            .I(N__51811));
    InMux I__12402 (
            .O(N__51859),
            .I(N__51806));
    InMux I__12401 (
            .O(N__51858),
            .I(N__51806));
    InMux I__12400 (
            .O(N__51857),
            .I(N__51803));
    InMux I__12399 (
            .O(N__51856),
            .I(N__51800));
    LocalMux I__12398 (
            .O(N__51853),
            .I(N__51789));
    LocalMux I__12397 (
            .O(N__51846),
            .I(N__51789));
    Span4Mux_v I__12396 (
            .O(N__51843),
            .I(N__51789));
    Span4Mux_v I__12395 (
            .O(N__51840),
            .I(N__51789));
    LocalMux I__12394 (
            .O(N__51833),
            .I(N__51789));
    Span12Mux_h I__12393 (
            .O(N__51828),
            .I(N__51786));
    Span4Mux_h I__12392 (
            .O(N__51823),
            .I(N__51783));
    LocalMux I__12391 (
            .O(N__51820),
            .I(\ADC_VDC.adc_state_0 ));
    Odrv4 I__12390 (
            .O(N__51817),
            .I(\ADC_VDC.adc_state_0 ));
    Odrv12 I__12389 (
            .O(N__51814),
            .I(\ADC_VDC.adc_state_0 ));
    LocalMux I__12388 (
            .O(N__51811),
            .I(\ADC_VDC.adc_state_0 ));
    LocalMux I__12387 (
            .O(N__51806),
            .I(\ADC_VDC.adc_state_0 ));
    LocalMux I__12386 (
            .O(N__51803),
            .I(\ADC_VDC.adc_state_0 ));
    LocalMux I__12385 (
            .O(N__51800),
            .I(\ADC_VDC.adc_state_0 ));
    Odrv4 I__12384 (
            .O(N__51789),
            .I(\ADC_VDC.adc_state_0 ));
    Odrv12 I__12383 (
            .O(N__51786),
            .I(\ADC_VDC.adc_state_0 ));
    Odrv4 I__12382 (
            .O(N__51783),
            .I(\ADC_VDC.adc_state_0 ));
    CascadeMux I__12381 (
            .O(N__51762),
            .I(N__51755));
    CascadeMux I__12380 (
            .O(N__51761),
            .I(N__51750));
    InMux I__12379 (
            .O(N__51760),
            .I(N__51747));
    CascadeMux I__12378 (
            .O(N__51759),
            .I(N__51741));
    CascadeMux I__12377 (
            .O(N__51758),
            .I(N__51738));
    InMux I__12376 (
            .O(N__51755),
            .I(N__51735));
    CascadeMux I__12375 (
            .O(N__51754),
            .I(N__51732));
    InMux I__12374 (
            .O(N__51753),
            .I(N__51729));
    InMux I__12373 (
            .O(N__51750),
            .I(N__51726));
    LocalMux I__12372 (
            .O(N__51747),
            .I(N__51723));
    InMux I__12371 (
            .O(N__51746),
            .I(N__51717));
    InMux I__12370 (
            .O(N__51745),
            .I(N__51714));
    InMux I__12369 (
            .O(N__51744),
            .I(N__51691));
    InMux I__12368 (
            .O(N__51741),
            .I(N__51691));
    InMux I__12367 (
            .O(N__51738),
            .I(N__51687));
    LocalMux I__12366 (
            .O(N__51735),
            .I(N__51684));
    InMux I__12365 (
            .O(N__51732),
            .I(N__51681));
    LocalMux I__12364 (
            .O(N__51729),
            .I(N__51674));
    LocalMux I__12363 (
            .O(N__51726),
            .I(N__51674));
    Span4Mux_v I__12362 (
            .O(N__51723),
            .I(N__51674));
    InMux I__12361 (
            .O(N__51722),
            .I(N__51669));
    InMux I__12360 (
            .O(N__51721),
            .I(N__51669));
    InMux I__12359 (
            .O(N__51720),
            .I(N__51666));
    LocalMux I__12358 (
            .O(N__51717),
            .I(N__51661));
    LocalMux I__12357 (
            .O(N__51714),
            .I(N__51661));
    InMux I__12356 (
            .O(N__51713),
            .I(N__51652));
    InMux I__12355 (
            .O(N__51712),
            .I(N__51652));
    InMux I__12354 (
            .O(N__51711),
            .I(N__51652));
    InMux I__12353 (
            .O(N__51710),
            .I(N__51652));
    CascadeMux I__12352 (
            .O(N__51709),
            .I(N__51649));
    CascadeMux I__12351 (
            .O(N__51708),
            .I(N__51645));
    CascadeMux I__12350 (
            .O(N__51707),
            .I(N__51642));
    InMux I__12349 (
            .O(N__51706),
            .I(N__51625));
    InMux I__12348 (
            .O(N__51705),
            .I(N__51625));
    InMux I__12347 (
            .O(N__51704),
            .I(N__51625));
    InMux I__12346 (
            .O(N__51703),
            .I(N__51625));
    InMux I__12345 (
            .O(N__51702),
            .I(N__51616));
    InMux I__12344 (
            .O(N__51701),
            .I(N__51616));
    InMux I__12343 (
            .O(N__51700),
            .I(N__51616));
    InMux I__12342 (
            .O(N__51699),
            .I(N__51616));
    InMux I__12341 (
            .O(N__51698),
            .I(N__51609));
    InMux I__12340 (
            .O(N__51697),
            .I(N__51609));
    InMux I__12339 (
            .O(N__51696),
            .I(N__51609));
    LocalMux I__12338 (
            .O(N__51691),
            .I(N__51606));
    InMux I__12337 (
            .O(N__51690),
            .I(N__51603));
    LocalMux I__12336 (
            .O(N__51687),
            .I(N__51596));
    Span4Mux_v I__12335 (
            .O(N__51684),
            .I(N__51593));
    LocalMux I__12334 (
            .O(N__51681),
            .I(N__51590));
    Span4Mux_h I__12333 (
            .O(N__51674),
            .I(N__51587));
    LocalMux I__12332 (
            .O(N__51669),
            .I(N__51578));
    LocalMux I__12331 (
            .O(N__51666),
            .I(N__51578));
    Span4Mux_v I__12330 (
            .O(N__51661),
            .I(N__51578));
    LocalMux I__12329 (
            .O(N__51652),
            .I(N__51578));
    InMux I__12328 (
            .O(N__51649),
            .I(N__51575));
    InMux I__12327 (
            .O(N__51648),
            .I(N__51560));
    InMux I__12326 (
            .O(N__51645),
            .I(N__51560));
    InMux I__12325 (
            .O(N__51642),
            .I(N__51560));
    InMux I__12324 (
            .O(N__51641),
            .I(N__51560));
    InMux I__12323 (
            .O(N__51640),
            .I(N__51560));
    InMux I__12322 (
            .O(N__51639),
            .I(N__51560));
    InMux I__12321 (
            .O(N__51638),
            .I(N__51560));
    InMux I__12320 (
            .O(N__51637),
            .I(N__51557));
    InMux I__12319 (
            .O(N__51636),
            .I(N__51550));
    InMux I__12318 (
            .O(N__51635),
            .I(N__51550));
    InMux I__12317 (
            .O(N__51634),
            .I(N__51550));
    LocalMux I__12316 (
            .O(N__51625),
            .I(N__51539));
    LocalMux I__12315 (
            .O(N__51616),
            .I(N__51539));
    LocalMux I__12314 (
            .O(N__51609),
            .I(N__51539));
    Span4Mux_v I__12313 (
            .O(N__51606),
            .I(N__51539));
    LocalMux I__12312 (
            .O(N__51603),
            .I(N__51539));
    InMux I__12311 (
            .O(N__51602),
            .I(N__51530));
    InMux I__12310 (
            .O(N__51601),
            .I(N__51530));
    InMux I__12309 (
            .O(N__51600),
            .I(N__51530));
    InMux I__12308 (
            .O(N__51599),
            .I(N__51530));
    Span4Mux_v I__12307 (
            .O(N__51596),
            .I(N__51521));
    Span4Mux_h I__12306 (
            .O(N__51593),
            .I(N__51521));
    Span4Mux_v I__12305 (
            .O(N__51590),
            .I(N__51521));
    Span4Mux_h I__12304 (
            .O(N__51587),
            .I(N__51521));
    Span4Mux_h I__12303 (
            .O(N__51578),
            .I(N__51518));
    LocalMux I__12302 (
            .O(N__51575),
            .I(adc_state_3));
    LocalMux I__12301 (
            .O(N__51560),
            .I(adc_state_3));
    LocalMux I__12300 (
            .O(N__51557),
            .I(adc_state_3));
    LocalMux I__12299 (
            .O(N__51550),
            .I(adc_state_3));
    Odrv4 I__12298 (
            .O(N__51539),
            .I(adc_state_3));
    LocalMux I__12297 (
            .O(N__51530),
            .I(adc_state_3));
    Odrv4 I__12296 (
            .O(N__51521),
            .I(adc_state_3));
    Odrv4 I__12295 (
            .O(N__51518),
            .I(adc_state_3));
    CascadeMux I__12294 (
            .O(N__51501),
            .I(N__51485));
    InMux I__12293 (
            .O(N__51500),
            .I(N__51470));
    InMux I__12292 (
            .O(N__51499),
            .I(N__51457));
    InMux I__12291 (
            .O(N__51498),
            .I(N__51457));
    InMux I__12290 (
            .O(N__51497),
            .I(N__51457));
    InMux I__12289 (
            .O(N__51496),
            .I(N__51457));
    InMux I__12288 (
            .O(N__51495),
            .I(N__51457));
    InMux I__12287 (
            .O(N__51494),
            .I(N__51457));
    InMux I__12286 (
            .O(N__51493),
            .I(N__51452));
    InMux I__12285 (
            .O(N__51492),
            .I(N__51449));
    CascadeMux I__12284 (
            .O(N__51491),
            .I(N__51446));
    CascadeMux I__12283 (
            .O(N__51490),
            .I(N__51443));
    InMux I__12282 (
            .O(N__51489),
            .I(N__51437));
    InMux I__12281 (
            .O(N__51488),
            .I(N__51437));
    InMux I__12280 (
            .O(N__51485),
            .I(N__51424));
    InMux I__12279 (
            .O(N__51484),
            .I(N__51424));
    InMux I__12278 (
            .O(N__51483),
            .I(N__51424));
    InMux I__12277 (
            .O(N__51482),
            .I(N__51424));
    InMux I__12276 (
            .O(N__51481),
            .I(N__51424));
    InMux I__12275 (
            .O(N__51480),
            .I(N__51424));
    InMux I__12274 (
            .O(N__51479),
            .I(N__51421));
    InMux I__12273 (
            .O(N__51478),
            .I(N__51416));
    InMux I__12272 (
            .O(N__51477),
            .I(N__51416));
    InMux I__12271 (
            .O(N__51476),
            .I(N__51409));
    InMux I__12270 (
            .O(N__51475),
            .I(N__51402));
    InMux I__12269 (
            .O(N__51474),
            .I(N__51402));
    InMux I__12268 (
            .O(N__51473),
            .I(N__51402));
    LocalMux I__12267 (
            .O(N__51470),
            .I(N__51399));
    LocalMux I__12266 (
            .O(N__51457),
            .I(N__51396));
    InMux I__12265 (
            .O(N__51456),
            .I(N__51391));
    InMux I__12264 (
            .O(N__51455),
            .I(N__51391));
    LocalMux I__12263 (
            .O(N__51452),
            .I(N__51386));
    LocalMux I__12262 (
            .O(N__51449),
            .I(N__51386));
    InMux I__12261 (
            .O(N__51446),
            .I(N__51380));
    InMux I__12260 (
            .O(N__51443),
            .I(N__51380));
    InMux I__12259 (
            .O(N__51442),
            .I(N__51377));
    LocalMux I__12258 (
            .O(N__51437),
            .I(N__51374));
    LocalMux I__12257 (
            .O(N__51424),
            .I(N__51371));
    LocalMux I__12256 (
            .O(N__51421),
            .I(N__51368));
    LocalMux I__12255 (
            .O(N__51416),
            .I(N__51365));
    CascadeMux I__12254 (
            .O(N__51415),
            .I(N__51358));
    CascadeMux I__12253 (
            .O(N__51414),
            .I(N__51352));
    InMux I__12252 (
            .O(N__51413),
            .I(N__51349));
    InMux I__12251 (
            .O(N__51412),
            .I(N__51346));
    LocalMux I__12250 (
            .O(N__51409),
            .I(N__51339));
    LocalMux I__12249 (
            .O(N__51402),
            .I(N__51339));
    Span4Mux_h I__12248 (
            .O(N__51399),
            .I(N__51332));
    Span4Mux_h I__12247 (
            .O(N__51396),
            .I(N__51332));
    LocalMux I__12246 (
            .O(N__51391),
            .I(N__51332));
    Span4Mux_h I__12245 (
            .O(N__51386),
            .I(N__51324));
    InMux I__12244 (
            .O(N__51385),
            .I(N__51321));
    LocalMux I__12243 (
            .O(N__51380),
            .I(N__51312));
    LocalMux I__12242 (
            .O(N__51377),
            .I(N__51312));
    Span4Mux_h I__12241 (
            .O(N__51374),
            .I(N__51312));
    Span4Mux_v I__12240 (
            .O(N__51371),
            .I(N__51312));
    Span4Mux_v I__12239 (
            .O(N__51368),
            .I(N__51309));
    Span4Mux_h I__12238 (
            .O(N__51365),
            .I(N__51306));
    InMux I__12237 (
            .O(N__51364),
            .I(N__51295));
    InMux I__12236 (
            .O(N__51363),
            .I(N__51295));
    InMux I__12235 (
            .O(N__51362),
            .I(N__51295));
    InMux I__12234 (
            .O(N__51361),
            .I(N__51295));
    InMux I__12233 (
            .O(N__51358),
            .I(N__51295));
    InMux I__12232 (
            .O(N__51357),
            .I(N__51286));
    InMux I__12231 (
            .O(N__51356),
            .I(N__51286));
    InMux I__12230 (
            .O(N__51355),
            .I(N__51286));
    InMux I__12229 (
            .O(N__51352),
            .I(N__51286));
    LocalMux I__12228 (
            .O(N__51349),
            .I(N__51281));
    LocalMux I__12227 (
            .O(N__51346),
            .I(N__51281));
    InMux I__12226 (
            .O(N__51345),
            .I(N__51278));
    InMux I__12225 (
            .O(N__51344),
            .I(N__51275));
    Span4Mux_v I__12224 (
            .O(N__51339),
            .I(N__51272));
    Span4Mux_v I__12223 (
            .O(N__51332),
            .I(N__51269));
    InMux I__12222 (
            .O(N__51331),
            .I(N__51264));
    InMux I__12221 (
            .O(N__51330),
            .I(N__51264));
    InMux I__12220 (
            .O(N__51329),
            .I(N__51257));
    InMux I__12219 (
            .O(N__51328),
            .I(N__51257));
    InMux I__12218 (
            .O(N__51327),
            .I(N__51257));
    Span4Mux_h I__12217 (
            .O(N__51324),
            .I(N__51254));
    LocalMux I__12216 (
            .O(N__51321),
            .I(N__51251));
    Span4Mux_v I__12215 (
            .O(N__51312),
            .I(N__51246));
    Span4Mux_h I__12214 (
            .O(N__51309),
            .I(N__51246));
    Span4Mux_v I__12213 (
            .O(N__51306),
            .I(N__51237));
    LocalMux I__12212 (
            .O(N__51295),
            .I(N__51237));
    LocalMux I__12211 (
            .O(N__51286),
            .I(N__51237));
    Span4Mux_h I__12210 (
            .O(N__51281),
            .I(N__51237));
    LocalMux I__12209 (
            .O(N__51278),
            .I(adc_state_2_adj_1500));
    LocalMux I__12208 (
            .O(N__51275),
            .I(adc_state_2_adj_1500));
    Odrv4 I__12207 (
            .O(N__51272),
            .I(adc_state_2_adj_1500));
    Odrv4 I__12206 (
            .O(N__51269),
            .I(adc_state_2_adj_1500));
    LocalMux I__12205 (
            .O(N__51264),
            .I(adc_state_2_adj_1500));
    LocalMux I__12204 (
            .O(N__51257),
            .I(adc_state_2_adj_1500));
    Odrv4 I__12203 (
            .O(N__51254),
            .I(adc_state_2_adj_1500));
    Odrv4 I__12202 (
            .O(N__51251),
            .I(adc_state_2_adj_1500));
    Odrv4 I__12201 (
            .O(N__51246),
            .I(adc_state_2_adj_1500));
    Odrv4 I__12200 (
            .O(N__51237),
            .I(adc_state_2_adj_1500));
    CascadeMux I__12199 (
            .O(N__51216),
            .I(\ADC_VDC.n52_cascade_ ));
    InMux I__12198 (
            .O(N__51213),
            .I(N__51205));
    InMux I__12197 (
            .O(N__51212),
            .I(N__51198));
    InMux I__12196 (
            .O(N__51211),
            .I(N__51198));
    InMux I__12195 (
            .O(N__51210),
            .I(N__51194));
    InMux I__12194 (
            .O(N__51209),
            .I(N__51191));
    InMux I__12193 (
            .O(N__51208),
            .I(N__51188));
    LocalMux I__12192 (
            .O(N__51205),
            .I(N__51185));
    InMux I__12191 (
            .O(N__51204),
            .I(N__51181));
    InMux I__12190 (
            .O(N__51203),
            .I(N__51176));
    LocalMux I__12189 (
            .O(N__51198),
            .I(N__51171));
    InMux I__12188 (
            .O(N__51197),
            .I(N__51168));
    LocalMux I__12187 (
            .O(N__51194),
            .I(N__51163));
    LocalMux I__12186 (
            .O(N__51191),
            .I(N__51163));
    LocalMux I__12185 (
            .O(N__51188),
            .I(N__51158));
    Span4Mux_h I__12184 (
            .O(N__51185),
            .I(N__51158));
    InMux I__12183 (
            .O(N__51184),
            .I(N__51155));
    LocalMux I__12182 (
            .O(N__51181),
            .I(N__51146));
    InMux I__12181 (
            .O(N__51180),
            .I(N__51142));
    InMux I__12180 (
            .O(N__51179),
            .I(N__51139));
    LocalMux I__12179 (
            .O(N__51176),
            .I(N__51136));
    InMux I__12178 (
            .O(N__51175),
            .I(N__51133));
    InMux I__12177 (
            .O(N__51174),
            .I(N__51130));
    Sp12to4 I__12176 (
            .O(N__51171),
            .I(N__51125));
    LocalMux I__12175 (
            .O(N__51168),
            .I(N__51125));
    Span4Mux_v I__12174 (
            .O(N__51163),
            .I(N__51118));
    Span4Mux_h I__12173 (
            .O(N__51158),
            .I(N__51118));
    LocalMux I__12172 (
            .O(N__51155),
            .I(N__51118));
    InMux I__12171 (
            .O(N__51154),
            .I(N__51111));
    InMux I__12170 (
            .O(N__51153),
            .I(N__51111));
    InMux I__12169 (
            .O(N__51152),
            .I(N__51111));
    InMux I__12168 (
            .O(N__51151),
            .I(N__51104));
    InMux I__12167 (
            .O(N__51150),
            .I(N__51104));
    InMux I__12166 (
            .O(N__51149),
            .I(N__51104));
    Span12Mux_h I__12165 (
            .O(N__51146),
            .I(N__51101));
    InMux I__12164 (
            .O(N__51145),
            .I(N__51098));
    LocalMux I__12163 (
            .O(N__51142),
            .I(\ADC_VDC.adc_state_1 ));
    LocalMux I__12162 (
            .O(N__51139),
            .I(\ADC_VDC.adc_state_1 ));
    Odrv4 I__12161 (
            .O(N__51136),
            .I(\ADC_VDC.adc_state_1 ));
    LocalMux I__12160 (
            .O(N__51133),
            .I(\ADC_VDC.adc_state_1 ));
    LocalMux I__12159 (
            .O(N__51130),
            .I(\ADC_VDC.adc_state_1 ));
    Odrv12 I__12158 (
            .O(N__51125),
            .I(\ADC_VDC.adc_state_1 ));
    Odrv4 I__12157 (
            .O(N__51118),
            .I(\ADC_VDC.adc_state_1 ));
    LocalMux I__12156 (
            .O(N__51111),
            .I(\ADC_VDC.adc_state_1 ));
    LocalMux I__12155 (
            .O(N__51104),
            .I(\ADC_VDC.adc_state_1 ));
    Odrv12 I__12154 (
            .O(N__51101),
            .I(\ADC_VDC.adc_state_1 ));
    LocalMux I__12153 (
            .O(N__51098),
            .I(\ADC_VDC.adc_state_1 ));
    CEMux I__12152 (
            .O(N__51075),
            .I(N__51072));
    LocalMux I__12151 (
            .O(N__51072),
            .I(N__51069));
    Span4Mux_h I__12150 (
            .O(N__51069),
            .I(N__51066));
    Odrv4 I__12149 (
            .O(N__51066),
            .I(\ADC_VDC.n11905 ));
    InMux I__12148 (
            .O(N__51063),
            .I(bfn_19_7_0_));
    InMux I__12147 (
            .O(N__51060),
            .I(\ADC_VDC.genclk.n19888 ));
    InMux I__12146 (
            .O(N__51057),
            .I(\ADC_VDC.genclk.n19889 ));
    InMux I__12145 (
            .O(N__51054),
            .I(\ADC_VDC.genclk.n19890 ));
    InMux I__12144 (
            .O(N__51051),
            .I(\ADC_VDC.genclk.n19891 ));
    InMux I__12143 (
            .O(N__51048),
            .I(\ADC_VDC.genclk.n19892 ));
    InMux I__12142 (
            .O(N__51045),
            .I(N__51041));
    InMux I__12141 (
            .O(N__51044),
            .I(N__51038));
    LocalMux I__12140 (
            .O(N__51041),
            .I(dds0_mclkcnt_5));
    LocalMux I__12139 (
            .O(N__51038),
            .I(dds0_mclkcnt_5));
    InMux I__12138 (
            .O(N__51033),
            .I(n19929));
    InMux I__12137 (
            .O(N__51030),
            .I(N__51027));
    LocalMux I__12136 (
            .O(N__51027),
            .I(n10_adj_1528));
    CascadeMux I__12135 (
            .O(N__51024),
            .I(N__51021));
    InMux I__12134 (
            .O(N__51021),
            .I(N__51015));
    InMux I__12133 (
            .O(N__51020),
            .I(N__51015));
    LocalMux I__12132 (
            .O(N__51015),
            .I(dds0_mclkcnt_6));
    InMux I__12131 (
            .O(N__51012),
            .I(n19930));
    InMux I__12130 (
            .O(N__51009),
            .I(n19931));
    InMux I__12129 (
            .O(N__51006),
            .I(N__51002));
    InMux I__12128 (
            .O(N__51005),
            .I(N__50999));
    LocalMux I__12127 (
            .O(N__51002),
            .I(dds0_mclkcnt_7));
    LocalMux I__12126 (
            .O(N__50999),
            .I(dds0_mclkcnt_7));
    InMux I__12125 (
            .O(N__50994),
            .I(N__50991));
    LocalMux I__12124 (
            .O(N__50991),
            .I(N__50987));
    CascadeMux I__12123 (
            .O(N__50990),
            .I(N__50984));
    Span4Mux_v I__12122 (
            .O(N__50987),
            .I(N__50977));
    InMux I__12121 (
            .O(N__50984),
            .I(N__50972));
    InMux I__12120 (
            .O(N__50983),
            .I(N__50972));
    InMux I__12119 (
            .O(N__50982),
            .I(N__50969));
    InMux I__12118 (
            .O(N__50981),
            .I(N__50966));
    CascadeMux I__12117 (
            .O(N__50980),
            .I(N__50963));
    Span4Mux_h I__12116 (
            .O(N__50977),
            .I(N__50960));
    LocalMux I__12115 (
            .O(N__50972),
            .I(N__50957));
    LocalMux I__12114 (
            .O(N__50969),
            .I(N__50954));
    LocalMux I__12113 (
            .O(N__50966),
            .I(N__50949));
    InMux I__12112 (
            .O(N__50963),
            .I(N__50946));
    Span4Mux_h I__12111 (
            .O(N__50960),
            .I(N__50941));
    Span4Mux_v I__12110 (
            .O(N__50957),
            .I(N__50941));
    Span4Mux_v I__12109 (
            .O(N__50954),
            .I(N__50938));
    InMux I__12108 (
            .O(N__50953),
            .I(N__50933));
    InMux I__12107 (
            .O(N__50952),
            .I(N__50933));
    Span4Mux_h I__12106 (
            .O(N__50949),
            .I(N__50928));
    LocalMux I__12105 (
            .O(N__50946),
            .I(N__50928));
    Span4Mux_h I__12104 (
            .O(N__50941),
            .I(N__50925));
    Span4Mux_h I__12103 (
            .O(N__50938),
            .I(N__50922));
    LocalMux I__12102 (
            .O(N__50933),
            .I(N__50919));
    Sp12to4 I__12101 (
            .O(N__50928),
            .I(N__50916));
    Span4Mux_v I__12100 (
            .O(N__50925),
            .I(N__50913));
    Span4Mux_h I__12099 (
            .O(N__50922),
            .I(N__50908));
    Span4Mux_v I__12098 (
            .O(N__50919),
            .I(N__50908));
    Span12Mux_v I__12097 (
            .O(N__50916),
            .I(N__50905));
    Span4Mux_h I__12096 (
            .O(N__50913),
            .I(N__50902));
    Span4Mux_h I__12095 (
            .O(N__50908),
            .I(N__50899));
    Odrv12 I__12094 (
            .O(N__50905),
            .I(n14716));
    Odrv4 I__12093 (
            .O(N__50902),
            .I(n14716));
    Odrv4 I__12092 (
            .O(N__50899),
            .I(n14716));
    InMux I__12091 (
            .O(N__50892),
            .I(N__50888));
    InMux I__12090 (
            .O(N__50891),
            .I(N__50885));
    LocalMux I__12089 (
            .O(N__50888),
            .I(N__50879));
    LocalMux I__12088 (
            .O(N__50885),
            .I(N__50879));
    InMux I__12087 (
            .O(N__50884),
            .I(N__50876));
    Span4Mux_v I__12086 (
            .O(N__50879),
            .I(N__50870));
    LocalMux I__12085 (
            .O(N__50876),
            .I(N__50870));
    InMux I__12084 (
            .O(N__50875),
            .I(N__50866));
    Span4Mux_v I__12083 (
            .O(N__50870),
            .I(N__50863));
    InMux I__12082 (
            .O(N__50869),
            .I(N__50860));
    LocalMux I__12081 (
            .O(N__50866),
            .I(N__50857));
    Span4Mux_h I__12080 (
            .O(N__50863),
            .I(N__50852));
    LocalMux I__12079 (
            .O(N__50860),
            .I(N__50852));
    Span4Mux_h I__12078 (
            .O(N__50857),
            .I(N__50849));
    Sp12to4 I__12077 (
            .O(N__50852),
            .I(N__50846));
    Sp12to4 I__12076 (
            .O(N__50849),
            .I(N__50843));
    Span12Mux_v I__12075 (
            .O(N__50846),
            .I(N__50840));
    Span12Mux_v I__12074 (
            .O(N__50843),
            .I(N__50837));
    Odrv12 I__12073 (
            .O(N__50840),
            .I(ICE_SPI_MOSI));
    Odrv12 I__12072 (
            .O(N__50837),
            .I(ICE_SPI_MOSI));
    SRMux I__12071 (
            .O(N__50832),
            .I(N__50829));
    LocalMux I__12070 (
            .O(N__50829),
            .I(N__50826));
    Span12Mux_h I__12069 (
            .O(N__50826),
            .I(N__50823));
    Odrv12 I__12068 (
            .O(N__50823),
            .I(\comm_spi.imosi_N_793 ));
    SRMux I__12067 (
            .O(N__50820),
            .I(N__50817));
    LocalMux I__12066 (
            .O(N__50817),
            .I(N__50814));
    Odrv12 I__12065 (
            .O(N__50814),
            .I(\comm_spi.data_tx_7__N_810 ));
    InMux I__12064 (
            .O(N__50811),
            .I(N__50807));
    InMux I__12063 (
            .O(N__50810),
            .I(N__50804));
    LocalMux I__12062 (
            .O(N__50807),
            .I(N__50800));
    LocalMux I__12061 (
            .O(N__50804),
            .I(N__50778));
    ClkMux I__12060 (
            .O(N__50803),
            .I(N__50733));
    Glb2LocalMux I__12059 (
            .O(N__50800),
            .I(N__50733));
    ClkMux I__12058 (
            .O(N__50799),
            .I(N__50733));
    ClkMux I__12057 (
            .O(N__50798),
            .I(N__50733));
    ClkMux I__12056 (
            .O(N__50797),
            .I(N__50733));
    ClkMux I__12055 (
            .O(N__50796),
            .I(N__50733));
    ClkMux I__12054 (
            .O(N__50795),
            .I(N__50733));
    ClkMux I__12053 (
            .O(N__50794),
            .I(N__50733));
    ClkMux I__12052 (
            .O(N__50793),
            .I(N__50733));
    ClkMux I__12051 (
            .O(N__50792),
            .I(N__50733));
    ClkMux I__12050 (
            .O(N__50791),
            .I(N__50733));
    ClkMux I__12049 (
            .O(N__50790),
            .I(N__50733));
    ClkMux I__12048 (
            .O(N__50789),
            .I(N__50733));
    ClkMux I__12047 (
            .O(N__50788),
            .I(N__50733));
    ClkMux I__12046 (
            .O(N__50787),
            .I(N__50733));
    ClkMux I__12045 (
            .O(N__50786),
            .I(N__50733));
    ClkMux I__12044 (
            .O(N__50785),
            .I(N__50733));
    ClkMux I__12043 (
            .O(N__50784),
            .I(N__50733));
    ClkMux I__12042 (
            .O(N__50783),
            .I(N__50733));
    ClkMux I__12041 (
            .O(N__50782),
            .I(N__50733));
    ClkMux I__12040 (
            .O(N__50781),
            .I(N__50733));
    Glb2LocalMux I__12039 (
            .O(N__50778),
            .I(N__50733));
    GlobalMux I__12038 (
            .O(N__50733),
            .I(clk_16MHz));
    InMux I__12037 (
            .O(N__50730),
            .I(N__50724));
    InMux I__12036 (
            .O(N__50729),
            .I(N__50724));
    LocalMux I__12035 (
            .O(N__50724),
            .I(dds0_mclk));
    InMux I__12034 (
            .O(N__50721),
            .I(N__50717));
    InMux I__12033 (
            .O(N__50720),
            .I(N__50714));
    LocalMux I__12032 (
            .O(N__50717),
            .I(N__50711));
    LocalMux I__12031 (
            .O(N__50714),
            .I(N__50707));
    Span4Mux_v I__12030 (
            .O(N__50711),
            .I(N__50704));
    InMux I__12029 (
            .O(N__50710),
            .I(N__50701));
    Span12Mux_v I__12028 (
            .O(N__50707),
            .I(N__50698));
    Odrv4 I__12027 (
            .O(N__50704),
            .I(buf_control_6));
    LocalMux I__12026 (
            .O(N__50701),
            .I(buf_control_6));
    Odrv12 I__12025 (
            .O(N__50698),
            .I(buf_control_6));
    IoInMux I__12024 (
            .O(N__50691),
            .I(N__50688));
    LocalMux I__12023 (
            .O(N__50688),
            .I(N__50685));
    Span4Mux_s3_v I__12022 (
            .O(N__50685),
            .I(N__50682));
    Span4Mux_h I__12021 (
            .O(N__50682),
            .I(N__50679));
    Span4Mux_v I__12020 (
            .O(N__50679),
            .I(N__50676));
    Span4Mux_v I__12019 (
            .O(N__50676),
            .I(N__50673));
    Odrv4 I__12018 (
            .O(N__50673),
            .I(DDS_MCLK));
    InMux I__12017 (
            .O(N__50670),
            .I(N__50667));
    LocalMux I__12016 (
            .O(N__50667),
            .I(N__50664));
    Span4Mux_v I__12015 (
            .O(N__50664),
            .I(N__50660));
    InMux I__12014 (
            .O(N__50663),
            .I(N__50657));
    Span4Mux_h I__12013 (
            .O(N__50660),
            .I(N__50654));
    LocalMux I__12012 (
            .O(N__50657),
            .I(acadc_skipcnt_10));
    Odrv4 I__12011 (
            .O(N__50654),
            .I(acadc_skipcnt_10));
    InMux I__12010 (
            .O(N__50649),
            .I(N__50645));
    InMux I__12009 (
            .O(N__50648),
            .I(N__50641));
    LocalMux I__12008 (
            .O(N__50645),
            .I(N__50638));
    InMux I__12007 (
            .O(N__50644),
            .I(N__50635));
    LocalMux I__12006 (
            .O(N__50641),
            .I(acadc_skipCount_12));
    Odrv4 I__12005 (
            .O(N__50638),
            .I(acadc_skipCount_12));
    LocalMux I__12004 (
            .O(N__50635),
            .I(acadc_skipCount_12));
    CascadeMux I__12003 (
            .O(N__50628),
            .I(N__50625));
    InMux I__12002 (
            .O(N__50625),
            .I(N__50622));
    LocalMux I__12001 (
            .O(N__50622),
            .I(N__50618));
    InMux I__12000 (
            .O(N__50621),
            .I(N__50615));
    Span12Mux_v I__11999 (
            .O(N__50618),
            .I(N__50612));
    LocalMux I__11998 (
            .O(N__50615),
            .I(acadc_skipcnt_12));
    Odrv12 I__11997 (
            .O(N__50612),
            .I(acadc_skipcnt_12));
    InMux I__11996 (
            .O(N__50607),
            .I(N__50600));
    InMux I__11995 (
            .O(N__50606),
            .I(N__50600));
    InMux I__11994 (
            .O(N__50605),
            .I(N__50597));
    LocalMux I__11993 (
            .O(N__50600),
            .I(acadc_skipCount_10));
    LocalMux I__11992 (
            .O(N__50597),
            .I(acadc_skipCount_10));
    InMux I__11991 (
            .O(N__50592),
            .I(N__50589));
    LocalMux I__11990 (
            .O(N__50589),
            .I(N__50586));
    Span4Mux_h I__11989 (
            .O(N__50586),
            .I(N__50583));
    Odrv4 I__11988 (
            .O(N__50583),
            .I(n21));
    CEMux I__11987 (
            .O(N__50580),
            .I(N__50577));
    LocalMux I__11986 (
            .O(N__50577),
            .I(N__50574));
    Span4Mux_v I__11985 (
            .O(N__50574),
            .I(N__50571));
    Odrv4 I__11984 (
            .O(N__50571),
            .I(n11590));
    InMux I__11983 (
            .O(N__50568),
            .I(N__50564));
    InMux I__11982 (
            .O(N__50567),
            .I(N__50561));
    LocalMux I__11981 (
            .O(N__50564),
            .I(dds0_mclkcnt_0));
    LocalMux I__11980 (
            .O(N__50561),
            .I(dds0_mclkcnt_0));
    InMux I__11979 (
            .O(N__50556),
            .I(bfn_18_16_0_));
    CascadeMux I__11978 (
            .O(N__50553),
            .I(N__50549));
    InMux I__11977 (
            .O(N__50552),
            .I(N__50546));
    InMux I__11976 (
            .O(N__50549),
            .I(N__50543));
    LocalMux I__11975 (
            .O(N__50546),
            .I(dds0_mclkcnt_1));
    LocalMux I__11974 (
            .O(N__50543),
            .I(dds0_mclkcnt_1));
    InMux I__11973 (
            .O(N__50538),
            .I(n19925));
    CascadeMux I__11972 (
            .O(N__50535),
            .I(N__50531));
    InMux I__11971 (
            .O(N__50534),
            .I(N__50528));
    InMux I__11970 (
            .O(N__50531),
            .I(N__50525));
    LocalMux I__11969 (
            .O(N__50528),
            .I(dds0_mclkcnt_2));
    LocalMux I__11968 (
            .O(N__50525),
            .I(dds0_mclkcnt_2));
    InMux I__11967 (
            .O(N__50520),
            .I(n19926));
    InMux I__11966 (
            .O(N__50517),
            .I(N__50513));
    InMux I__11965 (
            .O(N__50516),
            .I(N__50510));
    LocalMux I__11964 (
            .O(N__50513),
            .I(dds0_mclkcnt_3));
    LocalMux I__11963 (
            .O(N__50510),
            .I(dds0_mclkcnt_3));
    InMux I__11962 (
            .O(N__50505),
            .I(n19927));
    InMux I__11961 (
            .O(N__50502),
            .I(N__50498));
    InMux I__11960 (
            .O(N__50501),
            .I(N__50495));
    LocalMux I__11959 (
            .O(N__50498),
            .I(dds0_mclkcnt_4));
    LocalMux I__11958 (
            .O(N__50495),
            .I(dds0_mclkcnt_4));
    InMux I__11957 (
            .O(N__50490),
            .I(n19928));
    InMux I__11956 (
            .O(N__50487),
            .I(N__50484));
    LocalMux I__11955 (
            .O(N__50484),
            .I(N__50481));
    Odrv4 I__11954 (
            .O(N__50481),
            .I(n4_adj_1581));
    CascadeMux I__11953 (
            .O(N__50478),
            .I(n21282_cascade_));
    InMux I__11952 (
            .O(N__50475),
            .I(N__50472));
    LocalMux I__11951 (
            .O(N__50472),
            .I(N__50469));
    Odrv4 I__11950 (
            .O(N__50469),
            .I(n22548));
    InMux I__11949 (
            .O(N__50466),
            .I(N__50463));
    LocalMux I__11948 (
            .O(N__50463),
            .I(N__50459));
    InMux I__11947 (
            .O(N__50462),
            .I(N__50456));
    Span4Mux_v I__11946 (
            .O(N__50459),
            .I(N__50450));
    LocalMux I__11945 (
            .O(N__50456),
            .I(N__50450));
    InMux I__11944 (
            .O(N__50455),
            .I(N__50447));
    Span4Mux_v I__11943 (
            .O(N__50450),
            .I(N__50442));
    LocalMux I__11942 (
            .O(N__50447),
            .I(N__50442));
    Span4Mux_v I__11941 (
            .O(N__50442),
            .I(N__50439));
    Span4Mux_h I__11940 (
            .O(N__50439),
            .I(N__50436));
    Odrv4 I__11939 (
            .O(N__50436),
            .I(comm_tx_buf_6));
    InMux I__11938 (
            .O(N__50433),
            .I(N__50430));
    LocalMux I__11937 (
            .O(N__50430),
            .I(N__50427));
    Odrv12 I__11936 (
            .O(N__50427),
            .I(comm_buf_5_5));
    CascadeMux I__11935 (
            .O(N__50424),
            .I(N__50419));
    InMux I__11934 (
            .O(N__50423),
            .I(N__50415));
    InMux I__11933 (
            .O(N__50422),
            .I(N__50411));
    InMux I__11932 (
            .O(N__50419),
            .I(N__50406));
    InMux I__11931 (
            .O(N__50418),
            .I(N__50406));
    LocalMux I__11930 (
            .O(N__50415),
            .I(N__50403));
    InMux I__11929 (
            .O(N__50414),
            .I(N__50400));
    LocalMux I__11928 (
            .O(N__50411),
            .I(N__50397));
    LocalMux I__11927 (
            .O(N__50406),
            .I(N__50394));
    Span4Mux_v I__11926 (
            .O(N__50403),
            .I(N__50391));
    LocalMux I__11925 (
            .O(N__50400),
            .I(N__50388));
    Span4Mux_h I__11924 (
            .O(N__50397),
            .I(N__50385));
    Span4Mux_v I__11923 (
            .O(N__50394),
            .I(N__50382));
    Span4Mux_h I__11922 (
            .O(N__50391),
            .I(N__50375));
    Span4Mux_v I__11921 (
            .O(N__50388),
            .I(N__50375));
    Span4Mux_v I__11920 (
            .O(N__50385),
            .I(N__50375));
    Odrv4 I__11919 (
            .O(N__50382),
            .I(comm_buf_1_5));
    Odrv4 I__11918 (
            .O(N__50375),
            .I(comm_buf_1_5));
    InMux I__11917 (
            .O(N__50370),
            .I(N__50367));
    LocalMux I__11916 (
            .O(N__50367),
            .I(N__50364));
    Odrv4 I__11915 (
            .O(N__50364),
            .I(comm_buf_3_5));
    CascadeMux I__11914 (
            .O(N__50361),
            .I(n17698_cascade_));
    CascadeMux I__11913 (
            .O(N__50358),
            .I(n21270_cascade_));
    CEMux I__11912 (
            .O(N__50355),
            .I(N__50351));
    CEMux I__11911 (
            .O(N__50354),
            .I(N__50348));
    LocalMux I__11910 (
            .O(N__50351),
            .I(N__50343));
    LocalMux I__11909 (
            .O(N__50348),
            .I(N__50343));
    Span4Mux_v I__11908 (
            .O(N__50343),
            .I(N__50338));
    CEMux I__11907 (
            .O(N__50342),
            .I(N__50335));
    CEMux I__11906 (
            .O(N__50341),
            .I(N__50330));
    Span4Mux_h I__11905 (
            .O(N__50338),
            .I(N__50325));
    LocalMux I__11904 (
            .O(N__50335),
            .I(N__50325));
    CEMux I__11903 (
            .O(N__50334),
            .I(N__50322));
    CEMux I__11902 (
            .O(N__50333),
            .I(N__50318));
    LocalMux I__11901 (
            .O(N__50330),
            .I(N__50315));
    Span4Mux_h I__11900 (
            .O(N__50325),
            .I(N__50312));
    LocalMux I__11899 (
            .O(N__50322),
            .I(N__50309));
    InMux I__11898 (
            .O(N__50321),
            .I(N__50306));
    LocalMux I__11897 (
            .O(N__50318),
            .I(N__50302));
    Span4Mux_h I__11896 (
            .O(N__50315),
            .I(N__50299));
    Sp12to4 I__11895 (
            .O(N__50312),
            .I(N__50296));
    Span4Mux_v I__11894 (
            .O(N__50309),
            .I(N__50291));
    LocalMux I__11893 (
            .O(N__50306),
            .I(N__50291));
    CEMux I__11892 (
            .O(N__50305),
            .I(N__50288));
    Span12Mux_h I__11891 (
            .O(N__50302),
            .I(N__50285));
    Span4Mux_v I__11890 (
            .O(N__50299),
            .I(N__50282));
    Span12Mux_v I__11889 (
            .O(N__50296),
            .I(N__50279));
    Span4Mux_h I__11888 (
            .O(N__50291),
            .I(N__50276));
    LocalMux I__11887 (
            .O(N__50288),
            .I(n12541));
    Odrv12 I__11886 (
            .O(N__50285),
            .I(n12541));
    Odrv4 I__11885 (
            .O(N__50282),
            .I(n12541));
    Odrv12 I__11884 (
            .O(N__50279),
            .I(n12541));
    Odrv4 I__11883 (
            .O(N__50276),
            .I(n12541));
    SRMux I__11882 (
            .O(N__50265),
            .I(N__50262));
    LocalMux I__11881 (
            .O(N__50262),
            .I(N__50258));
    SRMux I__11880 (
            .O(N__50261),
            .I(N__50255));
    Span4Mux_h I__11879 (
            .O(N__50258),
            .I(N__50251));
    LocalMux I__11878 (
            .O(N__50255),
            .I(N__50247));
    SRMux I__11877 (
            .O(N__50254),
            .I(N__50244));
    Span4Mux_h I__11876 (
            .O(N__50251),
            .I(N__50240));
    SRMux I__11875 (
            .O(N__50250),
            .I(N__50237));
    Span4Mux_h I__11874 (
            .O(N__50247),
            .I(N__50232));
    LocalMux I__11873 (
            .O(N__50244),
            .I(N__50232));
    SRMux I__11872 (
            .O(N__50243),
            .I(N__50228));
    Span4Mux_v I__11871 (
            .O(N__50240),
            .I(N__50224));
    LocalMux I__11870 (
            .O(N__50237),
            .I(N__50219));
    Span4Mux_v I__11869 (
            .O(N__50232),
            .I(N__50219));
    SRMux I__11868 (
            .O(N__50231),
            .I(N__50216));
    LocalMux I__11867 (
            .O(N__50228),
            .I(N__50213));
    SRMux I__11866 (
            .O(N__50227),
            .I(N__50210));
    Sp12to4 I__11865 (
            .O(N__50224),
            .I(N__50207));
    Span4Mux_v I__11864 (
            .O(N__50219),
            .I(N__50204));
    LocalMux I__11863 (
            .O(N__50216),
            .I(N__50201));
    Span4Mux_h I__11862 (
            .O(N__50213),
            .I(N__50198));
    LocalMux I__11861 (
            .O(N__50210),
            .I(N__50191));
    Span12Mux_s10_h I__11860 (
            .O(N__50207),
            .I(N__50191));
    Sp12to4 I__11859 (
            .O(N__50204),
            .I(N__50191));
    Odrv12 I__11858 (
            .O(N__50201),
            .I(n15007));
    Odrv4 I__11857 (
            .O(N__50198),
            .I(n15007));
    Odrv12 I__11856 (
            .O(N__50191),
            .I(n15007));
    CascadeMux I__11855 (
            .O(N__50184),
            .I(n20996_cascade_));
    InMux I__11854 (
            .O(N__50181),
            .I(N__50178));
    LocalMux I__11853 (
            .O(N__50178),
            .I(n12_adj_1663));
    InMux I__11852 (
            .O(N__50175),
            .I(N__50172));
    LocalMux I__11851 (
            .O(N__50172),
            .I(n20996));
    CascadeMux I__11850 (
            .O(N__50169),
            .I(N__50166));
    InMux I__11849 (
            .O(N__50166),
            .I(N__50162));
    InMux I__11848 (
            .O(N__50165),
            .I(N__50159));
    LocalMux I__11847 (
            .O(N__50162),
            .I(N__50153));
    LocalMux I__11846 (
            .O(N__50159),
            .I(N__50150));
    InMux I__11845 (
            .O(N__50158),
            .I(N__50147));
    InMux I__11844 (
            .O(N__50157),
            .I(N__50142));
    InMux I__11843 (
            .O(N__50156),
            .I(N__50139));
    Span4Mux_v I__11842 (
            .O(N__50153),
            .I(N__50136));
    Span4Mux_h I__11841 (
            .O(N__50150),
            .I(N__50131));
    LocalMux I__11840 (
            .O(N__50147),
            .I(N__50131));
    InMux I__11839 (
            .O(N__50146),
            .I(N__50128));
    InMux I__11838 (
            .O(N__50145),
            .I(N__50125));
    LocalMux I__11837 (
            .O(N__50142),
            .I(N__50122));
    LocalMux I__11836 (
            .O(N__50139),
            .I(N__50119));
    Span4Mux_h I__11835 (
            .O(N__50136),
            .I(N__50114));
    Span4Mux_v I__11834 (
            .O(N__50131),
            .I(N__50114));
    LocalMux I__11833 (
            .O(N__50128),
            .I(N__50109));
    LocalMux I__11832 (
            .O(N__50125),
            .I(N__50109));
    Span4Mux_v I__11831 (
            .O(N__50122),
            .I(N__50105));
    Span4Mux_v I__11830 (
            .O(N__50119),
            .I(N__50098));
    Span4Mux_h I__11829 (
            .O(N__50114),
            .I(N__50098));
    Span4Mux_v I__11828 (
            .O(N__50109),
            .I(N__50098));
    InMux I__11827 (
            .O(N__50108),
            .I(N__50095));
    Span4Mux_h I__11826 (
            .O(N__50105),
            .I(N__50091));
    Sp12to4 I__11825 (
            .O(N__50098),
            .I(N__50088));
    LocalMux I__11824 (
            .O(N__50095),
            .I(N__50085));
    InMux I__11823 (
            .O(N__50094),
            .I(N__50082));
    Odrv4 I__11822 (
            .O(N__50091),
            .I(comm_rx_buf_2));
    Odrv12 I__11821 (
            .O(N__50088),
            .I(comm_rx_buf_2));
    Odrv12 I__11820 (
            .O(N__50085),
            .I(comm_rx_buf_2));
    LocalMux I__11819 (
            .O(N__50082),
            .I(comm_rx_buf_2));
    InMux I__11818 (
            .O(N__50073),
            .I(N__50069));
    InMux I__11817 (
            .O(N__50072),
            .I(N__50066));
    LocalMux I__11816 (
            .O(N__50069),
            .I(comm_buf_6_2));
    LocalMux I__11815 (
            .O(N__50066),
            .I(comm_buf_6_2));
    InMux I__11814 (
            .O(N__50061),
            .I(N__50058));
    LocalMux I__11813 (
            .O(N__50058),
            .I(N__50055));
    Span4Mux_v I__11812 (
            .O(N__50055),
            .I(N__50052));
    Odrv4 I__11811 (
            .O(N__50052),
            .I(comm_buf_5_0));
    InMux I__11810 (
            .O(N__50049),
            .I(N__50046));
    LocalMux I__11809 (
            .O(N__50046),
            .I(N__50043));
    Span4Mux_v I__11808 (
            .O(N__50043),
            .I(N__50040));
    Odrv4 I__11807 (
            .O(N__50040),
            .I(comm_buf_4_0));
    InMux I__11806 (
            .O(N__50037),
            .I(N__50034));
    LocalMux I__11805 (
            .O(N__50034),
            .I(n4_adj_1457));
    InMux I__11804 (
            .O(N__50031),
            .I(N__50028));
    LocalMux I__11803 (
            .O(N__50028),
            .I(N__50025));
    Span4Mux_v I__11802 (
            .O(N__50025),
            .I(N__50022));
    Odrv4 I__11801 (
            .O(N__50022),
            .I(comm_buf_5_1));
    InMux I__11800 (
            .O(N__50019),
            .I(N__50016));
    LocalMux I__11799 (
            .O(N__50016),
            .I(N__50013));
    Span4Mux_v I__11798 (
            .O(N__50013),
            .I(N__50010));
    Odrv4 I__11797 (
            .O(N__50010),
            .I(comm_buf_4_1));
    InMux I__11796 (
            .O(N__50007),
            .I(N__50004));
    LocalMux I__11795 (
            .O(N__50004),
            .I(N__49999));
    InMux I__11794 (
            .O(N__50003),
            .I(N__49994));
    InMux I__11793 (
            .O(N__50002),
            .I(N__49994));
    Span4Mux_v I__11792 (
            .O(N__49999),
            .I(N__49988));
    LocalMux I__11791 (
            .O(N__49994),
            .I(N__49988));
    InMux I__11790 (
            .O(N__49993),
            .I(N__49985));
    Span4Mux_h I__11789 (
            .O(N__49988),
            .I(N__49982));
    LocalMux I__11788 (
            .O(N__49985),
            .I(comm_cmd_7));
    Odrv4 I__11787 (
            .O(N__49982),
            .I(comm_cmd_7));
    InMux I__11786 (
            .O(N__49977),
            .I(N__49974));
    LocalMux I__11785 (
            .O(N__49974),
            .I(N__49970));
    InMux I__11784 (
            .O(N__49973),
            .I(N__49967));
    Span12Mux_h I__11783 (
            .O(N__49970),
            .I(N__49964));
    LocalMux I__11782 (
            .O(N__49967),
            .I(comm_buf_6_1));
    Odrv12 I__11781 (
            .O(N__49964),
            .I(comm_buf_6_1));
    InMux I__11780 (
            .O(N__49959),
            .I(N__49956));
    LocalMux I__11779 (
            .O(N__49956),
            .I(n4_adj_1588));
    CascadeMux I__11778 (
            .O(N__49953),
            .I(n21433_cascade_));
    CascadeMux I__11777 (
            .O(N__49950),
            .I(n22419_cascade_));
    InMux I__11776 (
            .O(N__49947),
            .I(N__49944));
    LocalMux I__11775 (
            .O(N__49944),
            .I(N__49939));
    InMux I__11774 (
            .O(N__49943),
            .I(N__49936));
    InMux I__11773 (
            .O(N__49942),
            .I(N__49933));
    Span4Mux_v I__11772 (
            .O(N__49939),
            .I(N__49928));
    LocalMux I__11771 (
            .O(N__49936),
            .I(N__49923));
    LocalMux I__11770 (
            .O(N__49933),
            .I(N__49923));
    InMux I__11769 (
            .O(N__49932),
            .I(N__49920));
    InMux I__11768 (
            .O(N__49931),
            .I(N__49917));
    Odrv4 I__11767 (
            .O(N__49928),
            .I(n21085));
    Odrv4 I__11766 (
            .O(N__49923),
            .I(n21085));
    LocalMux I__11765 (
            .O(N__49920),
            .I(n21085));
    LocalMux I__11764 (
            .O(N__49917),
            .I(n21085));
    CascadeMux I__11763 (
            .O(N__49908),
            .I(n7_adj_1458_cascade_));
    InMux I__11762 (
            .O(N__49905),
            .I(N__49902));
    LocalMux I__11761 (
            .O(N__49902),
            .I(N__49899));
    Span4Mux_h I__11760 (
            .O(N__49899),
            .I(N__49896));
    Span4Mux_v I__11759 (
            .O(N__49896),
            .I(N__49893));
    Odrv4 I__11758 (
            .O(N__49893),
            .I(buf_data_vac_20));
    InMux I__11757 (
            .O(N__49890),
            .I(N__49887));
    LocalMux I__11756 (
            .O(N__49887),
            .I(N__49884));
    Span4Mux_h I__11755 (
            .O(N__49884),
            .I(N__49881));
    Odrv4 I__11754 (
            .O(N__49881),
            .I(comm_buf_3_4));
    InMux I__11753 (
            .O(N__49878),
            .I(N__49872));
    InMux I__11752 (
            .O(N__49877),
            .I(N__49869));
    InMux I__11751 (
            .O(N__49876),
            .I(N__49864));
    InMux I__11750 (
            .O(N__49875),
            .I(N__49861));
    LocalMux I__11749 (
            .O(N__49872),
            .I(N__49857));
    LocalMux I__11748 (
            .O(N__49869),
            .I(N__49853));
    InMux I__11747 (
            .O(N__49868),
            .I(N__49850));
    InMux I__11746 (
            .O(N__49867),
            .I(N__49847));
    LocalMux I__11745 (
            .O(N__49864),
            .I(N__49844));
    LocalMux I__11744 (
            .O(N__49861),
            .I(N__49841));
    InMux I__11743 (
            .O(N__49860),
            .I(N__49838));
    Span4Mux_v I__11742 (
            .O(N__49857),
            .I(N__49835));
    InMux I__11741 (
            .O(N__49856),
            .I(N__49832));
    Span4Mux_v I__11740 (
            .O(N__49853),
            .I(N__49827));
    LocalMux I__11739 (
            .O(N__49850),
            .I(N__49827));
    LocalMux I__11738 (
            .O(N__49847),
            .I(N__49824));
    Span4Mux_h I__11737 (
            .O(N__49844),
            .I(N__49821));
    Span4Mux_h I__11736 (
            .O(N__49841),
            .I(N__49816));
    LocalMux I__11735 (
            .O(N__49838),
            .I(N__49816));
    Span4Mux_h I__11734 (
            .O(N__49835),
            .I(N__49811));
    LocalMux I__11733 (
            .O(N__49832),
            .I(N__49811));
    Span4Mux_v I__11732 (
            .O(N__49827),
            .I(N__49805));
    Span4Mux_v I__11731 (
            .O(N__49824),
            .I(N__49805));
    Span4Mux_h I__11730 (
            .O(N__49821),
            .I(N__49798));
    Span4Mux_v I__11729 (
            .O(N__49816),
            .I(N__49798));
    Span4Mux_h I__11728 (
            .O(N__49811),
            .I(N__49798));
    InMux I__11727 (
            .O(N__49810),
            .I(N__49795));
    Odrv4 I__11726 (
            .O(N__49805),
            .I(comm_rx_buf_3));
    Odrv4 I__11725 (
            .O(N__49798),
            .I(comm_rx_buf_3));
    LocalMux I__11724 (
            .O(N__49795),
            .I(comm_rx_buf_3));
    InMux I__11723 (
            .O(N__49788),
            .I(N__49785));
    LocalMux I__11722 (
            .O(N__49785),
            .I(N__49782));
    Span4Mux_v I__11721 (
            .O(N__49782),
            .I(N__49779));
    Odrv4 I__11720 (
            .O(N__49779),
            .I(buf_data_vac_19));
    CascadeMux I__11719 (
            .O(N__49776),
            .I(N__49773));
    InMux I__11718 (
            .O(N__49773),
            .I(N__49770));
    LocalMux I__11717 (
            .O(N__49770),
            .I(comm_buf_3_3));
    InMux I__11716 (
            .O(N__49767),
            .I(N__49764));
    LocalMux I__11715 (
            .O(N__49764),
            .I(N__49761));
    Span4Mux_h I__11714 (
            .O(N__49761),
            .I(N__49758));
    Odrv4 I__11713 (
            .O(N__49758),
            .I(buf_data_vac_18));
    CascadeMux I__11712 (
            .O(N__49755),
            .I(N__49752));
    InMux I__11711 (
            .O(N__49752),
            .I(N__49749));
    LocalMux I__11710 (
            .O(N__49749),
            .I(comm_buf_3_2));
    CascadeMux I__11709 (
            .O(N__49746),
            .I(N__49742));
    CascadeMux I__11708 (
            .O(N__49745),
            .I(N__49739));
    InMux I__11707 (
            .O(N__49742),
            .I(N__49736));
    InMux I__11706 (
            .O(N__49739),
            .I(N__49733));
    LocalMux I__11705 (
            .O(N__49736),
            .I(N__49730));
    LocalMux I__11704 (
            .O(N__49733),
            .I(N__49727));
    Span4Mux_h I__11703 (
            .O(N__49730),
            .I(N__49724));
    Span4Mux_v I__11702 (
            .O(N__49727),
            .I(N__49718));
    Span4Mux_h I__11701 (
            .O(N__49724),
            .I(N__49714));
    InMux I__11700 (
            .O(N__49723),
            .I(N__49711));
    InMux I__11699 (
            .O(N__49722),
            .I(N__49708));
    InMux I__11698 (
            .O(N__49721),
            .I(N__49705));
    Span4Mux_h I__11697 (
            .O(N__49718),
            .I(N__49701));
    InMux I__11696 (
            .O(N__49717),
            .I(N__49698));
    Span4Mux_h I__11695 (
            .O(N__49714),
            .I(N__49693));
    LocalMux I__11694 (
            .O(N__49711),
            .I(N__49693));
    LocalMux I__11693 (
            .O(N__49708),
            .I(N__49690));
    LocalMux I__11692 (
            .O(N__49705),
            .I(N__49687));
    InMux I__11691 (
            .O(N__49704),
            .I(N__49684));
    Span4Mux_h I__11690 (
            .O(N__49701),
            .I(N__49679));
    LocalMux I__11689 (
            .O(N__49698),
            .I(N__49679));
    Span4Mux_v I__11688 (
            .O(N__49693),
            .I(N__49675));
    Span4Mux_h I__11687 (
            .O(N__49690),
            .I(N__49672));
    Span4Mux_h I__11686 (
            .O(N__49687),
            .I(N__49669));
    LocalMux I__11685 (
            .O(N__49684),
            .I(N__49666));
    Span4Mux_h I__11684 (
            .O(N__49679),
            .I(N__49663));
    InMux I__11683 (
            .O(N__49678),
            .I(N__49660));
    Sp12to4 I__11682 (
            .O(N__49675),
            .I(N__49656));
    Span4Mux_v I__11681 (
            .O(N__49672),
            .I(N__49649));
    Span4Mux_h I__11680 (
            .O(N__49669),
            .I(N__49649));
    Span4Mux_h I__11679 (
            .O(N__49666),
            .I(N__49649));
    Span4Mux_v I__11678 (
            .O(N__49663),
            .I(N__49644));
    LocalMux I__11677 (
            .O(N__49660),
            .I(N__49644));
    InMux I__11676 (
            .O(N__49659),
            .I(N__49641));
    Odrv12 I__11675 (
            .O(N__49656),
            .I(comm_rx_buf_1));
    Odrv4 I__11674 (
            .O(N__49649),
            .I(comm_rx_buf_1));
    Odrv4 I__11673 (
            .O(N__49644),
            .I(comm_rx_buf_1));
    LocalMux I__11672 (
            .O(N__49641),
            .I(comm_rx_buf_1));
    InMux I__11671 (
            .O(N__49632),
            .I(N__49629));
    LocalMux I__11670 (
            .O(N__49629),
            .I(N__49626));
    Odrv12 I__11669 (
            .O(N__49626),
            .I(buf_data_vac_17));
    InMux I__11668 (
            .O(N__49623),
            .I(N__49620));
    LocalMux I__11667 (
            .O(N__49620),
            .I(N__49617));
    Odrv12 I__11666 (
            .O(N__49617),
            .I(comm_buf_5_6));
    InMux I__11665 (
            .O(N__49614),
            .I(N__49611));
    LocalMux I__11664 (
            .O(N__49611),
            .I(N__49608));
    Span4Mux_v I__11663 (
            .O(N__49608),
            .I(N__49605));
    Odrv4 I__11662 (
            .O(N__49605),
            .I(comm_buf_4_6));
    InMux I__11661 (
            .O(N__49602),
            .I(N__49599));
    LocalMux I__11660 (
            .O(N__49599),
            .I(comm_buf_2_6));
    CascadeMux I__11659 (
            .O(N__49596),
            .I(N__49593));
    InMux I__11658 (
            .O(N__49593),
            .I(N__49590));
    LocalMux I__11657 (
            .O(N__49590),
            .I(comm_buf_3_6));
    CascadeMux I__11656 (
            .O(N__49587),
            .I(N__49582));
    CascadeMux I__11655 (
            .O(N__49586),
            .I(N__49579));
    CascadeMux I__11654 (
            .O(N__49585),
            .I(N__49576));
    InMux I__11653 (
            .O(N__49582),
            .I(N__49573));
    InMux I__11652 (
            .O(N__49579),
            .I(N__49570));
    InMux I__11651 (
            .O(N__49576),
            .I(N__49564));
    LocalMux I__11650 (
            .O(N__49573),
            .I(N__49561));
    LocalMux I__11649 (
            .O(N__49570),
            .I(N__49558));
    CascadeMux I__11648 (
            .O(N__49569),
            .I(N__49554));
    InMux I__11647 (
            .O(N__49568),
            .I(N__49549));
    InMux I__11646 (
            .O(N__49567),
            .I(N__49549));
    LocalMux I__11645 (
            .O(N__49564),
            .I(N__49546));
    Span4Mux_v I__11644 (
            .O(N__49561),
            .I(N__49541));
    Span4Mux_v I__11643 (
            .O(N__49558),
            .I(N__49541));
    InMux I__11642 (
            .O(N__49557),
            .I(N__49538));
    InMux I__11641 (
            .O(N__49554),
            .I(N__49534));
    LocalMux I__11640 (
            .O(N__49549),
            .I(N__49531));
    Span4Mux_v I__11639 (
            .O(N__49546),
            .I(N__49524));
    Span4Mux_h I__11638 (
            .O(N__49541),
            .I(N__49524));
    LocalMux I__11637 (
            .O(N__49538),
            .I(N__49524));
    InMux I__11636 (
            .O(N__49537),
            .I(N__49521));
    LocalMux I__11635 (
            .O(N__49534),
            .I(N__49518));
    Span4Mux_h I__11634 (
            .O(N__49531),
            .I(N__49515));
    Span4Mux_h I__11633 (
            .O(N__49524),
            .I(N__49512));
    LocalMux I__11632 (
            .O(N__49521),
            .I(N__49505));
    Span4Mux_h I__11631 (
            .O(N__49518),
            .I(N__49505));
    Span4Mux_h I__11630 (
            .O(N__49515),
            .I(N__49505));
    Odrv4 I__11629 (
            .O(N__49512),
            .I(comm_buf_0_6));
    Odrv4 I__11628 (
            .O(N__49505),
            .I(comm_buf_0_6));
    CascadeMux I__11627 (
            .O(N__49500),
            .I(n22545_cascade_));
    CascadeMux I__11626 (
            .O(N__49497),
            .I(N__49491));
    InMux I__11625 (
            .O(N__49496),
            .I(N__49488));
    CascadeMux I__11624 (
            .O(N__49495),
            .I(N__49483));
    InMux I__11623 (
            .O(N__49494),
            .I(N__49480));
    InMux I__11622 (
            .O(N__49491),
            .I(N__49477));
    LocalMux I__11621 (
            .O(N__49488),
            .I(N__49474));
    CascadeMux I__11620 (
            .O(N__49487),
            .I(N__49471));
    InMux I__11619 (
            .O(N__49486),
            .I(N__49468));
    InMux I__11618 (
            .O(N__49483),
            .I(N__49465));
    LocalMux I__11617 (
            .O(N__49480),
            .I(N__49462));
    LocalMux I__11616 (
            .O(N__49477),
            .I(N__49459));
    Span4Mux_v I__11615 (
            .O(N__49474),
            .I(N__49456));
    InMux I__11614 (
            .O(N__49471),
            .I(N__49453));
    LocalMux I__11613 (
            .O(N__49468),
            .I(N__49450));
    LocalMux I__11612 (
            .O(N__49465),
            .I(N__49445));
    Span4Mux_h I__11611 (
            .O(N__49462),
            .I(N__49445));
    Span4Mux_h I__11610 (
            .O(N__49459),
            .I(N__49440));
    Span4Mux_h I__11609 (
            .O(N__49456),
            .I(N__49440));
    LocalMux I__11608 (
            .O(N__49453),
            .I(N__49433));
    Span4Mux_h I__11607 (
            .O(N__49450),
            .I(N__49433));
    Span4Mux_h I__11606 (
            .O(N__49445),
            .I(N__49433));
    Odrv4 I__11605 (
            .O(N__49440),
            .I(comm_buf_1_6));
    Odrv4 I__11604 (
            .O(N__49433),
            .I(comm_buf_1_6));
    CEMux I__11603 (
            .O(N__49428),
            .I(N__49425));
    LocalMux I__11602 (
            .O(N__49425),
            .I(N__49421));
    InMux I__11601 (
            .O(N__49424),
            .I(N__49418));
    Odrv4 I__11600 (
            .O(N__49421),
            .I(n12353));
    LocalMux I__11599 (
            .O(N__49418),
            .I(n12353));
    SRMux I__11598 (
            .O(N__49413),
            .I(N__49410));
    LocalMux I__11597 (
            .O(N__49410),
            .I(N__49407));
    Span4Mux_h I__11596 (
            .O(N__49407),
            .I(N__49404));
    Odrv4 I__11595 (
            .O(N__49404),
            .I(n14979));
    InMux I__11594 (
            .O(N__49401),
            .I(N__49398));
    LocalMux I__11593 (
            .O(N__49398),
            .I(N__49395));
    Odrv12 I__11592 (
            .O(N__49395),
            .I(n21588));
    CascadeMux I__11591 (
            .O(N__49392),
            .I(N__49379));
    CascadeMux I__11590 (
            .O(N__49391),
            .I(N__49371));
    CascadeMux I__11589 (
            .O(N__49390),
            .I(N__49366));
    CascadeMux I__11588 (
            .O(N__49389),
            .I(N__49362));
    InMux I__11587 (
            .O(N__49388),
            .I(N__49356));
    InMux I__11586 (
            .O(N__49387),
            .I(N__49356));
    CascadeMux I__11585 (
            .O(N__49386),
            .I(N__49352));
    InMux I__11584 (
            .O(N__49385),
            .I(N__49347));
    InMux I__11583 (
            .O(N__49384),
            .I(N__49342));
    InMux I__11582 (
            .O(N__49383),
            .I(N__49342));
    CascadeMux I__11581 (
            .O(N__49382),
            .I(N__49338));
    InMux I__11580 (
            .O(N__49379),
            .I(N__49332));
    InMux I__11579 (
            .O(N__49378),
            .I(N__49326));
    InMux I__11578 (
            .O(N__49377),
            .I(N__49326));
    CascadeMux I__11577 (
            .O(N__49376),
            .I(N__49319));
    CascadeMux I__11576 (
            .O(N__49375),
            .I(N__49313));
    InMux I__11575 (
            .O(N__49374),
            .I(N__49306));
    InMux I__11574 (
            .O(N__49371),
            .I(N__49298));
    CascadeMux I__11573 (
            .O(N__49370),
            .I(N__49294));
    InMux I__11572 (
            .O(N__49369),
            .I(N__49291));
    InMux I__11571 (
            .O(N__49366),
            .I(N__49284));
    InMux I__11570 (
            .O(N__49365),
            .I(N__49284));
    InMux I__11569 (
            .O(N__49362),
            .I(N__49284));
    CascadeMux I__11568 (
            .O(N__49361),
            .I(N__49281));
    LocalMux I__11567 (
            .O(N__49356),
            .I(N__49276));
    CascadeMux I__11566 (
            .O(N__49355),
            .I(N__49273));
    InMux I__11565 (
            .O(N__49352),
            .I(N__49269));
    InMux I__11564 (
            .O(N__49351),
            .I(N__49264));
    InMux I__11563 (
            .O(N__49350),
            .I(N__49264));
    LocalMux I__11562 (
            .O(N__49347),
            .I(N__49259));
    LocalMux I__11561 (
            .O(N__49342),
            .I(N__49259));
    CascadeMux I__11560 (
            .O(N__49341),
            .I(N__49255));
    InMux I__11559 (
            .O(N__49338),
            .I(N__49252));
    InMux I__11558 (
            .O(N__49337),
            .I(N__49249));
    InMux I__11557 (
            .O(N__49336),
            .I(N__49244));
    InMux I__11556 (
            .O(N__49335),
            .I(N__49244));
    LocalMux I__11555 (
            .O(N__49332),
            .I(N__49239));
    CascadeMux I__11554 (
            .O(N__49331),
            .I(N__49236));
    LocalMux I__11553 (
            .O(N__49326),
            .I(N__49231));
    InMux I__11552 (
            .O(N__49325),
            .I(N__49224));
    InMux I__11551 (
            .O(N__49324),
            .I(N__49224));
    InMux I__11550 (
            .O(N__49323),
            .I(N__49224));
    InMux I__11549 (
            .O(N__49322),
            .I(N__49221));
    InMux I__11548 (
            .O(N__49319),
            .I(N__49216));
    InMux I__11547 (
            .O(N__49318),
            .I(N__49216));
    CascadeMux I__11546 (
            .O(N__49317),
            .I(N__49211));
    CascadeMux I__11545 (
            .O(N__49316),
            .I(N__49204));
    InMux I__11544 (
            .O(N__49313),
            .I(N__49200));
    InMux I__11543 (
            .O(N__49312),
            .I(N__49197));
    InMux I__11542 (
            .O(N__49311),
            .I(N__49194));
    InMux I__11541 (
            .O(N__49310),
            .I(N__49191));
    InMux I__11540 (
            .O(N__49309),
            .I(N__49188));
    LocalMux I__11539 (
            .O(N__49306),
            .I(N__49185));
    InMux I__11538 (
            .O(N__49305),
            .I(N__49180));
    InMux I__11537 (
            .O(N__49304),
            .I(N__49180));
    InMux I__11536 (
            .O(N__49303),
            .I(N__49173));
    InMux I__11535 (
            .O(N__49302),
            .I(N__49173));
    InMux I__11534 (
            .O(N__49301),
            .I(N__49173));
    LocalMux I__11533 (
            .O(N__49298),
            .I(N__49170));
    InMux I__11532 (
            .O(N__49297),
            .I(N__49167));
    InMux I__11531 (
            .O(N__49294),
            .I(N__49164));
    LocalMux I__11530 (
            .O(N__49291),
            .I(N__49159));
    LocalMux I__11529 (
            .O(N__49284),
            .I(N__49159));
    InMux I__11528 (
            .O(N__49281),
            .I(N__49156));
    InMux I__11527 (
            .O(N__49280),
            .I(N__49151));
    InMux I__11526 (
            .O(N__49279),
            .I(N__49151));
    Span4Mux_h I__11525 (
            .O(N__49276),
            .I(N__49148));
    InMux I__11524 (
            .O(N__49273),
            .I(N__49143));
    InMux I__11523 (
            .O(N__49272),
            .I(N__49143));
    LocalMux I__11522 (
            .O(N__49269),
            .I(N__49140));
    LocalMux I__11521 (
            .O(N__49264),
            .I(N__49135));
    Span4Mux_h I__11520 (
            .O(N__49259),
            .I(N__49135));
    CascadeMux I__11519 (
            .O(N__49258),
            .I(N__49128));
    InMux I__11518 (
            .O(N__49255),
            .I(N__49120));
    LocalMux I__11517 (
            .O(N__49252),
            .I(N__49113));
    LocalMux I__11516 (
            .O(N__49249),
            .I(N__49113));
    LocalMux I__11515 (
            .O(N__49244),
            .I(N__49113));
    CascadeMux I__11514 (
            .O(N__49243),
            .I(N__49109));
    CascadeMux I__11513 (
            .O(N__49242),
            .I(N__49105));
    Span4Mux_h I__11512 (
            .O(N__49239),
            .I(N__49100));
    InMux I__11511 (
            .O(N__49236),
            .I(N__49093));
    InMux I__11510 (
            .O(N__49235),
            .I(N__49093));
    InMux I__11509 (
            .O(N__49234),
            .I(N__49093));
    Span4Mux_v I__11508 (
            .O(N__49231),
            .I(N__49088));
    LocalMux I__11507 (
            .O(N__49224),
            .I(N__49088));
    LocalMux I__11506 (
            .O(N__49221),
            .I(N__49083));
    LocalMux I__11505 (
            .O(N__49216),
            .I(N__49083));
    InMux I__11504 (
            .O(N__49215),
            .I(N__49070));
    InMux I__11503 (
            .O(N__49214),
            .I(N__49070));
    InMux I__11502 (
            .O(N__49211),
            .I(N__49070));
    InMux I__11501 (
            .O(N__49210),
            .I(N__49070));
    InMux I__11500 (
            .O(N__49209),
            .I(N__49070));
    InMux I__11499 (
            .O(N__49208),
            .I(N__49070));
    InMux I__11498 (
            .O(N__49207),
            .I(N__49063));
    InMux I__11497 (
            .O(N__49204),
            .I(N__49063));
    InMux I__11496 (
            .O(N__49203),
            .I(N__49063));
    LocalMux I__11495 (
            .O(N__49200),
            .I(N__49056));
    LocalMux I__11494 (
            .O(N__49197),
            .I(N__49053));
    LocalMux I__11493 (
            .O(N__49194),
            .I(N__49050));
    LocalMux I__11492 (
            .O(N__49191),
            .I(N__49043));
    LocalMux I__11491 (
            .O(N__49188),
            .I(N__49043));
    Span4Mux_v I__11490 (
            .O(N__49185),
            .I(N__49043));
    LocalMux I__11489 (
            .O(N__49180),
            .I(N__49030));
    LocalMux I__11488 (
            .O(N__49173),
            .I(N__49030));
    Span4Mux_v I__11487 (
            .O(N__49170),
            .I(N__49030));
    LocalMux I__11486 (
            .O(N__49167),
            .I(N__49030));
    LocalMux I__11485 (
            .O(N__49164),
            .I(N__49030));
    Span4Mux_v I__11484 (
            .O(N__49159),
            .I(N__49030));
    LocalMux I__11483 (
            .O(N__49156),
            .I(N__49021));
    LocalMux I__11482 (
            .O(N__49151),
            .I(N__49021));
    Span4Mux_v I__11481 (
            .O(N__49148),
            .I(N__49021));
    LocalMux I__11480 (
            .O(N__49143),
            .I(N__49021));
    Span4Mux_h I__11479 (
            .O(N__49140),
            .I(N__49016));
    Span4Mux_h I__11478 (
            .O(N__49135),
            .I(N__49016));
    InMux I__11477 (
            .O(N__49134),
            .I(N__49013));
    InMux I__11476 (
            .O(N__49133),
            .I(N__49008));
    InMux I__11475 (
            .O(N__49132),
            .I(N__49008));
    InMux I__11474 (
            .O(N__49131),
            .I(N__48999));
    InMux I__11473 (
            .O(N__49128),
            .I(N__48999));
    InMux I__11472 (
            .O(N__49127),
            .I(N__48999));
    InMux I__11471 (
            .O(N__49126),
            .I(N__48999));
    InMux I__11470 (
            .O(N__49125),
            .I(N__48992));
    InMux I__11469 (
            .O(N__49124),
            .I(N__48992));
    InMux I__11468 (
            .O(N__49123),
            .I(N__48992));
    LocalMux I__11467 (
            .O(N__49120),
            .I(N__48987));
    Span4Mux_v I__11466 (
            .O(N__49113),
            .I(N__48987));
    InMux I__11465 (
            .O(N__49112),
            .I(N__48984));
    InMux I__11464 (
            .O(N__49109),
            .I(N__48973));
    InMux I__11463 (
            .O(N__49108),
            .I(N__48973));
    InMux I__11462 (
            .O(N__49105),
            .I(N__48973));
    InMux I__11461 (
            .O(N__49104),
            .I(N__48973));
    InMux I__11460 (
            .O(N__49103),
            .I(N__48973));
    Span4Mux_v I__11459 (
            .O(N__49100),
            .I(N__48966));
    LocalMux I__11458 (
            .O(N__49093),
            .I(N__48966));
    Span4Mux_h I__11457 (
            .O(N__49088),
            .I(N__48966));
    Span4Mux_v I__11456 (
            .O(N__49083),
            .I(N__48959));
    LocalMux I__11455 (
            .O(N__49070),
            .I(N__48959));
    LocalMux I__11454 (
            .O(N__49063),
            .I(N__48959));
    InMux I__11453 (
            .O(N__49062),
            .I(N__48956));
    InMux I__11452 (
            .O(N__49061),
            .I(N__48949));
    InMux I__11451 (
            .O(N__49060),
            .I(N__48949));
    InMux I__11450 (
            .O(N__49059),
            .I(N__48949));
    Span12Mux_h I__11449 (
            .O(N__49056),
            .I(N__48946));
    Span12Mux_v I__11448 (
            .O(N__49053),
            .I(N__48943));
    Span4Mux_v I__11447 (
            .O(N__49050),
            .I(N__48936));
    Span4Mux_v I__11446 (
            .O(N__49043),
            .I(N__48936));
    Span4Mux_h I__11445 (
            .O(N__49030),
            .I(N__48936));
    Span4Mux_h I__11444 (
            .O(N__49021),
            .I(N__48931));
    Span4Mux_v I__11443 (
            .O(N__49016),
            .I(N__48931));
    LocalMux I__11442 (
            .O(N__49013),
            .I(N__48926));
    LocalMux I__11441 (
            .O(N__49008),
            .I(N__48926));
    LocalMux I__11440 (
            .O(N__48999),
            .I(N__48913));
    LocalMux I__11439 (
            .O(N__48992),
            .I(N__48913));
    Span4Mux_h I__11438 (
            .O(N__48987),
            .I(N__48913));
    LocalMux I__11437 (
            .O(N__48984),
            .I(N__48913));
    LocalMux I__11436 (
            .O(N__48973),
            .I(N__48913));
    Span4Mux_v I__11435 (
            .O(N__48966),
            .I(N__48913));
    Span4Mux_h I__11434 (
            .O(N__48959),
            .I(N__48910));
    LocalMux I__11433 (
            .O(N__48956),
            .I(n9342));
    LocalMux I__11432 (
            .O(N__48949),
            .I(n9342));
    Odrv12 I__11431 (
            .O(N__48946),
            .I(n9342));
    Odrv12 I__11430 (
            .O(N__48943),
            .I(n9342));
    Odrv4 I__11429 (
            .O(N__48936),
            .I(n9342));
    Odrv4 I__11428 (
            .O(N__48931),
            .I(n9342));
    Odrv4 I__11427 (
            .O(N__48926),
            .I(n9342));
    Odrv4 I__11426 (
            .O(N__48913),
            .I(n9342));
    Odrv4 I__11425 (
            .O(N__48910),
            .I(n9342));
    InMux I__11424 (
            .O(N__48891),
            .I(N__48888));
    LocalMux I__11423 (
            .O(N__48888),
            .I(N__48885));
    Span4Mux_h I__11422 (
            .O(N__48885),
            .I(N__48882));
    Odrv4 I__11421 (
            .O(N__48882),
            .I(n18070));
    CEMux I__11420 (
            .O(N__48879),
            .I(N__48876));
    LocalMux I__11419 (
            .O(N__48876),
            .I(N__48873));
    Odrv12 I__11418 (
            .O(N__48873),
            .I(n21033));
    InMux I__11417 (
            .O(N__48870),
            .I(N__48867));
    LocalMux I__11416 (
            .O(N__48867),
            .I(N__48864));
    Span12Mux_v I__11415 (
            .O(N__48864),
            .I(N__48861));
    Odrv12 I__11414 (
            .O(N__48861),
            .I(n7_adj_1650));
    InMux I__11413 (
            .O(N__48858),
            .I(N__48855));
    LocalMux I__11412 (
            .O(N__48855),
            .I(N__48852));
    Span4Mux_h I__11411 (
            .O(N__48852),
            .I(N__48848));
    InMux I__11410 (
            .O(N__48851),
            .I(N__48844));
    Span4Mux_h I__11409 (
            .O(N__48848),
            .I(N__48841));
    InMux I__11408 (
            .O(N__48847),
            .I(N__48838));
    LocalMux I__11407 (
            .O(N__48844),
            .I(comm_cmd_6));
    Odrv4 I__11406 (
            .O(N__48841),
            .I(comm_cmd_6));
    LocalMux I__11405 (
            .O(N__48838),
            .I(comm_cmd_6));
    InMux I__11404 (
            .O(N__48831),
            .I(N__48828));
    LocalMux I__11403 (
            .O(N__48828),
            .I(N__48825));
    Span4Mux_h I__11402 (
            .O(N__48825),
            .I(N__48822));
    Span4Mux_h I__11401 (
            .O(N__48822),
            .I(N__48817));
    InMux I__11400 (
            .O(N__48821),
            .I(N__48812));
    InMux I__11399 (
            .O(N__48820),
            .I(N__48812));
    Odrv4 I__11398 (
            .O(N__48817),
            .I(comm_cmd_5));
    LocalMux I__11397 (
            .O(N__48812),
            .I(comm_cmd_5));
    InMux I__11396 (
            .O(N__48807),
            .I(N__48804));
    LocalMux I__11395 (
            .O(N__48804),
            .I(N__48801));
    Span4Mux_h I__11394 (
            .O(N__48801),
            .I(N__48798));
    Span4Mux_h I__11393 (
            .O(N__48798),
            .I(N__48795));
    Odrv4 I__11392 (
            .O(N__48795),
            .I(n4_adj_1455));
    InMux I__11391 (
            .O(N__48792),
            .I(N__48788));
    InMux I__11390 (
            .O(N__48791),
            .I(N__48785));
    LocalMux I__11389 (
            .O(N__48788),
            .I(N__48782));
    LocalMux I__11388 (
            .O(N__48785),
            .I(N__48779));
    Span4Mux_h I__11387 (
            .O(N__48782),
            .I(N__48776));
    Span4Mux_h I__11386 (
            .O(N__48779),
            .I(N__48773));
    Odrv4 I__11385 (
            .O(N__48776),
            .I(n21147));
    Odrv4 I__11384 (
            .O(N__48773),
            .I(n21147));
    CascadeMux I__11383 (
            .O(N__48768),
            .I(n21219_cascade_));
    InMux I__11382 (
            .O(N__48765),
            .I(N__48758));
    InMux I__11381 (
            .O(N__48764),
            .I(N__48758));
    InMux I__11380 (
            .O(N__48763),
            .I(N__48755));
    LocalMux I__11379 (
            .O(N__48758),
            .I(n21089));
    LocalMux I__11378 (
            .O(N__48755),
            .I(n21089));
    InMux I__11377 (
            .O(N__48750),
            .I(N__48746));
    InMux I__11376 (
            .O(N__48749),
            .I(N__48743));
    LocalMux I__11375 (
            .O(N__48746),
            .I(N__48738));
    LocalMux I__11374 (
            .O(N__48743),
            .I(N__48735));
    InMux I__11373 (
            .O(N__48742),
            .I(N__48732));
    InMux I__11372 (
            .O(N__48741),
            .I(N__48729));
    Odrv4 I__11371 (
            .O(N__48738),
            .I(n21043));
    Odrv4 I__11370 (
            .O(N__48735),
            .I(n21043));
    LocalMux I__11369 (
            .O(N__48732),
            .I(n21043));
    LocalMux I__11368 (
            .O(N__48729),
            .I(n21043));
    InMux I__11367 (
            .O(N__48720),
            .I(N__48717));
    LocalMux I__11366 (
            .O(N__48717),
            .I(N__48714));
    Span4Mux_h I__11365 (
            .O(N__48714),
            .I(N__48711));
    Odrv4 I__11364 (
            .O(N__48711),
            .I(buf_data_vac_16));
    InMux I__11363 (
            .O(N__48708),
            .I(N__48704));
    InMux I__11362 (
            .O(N__48707),
            .I(N__48700));
    LocalMux I__11361 (
            .O(N__48704),
            .I(N__48693));
    InMux I__11360 (
            .O(N__48703),
            .I(N__48690));
    LocalMux I__11359 (
            .O(N__48700),
            .I(N__48687));
    InMux I__11358 (
            .O(N__48699),
            .I(N__48684));
    InMux I__11357 (
            .O(N__48698),
            .I(N__48681));
    InMux I__11356 (
            .O(N__48697),
            .I(N__48678));
    InMux I__11355 (
            .O(N__48696),
            .I(N__48673));
    Span4Mux_h I__11354 (
            .O(N__48693),
            .I(N__48668));
    LocalMux I__11353 (
            .O(N__48690),
            .I(N__48668));
    Span4Mux_h I__11352 (
            .O(N__48687),
            .I(N__48659));
    LocalMux I__11351 (
            .O(N__48684),
            .I(N__48659));
    LocalMux I__11350 (
            .O(N__48681),
            .I(N__48659));
    LocalMux I__11349 (
            .O(N__48678),
            .I(N__48659));
    InMux I__11348 (
            .O(N__48677),
            .I(N__48656));
    InMux I__11347 (
            .O(N__48676),
            .I(N__48653));
    LocalMux I__11346 (
            .O(N__48673),
            .I(N__48650));
    Span4Mux_v I__11345 (
            .O(N__48668),
            .I(N__48645));
    Span4Mux_v I__11344 (
            .O(N__48659),
            .I(N__48645));
    LocalMux I__11343 (
            .O(N__48656),
            .I(N__48640));
    LocalMux I__11342 (
            .O(N__48653),
            .I(N__48640));
    Span4Mux_h I__11341 (
            .O(N__48650),
            .I(N__48635));
    Span4Mux_h I__11340 (
            .O(N__48645),
            .I(N__48635));
    Span12Mux_v I__11339 (
            .O(N__48640),
            .I(N__48632));
    Span4Mux_v I__11338 (
            .O(N__48635),
            .I(N__48629));
    Odrv12 I__11337 (
            .O(N__48632),
            .I(comm_rx_buf_0));
    Odrv4 I__11336 (
            .O(N__48629),
            .I(comm_rx_buf_0));
    CascadeMux I__11335 (
            .O(N__48624),
            .I(N__48621));
    InMux I__11334 (
            .O(N__48621),
            .I(N__48618));
    LocalMux I__11333 (
            .O(N__48618),
            .I(comm_buf_3_0));
    InMux I__11332 (
            .O(N__48615),
            .I(N__48612));
    LocalMux I__11331 (
            .O(N__48612),
            .I(N__48609));
    Sp12to4 I__11330 (
            .O(N__48609),
            .I(N__48606));
    Span12Mux_v I__11329 (
            .O(N__48606),
            .I(N__48603));
    Odrv12 I__11328 (
            .O(N__48603),
            .I(buf_data_vac_23));
    InMux I__11327 (
            .O(N__48600),
            .I(N__48592));
    InMux I__11326 (
            .O(N__48599),
            .I(N__48589));
    CascadeMux I__11325 (
            .O(N__48598),
            .I(N__48585));
    CascadeMux I__11324 (
            .O(N__48597),
            .I(N__48582));
    CascadeMux I__11323 (
            .O(N__48596),
            .I(N__48579));
    InMux I__11322 (
            .O(N__48595),
            .I(N__48576));
    LocalMux I__11321 (
            .O(N__48592),
            .I(N__48573));
    LocalMux I__11320 (
            .O(N__48589),
            .I(N__48569));
    InMux I__11319 (
            .O(N__48588),
            .I(N__48566));
    InMux I__11318 (
            .O(N__48585),
            .I(N__48563));
    InMux I__11317 (
            .O(N__48582),
            .I(N__48560));
    InMux I__11316 (
            .O(N__48579),
            .I(N__48557));
    LocalMux I__11315 (
            .O(N__48576),
            .I(N__48554));
    Span4Mux_v I__11314 (
            .O(N__48573),
            .I(N__48551));
    InMux I__11313 (
            .O(N__48572),
            .I(N__48548));
    Span4Mux_v I__11312 (
            .O(N__48569),
            .I(N__48543));
    LocalMux I__11311 (
            .O(N__48566),
            .I(N__48543));
    LocalMux I__11310 (
            .O(N__48563),
            .I(N__48540));
    LocalMux I__11309 (
            .O(N__48560),
            .I(N__48535));
    LocalMux I__11308 (
            .O(N__48557),
            .I(N__48535));
    Span4Mux_h I__11307 (
            .O(N__48554),
            .I(N__48528));
    Span4Mux_h I__11306 (
            .O(N__48551),
            .I(N__48528));
    LocalMux I__11305 (
            .O(N__48548),
            .I(N__48528));
    Span4Mux_v I__11304 (
            .O(N__48543),
            .I(N__48525));
    Span4Mux_v I__11303 (
            .O(N__48540),
            .I(N__48520));
    Span4Mux_v I__11302 (
            .O(N__48535),
            .I(N__48520));
    Span4Mux_v I__11301 (
            .O(N__48528),
            .I(N__48517));
    Odrv4 I__11300 (
            .O(N__48525),
            .I(comm_rx_buf_7));
    Odrv4 I__11299 (
            .O(N__48520),
            .I(comm_rx_buf_7));
    Odrv4 I__11298 (
            .O(N__48517),
            .I(comm_rx_buf_7));
    CascadeMux I__11297 (
            .O(N__48510),
            .I(N__48507));
    InMux I__11296 (
            .O(N__48507),
            .I(N__48504));
    LocalMux I__11295 (
            .O(N__48504),
            .I(N__48501));
    Span4Mux_h I__11294 (
            .O(N__48501),
            .I(N__48498));
    Span4Mux_h I__11293 (
            .O(N__48498),
            .I(N__48495));
    Odrv4 I__11292 (
            .O(N__48495),
            .I(comm_buf_3_7));
    InMux I__11291 (
            .O(N__48492),
            .I(N__48489));
    LocalMux I__11290 (
            .O(N__48489),
            .I(N__48486));
    Sp12to4 I__11289 (
            .O(N__48486),
            .I(N__48483));
    Span12Mux_v I__11288 (
            .O(N__48483),
            .I(N__48480));
    Odrv12 I__11287 (
            .O(N__48480),
            .I(buf_data_vac_22));
    InMux I__11286 (
            .O(N__48477),
            .I(N__48474));
    LocalMux I__11285 (
            .O(N__48474),
            .I(N__48471));
    Span4Mux_v I__11284 (
            .O(N__48471),
            .I(N__48468));
    Span4Mux_v I__11283 (
            .O(N__48468),
            .I(N__48465));
    Odrv4 I__11282 (
            .O(N__48465),
            .I(buf_data_vac_21));
    InMux I__11281 (
            .O(N__48462),
            .I(N__48459));
    LocalMux I__11280 (
            .O(N__48459),
            .I(n4));
    CascadeMux I__11279 (
            .O(N__48456),
            .I(n21013_cascade_));
    CEMux I__11278 (
            .O(N__48453),
            .I(N__48450));
    LocalMux I__11277 (
            .O(N__48450),
            .I(N__48447));
    Odrv4 I__11276 (
            .O(N__48447),
            .I(n21035));
    CascadeMux I__11275 (
            .O(N__48444),
            .I(N__48441));
    InMux I__11274 (
            .O(N__48441),
            .I(N__48438));
    LocalMux I__11273 (
            .O(N__48438),
            .I(N__48435));
    Span4Mux_v I__11272 (
            .O(N__48435),
            .I(N__48432));
    Odrv4 I__11271 (
            .O(N__48432),
            .I(comm_length_0));
    InMux I__11270 (
            .O(N__48429),
            .I(N__48426));
    LocalMux I__11269 (
            .O(N__48426),
            .I(N__48423));
    Span4Mux_v I__11268 (
            .O(N__48423),
            .I(N__48420));
    Odrv4 I__11267 (
            .O(N__48420),
            .I(n4_adj_1623));
    InMux I__11266 (
            .O(N__48417),
            .I(N__48414));
    LocalMux I__11265 (
            .O(N__48414),
            .I(n3));
    InMux I__11264 (
            .O(N__48411),
            .I(N__48404));
    InMux I__11263 (
            .O(N__48410),
            .I(N__48401));
    InMux I__11262 (
            .O(N__48409),
            .I(N__48398));
    CascadeMux I__11261 (
            .O(N__48408),
            .I(N__48395));
    InMux I__11260 (
            .O(N__48407),
            .I(N__48392));
    LocalMux I__11259 (
            .O(N__48404),
            .I(N__48389));
    LocalMux I__11258 (
            .O(N__48401),
            .I(N__48384));
    LocalMux I__11257 (
            .O(N__48398),
            .I(N__48384));
    InMux I__11256 (
            .O(N__48395),
            .I(N__48381));
    LocalMux I__11255 (
            .O(N__48392),
            .I(N__48378));
    Span4Mux_v I__11254 (
            .O(N__48389),
            .I(N__48375));
    Span4Mux_v I__11253 (
            .O(N__48384),
            .I(N__48370));
    LocalMux I__11252 (
            .O(N__48381),
            .I(N__48370));
    Odrv12 I__11251 (
            .O(N__48378),
            .I(n21110));
    Odrv4 I__11250 (
            .O(N__48375),
            .I(n21110));
    Odrv4 I__11249 (
            .O(N__48370),
            .I(n21110));
    CascadeMux I__11248 (
            .O(N__48363),
            .I(n3_cascade_));
    InMux I__11247 (
            .O(N__48360),
            .I(N__48355));
    InMux I__11246 (
            .O(N__48359),
            .I(N__48350));
    InMux I__11245 (
            .O(N__48358),
            .I(N__48350));
    LocalMux I__11244 (
            .O(N__48355),
            .I(N__48345));
    LocalMux I__11243 (
            .O(N__48350),
            .I(N__48345));
    Span4Mux_h I__11242 (
            .O(N__48345),
            .I(N__48342));
    Span4Mux_h I__11241 (
            .O(N__48342),
            .I(N__48338));
    InMux I__11240 (
            .O(N__48341),
            .I(N__48335));
    Odrv4 I__11239 (
            .O(N__48338),
            .I(n12442));
    LocalMux I__11238 (
            .O(N__48335),
            .I(n12442));
    InMux I__11237 (
            .O(N__48330),
            .I(N__48327));
    LocalMux I__11236 (
            .O(N__48327),
            .I(n4_adj_1589));
    CascadeMux I__11235 (
            .O(N__48324),
            .I(n20095_cascade_));
    InMux I__11234 (
            .O(N__48321),
            .I(N__48318));
    LocalMux I__11233 (
            .O(N__48318),
            .I(n21013));
    InMux I__11232 (
            .O(N__48315),
            .I(N__48312));
    LocalMux I__11231 (
            .O(N__48312),
            .I(n11619));
    CascadeMux I__11230 (
            .O(N__48309),
            .I(N__48306));
    InMux I__11229 (
            .O(N__48306),
            .I(N__48303));
    LocalMux I__11228 (
            .O(N__48303),
            .I(N__48300));
    Odrv4 I__11227 (
            .O(N__48300),
            .I(buf_data_vac_1));
    CEMux I__11226 (
            .O(N__48297),
            .I(N__48294));
    LocalMux I__11225 (
            .O(N__48294),
            .I(N__48290));
    InMux I__11224 (
            .O(N__48293),
            .I(N__48287));
    Span4Mux_h I__11223 (
            .O(N__48290),
            .I(N__48284));
    LocalMux I__11222 (
            .O(N__48287),
            .I(N__48281));
    Odrv4 I__11221 (
            .O(N__48284),
            .I(n12431));
    Odrv4 I__11220 (
            .O(N__48281),
            .I(n12431));
    SRMux I__11219 (
            .O(N__48276),
            .I(N__48273));
    LocalMux I__11218 (
            .O(N__48273),
            .I(N__48270));
    Odrv4 I__11217 (
            .O(N__48270),
            .I(n14993));
    InMux I__11216 (
            .O(N__48267),
            .I(N__48263));
    InMux I__11215 (
            .O(N__48266),
            .I(N__48260));
    LocalMux I__11214 (
            .O(N__48263),
            .I(N__48254));
    LocalMux I__11213 (
            .O(N__48260),
            .I(N__48251));
    InMux I__11212 (
            .O(N__48259),
            .I(N__48248));
    InMux I__11211 (
            .O(N__48258),
            .I(N__48245));
    InMux I__11210 (
            .O(N__48257),
            .I(N__48242));
    Span4Mux_h I__11209 (
            .O(N__48254),
            .I(N__48238));
    Span4Mux_h I__11208 (
            .O(N__48251),
            .I(N__48232));
    LocalMux I__11207 (
            .O(N__48248),
            .I(N__48232));
    LocalMux I__11206 (
            .O(N__48245),
            .I(N__48229));
    LocalMux I__11205 (
            .O(N__48242),
            .I(N__48226));
    InMux I__11204 (
            .O(N__48241),
            .I(N__48223));
    Span4Mux_h I__11203 (
            .O(N__48238),
            .I(N__48220));
    InMux I__11202 (
            .O(N__48237),
            .I(N__48217));
    Span4Mux_v I__11201 (
            .O(N__48232),
            .I(N__48208));
    Span4Mux_v I__11200 (
            .O(N__48229),
            .I(N__48208));
    Span4Mux_h I__11199 (
            .O(N__48226),
            .I(N__48208));
    LocalMux I__11198 (
            .O(N__48223),
            .I(N__48208));
    Odrv4 I__11197 (
            .O(N__48220),
            .I(n11652));
    LocalMux I__11196 (
            .O(N__48217),
            .I(n11652));
    Odrv4 I__11195 (
            .O(N__48208),
            .I(n11652));
    CascadeMux I__11194 (
            .O(N__48201),
            .I(n2_adj_1576_cascade_));
    InMux I__11193 (
            .O(N__48198),
            .I(N__48195));
    LocalMux I__11192 (
            .O(N__48195),
            .I(n22611));
    InMux I__11191 (
            .O(N__48192),
            .I(N__48189));
    LocalMux I__11190 (
            .O(N__48189),
            .I(N__48185));
    InMux I__11189 (
            .O(N__48188),
            .I(N__48182));
    Span4Mux_v I__11188 (
            .O(N__48185),
            .I(N__48177));
    LocalMux I__11187 (
            .O(N__48182),
            .I(N__48177));
    Span4Mux_h I__11186 (
            .O(N__48177),
            .I(N__48174));
    Span4Mux_h I__11185 (
            .O(N__48174),
            .I(N__48171));
    Odrv4 I__11184 (
            .O(N__48171),
            .I(comm_state_3_N_460_3));
    CascadeMux I__11183 (
            .O(N__48168),
            .I(n1348_cascade_));
    CascadeMux I__11182 (
            .O(N__48165),
            .I(n21139_cascade_));
    InMux I__11181 (
            .O(N__48162),
            .I(N__48156));
    InMux I__11180 (
            .O(N__48161),
            .I(N__48156));
    LocalMux I__11179 (
            .O(N__48156),
            .I(n1348));
    InMux I__11178 (
            .O(N__48153),
            .I(N__48150));
    LocalMux I__11177 (
            .O(N__48150),
            .I(n8_adj_1577));
    InMux I__11176 (
            .O(N__48147),
            .I(N__48144));
    LocalMux I__11175 (
            .O(N__48144),
            .I(n22614));
    InMux I__11174 (
            .O(N__48141),
            .I(N__48134));
    InMux I__11173 (
            .O(N__48140),
            .I(N__48131));
    InMux I__11172 (
            .O(N__48139),
            .I(N__48128));
    InMux I__11171 (
            .O(N__48138),
            .I(N__48125));
    InMux I__11170 (
            .O(N__48137),
            .I(N__48122));
    LocalMux I__11169 (
            .O(N__48134),
            .I(N__48117));
    LocalMux I__11168 (
            .O(N__48131),
            .I(N__48117));
    LocalMux I__11167 (
            .O(N__48128),
            .I(N__48110));
    LocalMux I__11166 (
            .O(N__48125),
            .I(N__48110));
    LocalMux I__11165 (
            .O(N__48122),
            .I(N__48110));
    Span4Mux_v I__11164 (
            .O(N__48117),
            .I(N__48107));
    Span4Mux_v I__11163 (
            .O(N__48110),
            .I(N__48104));
    Sp12to4 I__11162 (
            .O(N__48107),
            .I(N__48099));
    Sp12to4 I__11161 (
            .O(N__48104),
            .I(N__48099));
    Span12Mux_h I__11160 (
            .O(N__48099),
            .I(N__48096));
    Span12Mux_v I__11159 (
            .O(N__48096),
            .I(N__48093));
    Odrv12 I__11158 (
            .O(N__48093),
            .I(ICE_SPI_SCLK));
    SRMux I__11157 (
            .O(N__48090),
            .I(N__48087));
    LocalMux I__11156 (
            .O(N__48087),
            .I(N__48084));
    Span4Mux_v I__11155 (
            .O(N__48084),
            .I(N__48081));
    Odrv4 I__11154 (
            .O(N__48081),
            .I(\comm_spi.iclk_N_803 ));
    InMux I__11153 (
            .O(N__48078),
            .I(N__48075));
    LocalMux I__11152 (
            .O(N__48075),
            .I(N__48072));
    Span4Mux_h I__11151 (
            .O(N__48072),
            .I(N__48069));
    Odrv4 I__11150 (
            .O(N__48069),
            .I(buf_data_vac_0));
    InMux I__11149 (
            .O(N__48066),
            .I(N__48063));
    LocalMux I__11148 (
            .O(N__48063),
            .I(N__48060));
    Span4Mux_v I__11147 (
            .O(N__48060),
            .I(N__48057));
    Span4Mux_h I__11146 (
            .O(N__48057),
            .I(N__48054));
    Sp12to4 I__11145 (
            .O(N__48054),
            .I(N__48051));
    Odrv12 I__11144 (
            .O(N__48051),
            .I(buf_data_vac_7));
    InMux I__11143 (
            .O(N__48048),
            .I(N__48045));
    LocalMux I__11142 (
            .O(N__48045),
            .I(N__48042));
    Span4Mux_h I__11141 (
            .O(N__48042),
            .I(N__48039));
    Odrv4 I__11140 (
            .O(N__48039),
            .I(comm_buf_5_7));
    InMux I__11139 (
            .O(N__48036),
            .I(N__48033));
    LocalMux I__11138 (
            .O(N__48033),
            .I(N__48030));
    Span12Mux_v I__11137 (
            .O(N__48030),
            .I(N__48027));
    Span12Mux_h I__11136 (
            .O(N__48027),
            .I(N__48024));
    Odrv12 I__11135 (
            .O(N__48024),
            .I(buf_data_vac_6));
    InMux I__11134 (
            .O(N__48021),
            .I(N__48018));
    LocalMux I__11133 (
            .O(N__48018),
            .I(N__48015));
    Span4Mux_h I__11132 (
            .O(N__48015),
            .I(N__48012));
    Span4Mux_h I__11131 (
            .O(N__48012),
            .I(N__48009));
    Span4Mux_h I__11130 (
            .O(N__48009),
            .I(N__48006));
    Odrv4 I__11129 (
            .O(N__48006),
            .I(buf_data_vac_5));
    InMux I__11128 (
            .O(N__48003),
            .I(N__48000));
    LocalMux I__11127 (
            .O(N__48000),
            .I(N__47997));
    Span4Mux_v I__11126 (
            .O(N__47997),
            .I(N__47994));
    Span4Mux_h I__11125 (
            .O(N__47994),
            .I(N__47991));
    Sp12to4 I__11124 (
            .O(N__47991),
            .I(N__47988));
    Odrv12 I__11123 (
            .O(N__47988),
            .I(buf_data_vac_4));
    InMux I__11122 (
            .O(N__47985),
            .I(N__47982));
    LocalMux I__11121 (
            .O(N__47982),
            .I(N__47979));
    Span4Mux_h I__11120 (
            .O(N__47979),
            .I(N__47976));
    Odrv4 I__11119 (
            .O(N__47976),
            .I(comm_buf_5_4));
    InMux I__11118 (
            .O(N__47973),
            .I(N__47970));
    LocalMux I__11117 (
            .O(N__47970),
            .I(N__47967));
    Span4Mux_h I__11116 (
            .O(N__47967),
            .I(N__47964));
    Odrv4 I__11115 (
            .O(N__47964),
            .I(buf_data_vac_3));
    CascadeMux I__11114 (
            .O(N__47961),
            .I(N__47958));
    InMux I__11113 (
            .O(N__47958),
            .I(N__47955));
    LocalMux I__11112 (
            .O(N__47955),
            .I(N__47952));
    Odrv4 I__11111 (
            .O(N__47952),
            .I(comm_buf_5_3));
    InMux I__11110 (
            .O(N__47949),
            .I(N__47946));
    LocalMux I__11109 (
            .O(N__47946),
            .I(N__47943));
    Span4Mux_v I__11108 (
            .O(N__47943),
            .I(N__47940));
    Odrv4 I__11107 (
            .O(N__47940),
            .I(buf_data_vac_2));
    InMux I__11106 (
            .O(N__47937),
            .I(N__47934));
    LocalMux I__11105 (
            .O(N__47934),
            .I(N__47931));
    Span4Mux_v I__11104 (
            .O(N__47931),
            .I(N__47928));
    Odrv4 I__11103 (
            .O(N__47928),
            .I(comm_buf_5_2));
    InMux I__11102 (
            .O(N__47925),
            .I(N__47917));
    InMux I__11101 (
            .O(N__47924),
            .I(N__47911));
    InMux I__11100 (
            .O(N__47923),
            .I(N__47911));
    CascadeMux I__11099 (
            .O(N__47922),
            .I(N__47902));
    CascadeMux I__11098 (
            .O(N__47921),
            .I(N__47899));
    InMux I__11097 (
            .O(N__47920),
            .I(N__47896));
    LocalMux I__11096 (
            .O(N__47917),
            .I(N__47893));
    InMux I__11095 (
            .O(N__47916),
            .I(N__47890));
    LocalMux I__11094 (
            .O(N__47911),
            .I(N__47887));
    InMux I__11093 (
            .O(N__47910),
            .I(N__47882));
    InMux I__11092 (
            .O(N__47909),
            .I(N__47882));
    InMux I__11091 (
            .O(N__47908),
            .I(N__47873));
    InMux I__11090 (
            .O(N__47907),
            .I(N__47873));
    InMux I__11089 (
            .O(N__47906),
            .I(N__47873));
    InMux I__11088 (
            .O(N__47905),
            .I(N__47873));
    InMux I__11087 (
            .O(N__47902),
            .I(N__47868));
    InMux I__11086 (
            .O(N__47899),
            .I(N__47868));
    LocalMux I__11085 (
            .O(N__47896),
            .I(N__47865));
    Span4Mux_h I__11084 (
            .O(N__47893),
            .I(N__47859));
    LocalMux I__11083 (
            .O(N__47890),
            .I(N__47856));
    Span4Mux_v I__11082 (
            .O(N__47887),
            .I(N__47847));
    LocalMux I__11081 (
            .O(N__47882),
            .I(N__47847));
    LocalMux I__11080 (
            .O(N__47873),
            .I(N__47847));
    LocalMux I__11079 (
            .O(N__47868),
            .I(N__47847));
    Span12Mux_v I__11078 (
            .O(N__47865),
            .I(N__47844));
    InMux I__11077 (
            .O(N__47864),
            .I(N__47841));
    InMux I__11076 (
            .O(N__47863),
            .I(N__47836));
    InMux I__11075 (
            .O(N__47862),
            .I(N__47836));
    Span4Mux_h I__11074 (
            .O(N__47859),
            .I(N__47829));
    Span4Mux_v I__11073 (
            .O(N__47856),
            .I(N__47829));
    Span4Mux_v I__11072 (
            .O(N__47847),
            .I(N__47829));
    Odrv12 I__11071 (
            .O(N__47844),
            .I(n12654));
    LocalMux I__11070 (
            .O(N__47841),
            .I(n12654));
    LocalMux I__11069 (
            .O(N__47836),
            .I(n12654));
    Odrv4 I__11068 (
            .O(N__47829),
            .I(n12654));
    CascadeMux I__11067 (
            .O(N__47820),
            .I(N__47816));
    CascadeMux I__11066 (
            .O(N__47819),
            .I(N__47812));
    InMux I__11065 (
            .O(N__47816),
            .I(N__47809));
    CascadeMux I__11064 (
            .O(N__47815),
            .I(N__47806));
    InMux I__11063 (
            .O(N__47812),
            .I(N__47803));
    LocalMux I__11062 (
            .O(N__47809),
            .I(N__47800));
    InMux I__11061 (
            .O(N__47806),
            .I(N__47796));
    LocalMux I__11060 (
            .O(N__47803),
            .I(N__47791));
    Span4Mux_v I__11059 (
            .O(N__47800),
            .I(N__47791));
    InMux I__11058 (
            .O(N__47799),
            .I(N__47788));
    LocalMux I__11057 (
            .O(N__47796),
            .I(N__47783));
    Span4Mux_v I__11056 (
            .O(N__47791),
            .I(N__47778));
    LocalMux I__11055 (
            .O(N__47788),
            .I(N__47778));
    InMux I__11054 (
            .O(N__47787),
            .I(N__47775));
    InMux I__11053 (
            .O(N__47786),
            .I(N__47771));
    Span4Mux_v I__11052 (
            .O(N__47783),
            .I(N__47768));
    Span4Mux_v I__11051 (
            .O(N__47778),
            .I(N__47763));
    LocalMux I__11050 (
            .O(N__47775),
            .I(N__47763));
    InMux I__11049 (
            .O(N__47774),
            .I(N__47760));
    LocalMux I__11048 (
            .O(N__47771),
            .I(N__47756));
    Span4Mux_v I__11047 (
            .O(N__47768),
            .I(N__47751));
    Span4Mux_h I__11046 (
            .O(N__47763),
            .I(N__47751));
    LocalMux I__11045 (
            .O(N__47760),
            .I(N__47748));
    InMux I__11044 (
            .O(N__47759),
            .I(N__47745));
    Span4Mux_h I__11043 (
            .O(N__47756),
            .I(N__47742));
    Odrv4 I__11042 (
            .O(N__47751),
            .I(comm_buf_0_4));
    Odrv12 I__11041 (
            .O(N__47748),
            .I(comm_buf_0_4));
    LocalMux I__11040 (
            .O(N__47745),
            .I(comm_buf_0_4));
    Odrv4 I__11039 (
            .O(N__47742),
            .I(comm_buf_0_4));
    InMux I__11038 (
            .O(N__47733),
            .I(N__47730));
    LocalMux I__11037 (
            .O(N__47730),
            .I(N__47725));
    InMux I__11036 (
            .O(N__47729),
            .I(N__47718));
    CascadeMux I__11035 (
            .O(N__47728),
            .I(N__47713));
    Span4Mux_h I__11034 (
            .O(N__47725),
            .I(N__47688));
    InMux I__11033 (
            .O(N__47724),
            .I(N__47679));
    InMux I__11032 (
            .O(N__47723),
            .I(N__47679));
    InMux I__11031 (
            .O(N__47722),
            .I(N__47679));
    InMux I__11030 (
            .O(N__47721),
            .I(N__47679));
    LocalMux I__11029 (
            .O(N__47718),
            .I(N__47668));
    InMux I__11028 (
            .O(N__47717),
            .I(N__47658));
    InMux I__11027 (
            .O(N__47716),
            .I(N__47649));
    InMux I__11026 (
            .O(N__47713),
            .I(N__47649));
    InMux I__11025 (
            .O(N__47712),
            .I(N__47649));
    InMux I__11024 (
            .O(N__47711),
            .I(N__47649));
    InMux I__11023 (
            .O(N__47710),
            .I(N__47644));
    InMux I__11022 (
            .O(N__47709),
            .I(N__47644));
    CascadeMux I__11021 (
            .O(N__47708),
            .I(N__47639));
    InMux I__11020 (
            .O(N__47707),
            .I(N__47628));
    InMux I__11019 (
            .O(N__47706),
            .I(N__47628));
    InMux I__11018 (
            .O(N__47705),
            .I(N__47628));
    InMux I__11017 (
            .O(N__47704),
            .I(N__47628));
    InMux I__11016 (
            .O(N__47703),
            .I(N__47625));
    InMux I__11015 (
            .O(N__47702),
            .I(N__47622));
    InMux I__11014 (
            .O(N__47701),
            .I(N__47613));
    InMux I__11013 (
            .O(N__47700),
            .I(N__47613));
    InMux I__11012 (
            .O(N__47699),
            .I(N__47613));
    InMux I__11011 (
            .O(N__47698),
            .I(N__47613));
    InMux I__11010 (
            .O(N__47697),
            .I(N__47608));
    InMux I__11009 (
            .O(N__47696),
            .I(N__47608));
    InMux I__11008 (
            .O(N__47695),
            .I(N__47605));
    InMux I__11007 (
            .O(N__47694),
            .I(N__47602));
    InMux I__11006 (
            .O(N__47693),
            .I(N__47594));
    InMux I__11005 (
            .O(N__47692),
            .I(N__47594));
    InMux I__11004 (
            .O(N__47691),
            .I(N__47594));
    Span4Mux_v I__11003 (
            .O(N__47688),
            .I(N__47589));
    LocalMux I__11002 (
            .O(N__47679),
            .I(N__47589));
    InMux I__11001 (
            .O(N__47678),
            .I(N__47578));
    InMux I__11000 (
            .O(N__47677),
            .I(N__47578));
    InMux I__10999 (
            .O(N__47676),
            .I(N__47578));
    InMux I__10998 (
            .O(N__47675),
            .I(N__47578));
    InMux I__10997 (
            .O(N__47674),
            .I(N__47578));
    InMux I__10996 (
            .O(N__47673),
            .I(N__47571));
    InMux I__10995 (
            .O(N__47672),
            .I(N__47571));
    InMux I__10994 (
            .O(N__47671),
            .I(N__47571));
    Span4Mux_h I__10993 (
            .O(N__47668),
            .I(N__47568));
    InMux I__10992 (
            .O(N__47667),
            .I(N__47565));
    InMux I__10991 (
            .O(N__47666),
            .I(N__47560));
    InMux I__10990 (
            .O(N__47665),
            .I(N__47557));
    InMux I__10989 (
            .O(N__47664),
            .I(N__47548));
    InMux I__10988 (
            .O(N__47663),
            .I(N__47548));
    InMux I__10987 (
            .O(N__47662),
            .I(N__47548));
    InMux I__10986 (
            .O(N__47661),
            .I(N__47548));
    LocalMux I__10985 (
            .O(N__47658),
            .I(N__47541));
    LocalMux I__10984 (
            .O(N__47649),
            .I(N__47541));
    LocalMux I__10983 (
            .O(N__47644),
            .I(N__47541));
    InMux I__10982 (
            .O(N__47643),
            .I(N__47538));
    InMux I__10981 (
            .O(N__47642),
            .I(N__47533));
    InMux I__10980 (
            .O(N__47639),
            .I(N__47524));
    InMux I__10979 (
            .O(N__47638),
            .I(N__47524));
    InMux I__10978 (
            .O(N__47637),
            .I(N__47521));
    LocalMux I__10977 (
            .O(N__47628),
            .I(N__47510));
    LocalMux I__10976 (
            .O(N__47625),
            .I(N__47510));
    LocalMux I__10975 (
            .O(N__47622),
            .I(N__47507));
    LocalMux I__10974 (
            .O(N__47613),
            .I(N__47502));
    LocalMux I__10973 (
            .O(N__47608),
            .I(N__47502));
    LocalMux I__10972 (
            .O(N__47605),
            .I(N__47495));
    LocalMux I__10971 (
            .O(N__47602),
            .I(N__47495));
    InMux I__10970 (
            .O(N__47601),
            .I(N__47492));
    LocalMux I__10969 (
            .O(N__47594),
            .I(N__47485));
    Span4Mux_v I__10968 (
            .O(N__47589),
            .I(N__47485));
    LocalMux I__10967 (
            .O(N__47578),
            .I(N__47485));
    LocalMux I__10966 (
            .O(N__47571),
            .I(N__47478));
    Span4Mux_h I__10965 (
            .O(N__47568),
            .I(N__47478));
    LocalMux I__10964 (
            .O(N__47565),
            .I(N__47478));
    InMux I__10963 (
            .O(N__47564),
            .I(N__47473));
    InMux I__10962 (
            .O(N__47563),
            .I(N__47473));
    LocalMux I__10961 (
            .O(N__47560),
            .I(N__47468));
    LocalMux I__10960 (
            .O(N__47557),
            .I(N__47468));
    LocalMux I__10959 (
            .O(N__47548),
            .I(N__47461));
    Span4Mux_v I__10958 (
            .O(N__47541),
            .I(N__47461));
    LocalMux I__10957 (
            .O(N__47538),
            .I(N__47461));
    CascadeMux I__10956 (
            .O(N__47537),
            .I(N__47458));
    InMux I__10955 (
            .O(N__47536),
            .I(N__47454));
    LocalMux I__10954 (
            .O(N__47533),
            .I(N__47446));
    InMux I__10953 (
            .O(N__47532),
            .I(N__47443));
    InMux I__10952 (
            .O(N__47531),
            .I(N__47436));
    InMux I__10951 (
            .O(N__47530),
            .I(N__47436));
    InMux I__10950 (
            .O(N__47529),
            .I(N__47436));
    LocalMux I__10949 (
            .O(N__47524),
            .I(N__47431));
    LocalMux I__10948 (
            .O(N__47521),
            .I(N__47431));
    InMux I__10947 (
            .O(N__47520),
            .I(N__47424));
    InMux I__10946 (
            .O(N__47519),
            .I(N__47424));
    InMux I__10945 (
            .O(N__47518),
            .I(N__47424));
    InMux I__10944 (
            .O(N__47517),
            .I(N__47419));
    InMux I__10943 (
            .O(N__47516),
            .I(N__47419));
    InMux I__10942 (
            .O(N__47515),
            .I(N__47416));
    Span4Mux_v I__10941 (
            .O(N__47510),
            .I(N__47409));
    Span4Mux_v I__10940 (
            .O(N__47507),
            .I(N__47409));
    Span4Mux_v I__10939 (
            .O(N__47502),
            .I(N__47409));
    InMux I__10938 (
            .O(N__47501),
            .I(N__47404));
    InMux I__10937 (
            .O(N__47500),
            .I(N__47404));
    Span4Mux_h I__10936 (
            .O(N__47495),
            .I(N__47397));
    LocalMux I__10935 (
            .O(N__47492),
            .I(N__47397));
    Span4Mux_h I__10934 (
            .O(N__47485),
            .I(N__47397));
    Span4Mux_v I__10933 (
            .O(N__47478),
            .I(N__47394));
    LocalMux I__10932 (
            .O(N__47473),
            .I(N__47387));
    Span4Mux_v I__10931 (
            .O(N__47468),
            .I(N__47387));
    Span4Mux_h I__10930 (
            .O(N__47461),
            .I(N__47387));
    InMux I__10929 (
            .O(N__47458),
            .I(N__47384));
    InMux I__10928 (
            .O(N__47457),
            .I(N__47381));
    LocalMux I__10927 (
            .O(N__47454),
            .I(N__47378));
    InMux I__10926 (
            .O(N__47453),
            .I(N__47375));
    InMux I__10925 (
            .O(N__47452),
            .I(N__47370));
    InMux I__10924 (
            .O(N__47451),
            .I(N__47370));
    InMux I__10923 (
            .O(N__47450),
            .I(N__47365));
    InMux I__10922 (
            .O(N__47449),
            .I(N__47365));
    Span12Mux_h I__10921 (
            .O(N__47446),
            .I(N__47360));
    LocalMux I__10920 (
            .O(N__47443),
            .I(N__47360));
    LocalMux I__10919 (
            .O(N__47436),
            .I(N__47347));
    Span12Mux_v I__10918 (
            .O(N__47431),
            .I(N__47347));
    LocalMux I__10917 (
            .O(N__47424),
            .I(N__47347));
    LocalMux I__10916 (
            .O(N__47419),
            .I(N__47347));
    LocalMux I__10915 (
            .O(N__47416),
            .I(N__47347));
    Sp12to4 I__10914 (
            .O(N__47409),
            .I(N__47347));
    LocalMux I__10913 (
            .O(N__47404),
            .I(N__47342));
    Span4Mux_h I__10912 (
            .O(N__47397),
            .I(N__47342));
    Span4Mux_h I__10911 (
            .O(N__47394),
            .I(N__47337));
    Span4Mux_h I__10910 (
            .O(N__47387),
            .I(N__47337));
    LocalMux I__10909 (
            .O(N__47384),
            .I(comm_cmd_2));
    LocalMux I__10908 (
            .O(N__47381),
            .I(comm_cmd_2));
    Odrv4 I__10907 (
            .O(N__47378),
            .I(comm_cmd_2));
    LocalMux I__10906 (
            .O(N__47375),
            .I(comm_cmd_2));
    LocalMux I__10905 (
            .O(N__47370),
            .I(comm_cmd_2));
    LocalMux I__10904 (
            .O(N__47365),
            .I(comm_cmd_2));
    Odrv12 I__10903 (
            .O(N__47360),
            .I(comm_cmd_2));
    Odrv12 I__10902 (
            .O(N__47347),
            .I(comm_cmd_2));
    Odrv4 I__10901 (
            .O(N__47342),
            .I(comm_cmd_2));
    Odrv4 I__10900 (
            .O(N__47337),
            .I(comm_cmd_2));
    CascadeMux I__10899 (
            .O(N__47316),
            .I(N__47313));
    InMux I__10898 (
            .O(N__47313),
            .I(N__47310));
    LocalMux I__10897 (
            .O(N__47310),
            .I(n21368));
    InMux I__10896 (
            .O(N__47307),
            .I(N__47304));
    LocalMux I__10895 (
            .O(N__47304),
            .I(n21369));
    InMux I__10894 (
            .O(N__47301),
            .I(N__47298));
    LocalMux I__10893 (
            .O(N__47298),
            .I(N__47295));
    Odrv4 I__10892 (
            .O(N__47295),
            .I(n21362));
    InMux I__10891 (
            .O(N__47292),
            .I(N__47289));
    LocalMux I__10890 (
            .O(N__47289),
            .I(N__47286));
    Span4Mux_h I__10889 (
            .O(N__47286),
            .I(N__47283));
    Span4Mux_h I__10888 (
            .O(N__47283),
            .I(N__47280));
    Span4Mux_h I__10887 (
            .O(N__47280),
            .I(N__47277));
    Odrv4 I__10886 (
            .O(N__47277),
            .I(n21363));
    CascadeMux I__10885 (
            .O(N__47274),
            .I(n22599_cascade_));
    InMux I__10884 (
            .O(N__47271),
            .I(N__47264));
    InMux I__10883 (
            .O(N__47270),
            .I(N__47259));
    InMux I__10882 (
            .O(N__47269),
            .I(N__47246));
    InMux I__10881 (
            .O(N__47268),
            .I(N__47240));
    InMux I__10880 (
            .O(N__47267),
            .I(N__47237));
    LocalMux I__10879 (
            .O(N__47264),
            .I(N__47234));
    InMux I__10878 (
            .O(N__47263),
            .I(N__47227));
    InMux I__10877 (
            .O(N__47262),
            .I(N__47227));
    LocalMux I__10876 (
            .O(N__47259),
            .I(N__47224));
    InMux I__10875 (
            .O(N__47258),
            .I(N__47221));
    InMux I__10874 (
            .O(N__47257),
            .I(N__47218));
    InMux I__10873 (
            .O(N__47256),
            .I(N__47215));
    InMux I__10872 (
            .O(N__47255),
            .I(N__47212));
    InMux I__10871 (
            .O(N__47254),
            .I(N__47209));
    InMux I__10870 (
            .O(N__47253),
            .I(N__47204));
    InMux I__10869 (
            .O(N__47252),
            .I(N__47204));
    InMux I__10868 (
            .O(N__47251),
            .I(N__47197));
    InMux I__10867 (
            .O(N__47250),
            .I(N__47197));
    InMux I__10866 (
            .O(N__47249),
            .I(N__47197));
    LocalMux I__10865 (
            .O(N__47246),
            .I(N__47187));
    InMux I__10864 (
            .O(N__47245),
            .I(N__47182));
    InMux I__10863 (
            .O(N__47244),
            .I(N__47182));
    InMux I__10862 (
            .O(N__47243),
            .I(N__47179));
    LocalMux I__10861 (
            .O(N__47240),
            .I(N__47176));
    LocalMux I__10860 (
            .O(N__47237),
            .I(N__47171));
    Span4Mux_v I__10859 (
            .O(N__47234),
            .I(N__47171));
    InMux I__10858 (
            .O(N__47233),
            .I(N__47166));
    InMux I__10857 (
            .O(N__47232),
            .I(N__47166));
    LocalMux I__10856 (
            .O(N__47227),
            .I(N__47160));
    Span4Mux_v I__10855 (
            .O(N__47224),
            .I(N__47155));
    LocalMux I__10854 (
            .O(N__47221),
            .I(N__47150));
    LocalMux I__10853 (
            .O(N__47218),
            .I(N__47137));
    LocalMux I__10852 (
            .O(N__47215),
            .I(N__47137));
    LocalMux I__10851 (
            .O(N__47212),
            .I(N__47137));
    LocalMux I__10850 (
            .O(N__47209),
            .I(N__47137));
    LocalMux I__10849 (
            .O(N__47204),
            .I(N__47137));
    LocalMux I__10848 (
            .O(N__47197),
            .I(N__47137));
    InMux I__10847 (
            .O(N__47196),
            .I(N__47128));
    InMux I__10846 (
            .O(N__47195),
            .I(N__47123));
    InMux I__10845 (
            .O(N__47194),
            .I(N__47123));
    InMux I__10844 (
            .O(N__47193),
            .I(N__47120));
    InMux I__10843 (
            .O(N__47192),
            .I(N__47117));
    InMux I__10842 (
            .O(N__47191),
            .I(N__47112));
    InMux I__10841 (
            .O(N__47190),
            .I(N__47112));
    Span4Mux_h I__10840 (
            .O(N__47187),
            .I(N__47107));
    LocalMux I__10839 (
            .O(N__47182),
            .I(N__47107));
    LocalMux I__10838 (
            .O(N__47179),
            .I(N__47098));
    Span4Mux_h I__10837 (
            .O(N__47176),
            .I(N__47098));
    Span4Mux_v I__10836 (
            .O(N__47171),
            .I(N__47098));
    LocalMux I__10835 (
            .O(N__47166),
            .I(N__47098));
    InMux I__10834 (
            .O(N__47165),
            .I(N__47095));
    InMux I__10833 (
            .O(N__47164),
            .I(N__47092));
    InMux I__10832 (
            .O(N__47163),
            .I(N__47088));
    Sp12to4 I__10831 (
            .O(N__47160),
            .I(N__47085));
    InMux I__10830 (
            .O(N__47159),
            .I(N__47080));
    InMux I__10829 (
            .O(N__47158),
            .I(N__47080));
    Span4Mux_v I__10828 (
            .O(N__47155),
            .I(N__47077));
    InMux I__10827 (
            .O(N__47154),
            .I(N__47072));
    InMux I__10826 (
            .O(N__47153),
            .I(N__47072));
    Span4Mux_v I__10825 (
            .O(N__47150),
            .I(N__47067));
    Span4Mux_v I__10824 (
            .O(N__47137),
            .I(N__47067));
    InMux I__10823 (
            .O(N__47136),
            .I(N__47058));
    InMux I__10822 (
            .O(N__47135),
            .I(N__47058));
    InMux I__10821 (
            .O(N__47134),
            .I(N__47058));
    InMux I__10820 (
            .O(N__47133),
            .I(N__47058));
    InMux I__10819 (
            .O(N__47132),
            .I(N__47055));
    CascadeMux I__10818 (
            .O(N__47131),
            .I(N__47052));
    LocalMux I__10817 (
            .O(N__47128),
            .I(N__47049));
    LocalMux I__10816 (
            .O(N__47123),
            .I(N__47041));
    LocalMux I__10815 (
            .O(N__47120),
            .I(N__47041));
    LocalMux I__10814 (
            .O(N__47117),
            .I(N__47041));
    LocalMux I__10813 (
            .O(N__47112),
            .I(N__47034));
    Span4Mux_v I__10812 (
            .O(N__47107),
            .I(N__47034));
    Span4Mux_h I__10811 (
            .O(N__47098),
            .I(N__47034));
    LocalMux I__10810 (
            .O(N__47095),
            .I(N__47029));
    LocalMux I__10809 (
            .O(N__47092),
            .I(N__47029));
    InMux I__10808 (
            .O(N__47091),
            .I(N__47026));
    LocalMux I__10807 (
            .O(N__47088),
            .I(N__47009));
    Span12Mux_v I__10806 (
            .O(N__47085),
            .I(N__47009));
    LocalMux I__10805 (
            .O(N__47080),
            .I(N__47009));
    Sp12to4 I__10804 (
            .O(N__47077),
            .I(N__47009));
    LocalMux I__10803 (
            .O(N__47072),
            .I(N__47009));
    Sp12to4 I__10802 (
            .O(N__47067),
            .I(N__47009));
    LocalMux I__10801 (
            .O(N__47058),
            .I(N__47009));
    LocalMux I__10800 (
            .O(N__47055),
            .I(N__47009));
    InMux I__10799 (
            .O(N__47052),
            .I(N__47006));
    Span12Mux_h I__10798 (
            .O(N__47049),
            .I(N__47003));
    InMux I__10797 (
            .O(N__47048),
            .I(N__47000));
    Span12Mux_h I__10796 (
            .O(N__47041),
            .I(N__46997));
    Span4Mux_h I__10795 (
            .O(N__47034),
            .I(N__46994));
    Span4Mux_h I__10794 (
            .O(N__47029),
            .I(N__46991));
    LocalMux I__10793 (
            .O(N__47026),
            .I(N__46986));
    Span12Mux_h I__10792 (
            .O(N__47009),
            .I(N__46986));
    LocalMux I__10791 (
            .O(N__47006),
            .I(comm_cmd_3));
    Odrv12 I__10790 (
            .O(N__47003),
            .I(comm_cmd_3));
    LocalMux I__10789 (
            .O(N__47000),
            .I(comm_cmd_3));
    Odrv12 I__10788 (
            .O(N__46997),
            .I(comm_cmd_3));
    Odrv4 I__10787 (
            .O(N__46994),
            .I(comm_cmd_3));
    Odrv4 I__10786 (
            .O(N__46991),
            .I(comm_cmd_3));
    Odrv12 I__10785 (
            .O(N__46986),
            .I(comm_cmd_3));
    InMux I__10784 (
            .O(N__46971),
            .I(N__46968));
    LocalMux I__10783 (
            .O(N__46968),
            .I(n22602));
    InMux I__10782 (
            .O(N__46965),
            .I(N__46962));
    LocalMux I__10781 (
            .O(N__46962),
            .I(N__46959));
    Span4Mux_v I__10780 (
            .O(N__46959),
            .I(N__46954));
    InMux I__10779 (
            .O(N__46958),
            .I(N__46951));
    InMux I__10778 (
            .O(N__46957),
            .I(N__46948));
    Sp12to4 I__10777 (
            .O(N__46954),
            .I(N__46943));
    LocalMux I__10776 (
            .O(N__46951),
            .I(N__46943));
    LocalMux I__10775 (
            .O(N__46948),
            .I(buf_dds1_6));
    Odrv12 I__10774 (
            .O(N__46943),
            .I(buf_dds1_6));
    InMux I__10773 (
            .O(N__46938),
            .I(N__46935));
    LocalMux I__10772 (
            .O(N__46935),
            .I(N__46931));
    CascadeMux I__10771 (
            .O(N__46934),
            .I(N__46928));
    Span4Mux_h I__10770 (
            .O(N__46931),
            .I(N__46925));
    InMux I__10769 (
            .O(N__46928),
            .I(N__46922));
    Odrv4 I__10768 (
            .O(N__46925),
            .I(n68));
    LocalMux I__10767 (
            .O(N__46922),
            .I(n68));
    CascadeMux I__10766 (
            .O(N__46917),
            .I(N__46911));
    InMux I__10765 (
            .O(N__46916),
            .I(N__46906));
    InMux I__10764 (
            .O(N__46915),
            .I(N__46903));
    InMux I__10763 (
            .O(N__46914),
            .I(N__46900));
    InMux I__10762 (
            .O(N__46911),
            .I(N__46895));
    CascadeMux I__10761 (
            .O(N__46910),
            .I(N__46891));
    InMux I__10760 (
            .O(N__46909),
            .I(N__46886));
    LocalMux I__10759 (
            .O(N__46906),
            .I(N__46878));
    LocalMux I__10758 (
            .O(N__46903),
            .I(N__46878));
    LocalMux I__10757 (
            .O(N__46900),
            .I(N__46878));
    CascadeMux I__10756 (
            .O(N__46899),
            .I(N__46875));
    InMux I__10755 (
            .O(N__46898),
            .I(N__46869));
    LocalMux I__10754 (
            .O(N__46895),
            .I(N__46866));
    InMux I__10753 (
            .O(N__46894),
            .I(N__46859));
    InMux I__10752 (
            .O(N__46891),
            .I(N__46859));
    InMux I__10751 (
            .O(N__46890),
            .I(N__46859));
    InMux I__10750 (
            .O(N__46889),
            .I(N__46856));
    LocalMux I__10749 (
            .O(N__46886),
            .I(N__46853));
    InMux I__10748 (
            .O(N__46885),
            .I(N__46850));
    Span4Mux_v I__10747 (
            .O(N__46878),
            .I(N__46847));
    InMux I__10746 (
            .O(N__46875),
            .I(N__46842));
    InMux I__10745 (
            .O(N__46874),
            .I(N__46842));
    InMux I__10744 (
            .O(N__46873),
            .I(N__46839));
    InMux I__10743 (
            .O(N__46872),
            .I(N__46836));
    LocalMux I__10742 (
            .O(N__46869),
            .I(N__46833));
    Span4Mux_h I__10741 (
            .O(N__46866),
            .I(N__46828));
    LocalMux I__10740 (
            .O(N__46859),
            .I(N__46828));
    LocalMux I__10739 (
            .O(N__46856),
            .I(N__46823));
    Span4Mux_h I__10738 (
            .O(N__46853),
            .I(N__46823));
    LocalMux I__10737 (
            .O(N__46850),
            .I(N__46818));
    Span4Mux_h I__10736 (
            .O(N__46847),
            .I(N__46818));
    LocalMux I__10735 (
            .O(N__46842),
            .I(N__46811));
    LocalMux I__10734 (
            .O(N__46839),
            .I(N__46811));
    LocalMux I__10733 (
            .O(N__46836),
            .I(N__46811));
    Span4Mux_h I__10732 (
            .O(N__46833),
            .I(N__46807));
    Span4Mux_v I__10731 (
            .O(N__46828),
            .I(N__46804));
    Span4Mux_h I__10730 (
            .O(N__46823),
            .I(N__46801));
    Span4Mux_h I__10729 (
            .O(N__46818),
            .I(N__46796));
    Span4Mux_v I__10728 (
            .O(N__46811),
            .I(N__46796));
    InMux I__10727 (
            .O(N__46810),
            .I(N__46793));
    Span4Mux_v I__10726 (
            .O(N__46807),
            .I(N__46790));
    Span4Mux_h I__10725 (
            .O(N__46804),
            .I(N__46787));
    Span4Mux_h I__10724 (
            .O(N__46801),
            .I(N__46784));
    Span4Mux_h I__10723 (
            .O(N__46796),
            .I(N__46781));
    LocalMux I__10722 (
            .O(N__46793),
            .I(n12048));
    Odrv4 I__10721 (
            .O(N__46790),
            .I(n12048));
    Odrv4 I__10720 (
            .O(N__46787),
            .I(n12048));
    Odrv4 I__10719 (
            .O(N__46784),
            .I(n12048));
    Odrv4 I__10718 (
            .O(N__46781),
            .I(n12048));
    CascadeMux I__10717 (
            .O(N__46770),
            .I(n12048_cascade_));
    CascadeMux I__10716 (
            .O(N__46767),
            .I(N__46760));
    InMux I__10715 (
            .O(N__46766),
            .I(N__46757));
    InMux I__10714 (
            .O(N__46765),
            .I(N__46747));
    InMux I__10713 (
            .O(N__46764),
            .I(N__46747));
    InMux I__10712 (
            .O(N__46763),
            .I(N__46747));
    InMux I__10711 (
            .O(N__46760),
            .I(N__46742));
    LocalMux I__10710 (
            .O(N__46757),
            .I(N__46739));
    InMux I__10709 (
            .O(N__46756),
            .I(N__46734));
    InMux I__10708 (
            .O(N__46755),
            .I(N__46734));
    InMux I__10707 (
            .O(N__46754),
            .I(N__46729));
    LocalMux I__10706 (
            .O(N__46747),
            .I(N__46726));
    InMux I__10705 (
            .O(N__46746),
            .I(N__46723));
    InMux I__10704 (
            .O(N__46745),
            .I(N__46720));
    LocalMux I__10703 (
            .O(N__46742),
            .I(N__46717));
    Span4Mux_v I__10702 (
            .O(N__46739),
            .I(N__46712));
    LocalMux I__10701 (
            .O(N__46734),
            .I(N__46712));
    InMux I__10700 (
            .O(N__46733),
            .I(N__46709));
    InMux I__10699 (
            .O(N__46732),
            .I(N__46706));
    LocalMux I__10698 (
            .O(N__46729),
            .I(N__46703));
    Span4Mux_v I__10697 (
            .O(N__46726),
            .I(N__46700));
    LocalMux I__10696 (
            .O(N__46723),
            .I(N__46697));
    LocalMux I__10695 (
            .O(N__46720),
            .I(N__46689));
    Span4Mux_v I__10694 (
            .O(N__46717),
            .I(N__46689));
    Span4Mux_h I__10693 (
            .O(N__46712),
            .I(N__46689));
    LocalMux I__10692 (
            .O(N__46709),
            .I(N__46686));
    LocalMux I__10691 (
            .O(N__46706),
            .I(N__46681));
    Span4Mux_v I__10690 (
            .O(N__46703),
            .I(N__46681));
    Span4Mux_h I__10689 (
            .O(N__46700),
            .I(N__46676));
    Span4Mux_h I__10688 (
            .O(N__46697),
            .I(N__46676));
    InMux I__10687 (
            .O(N__46696),
            .I(N__46673));
    Span4Mux_h I__10686 (
            .O(N__46689),
            .I(N__46670));
    Span12Mux_v I__10685 (
            .O(N__46686),
            .I(N__46665));
    Sp12to4 I__10684 (
            .O(N__46681),
            .I(N__46665));
    Span4Mux_v I__10683 (
            .O(N__46676),
            .I(N__46662));
    LocalMux I__10682 (
            .O(N__46673),
            .I(n16971));
    Odrv4 I__10681 (
            .O(N__46670),
            .I(n16971));
    Odrv12 I__10680 (
            .O(N__46665),
            .I(n16971));
    Odrv4 I__10679 (
            .O(N__46662),
            .I(n16971));
    InMux I__10678 (
            .O(N__46653),
            .I(N__46650));
    LocalMux I__10677 (
            .O(N__46650),
            .I(\comm_spi.n14805 ));
    SRMux I__10676 (
            .O(N__46647),
            .I(N__46644));
    LocalMux I__10675 (
            .O(N__46644),
            .I(\comm_spi.iclk_N_802 ));
    CascadeMux I__10674 (
            .O(N__46641),
            .I(N__46637));
    CascadeMux I__10673 (
            .O(N__46640),
            .I(N__46634));
    InMux I__10672 (
            .O(N__46637),
            .I(N__46631));
    InMux I__10671 (
            .O(N__46634),
            .I(N__46628));
    LocalMux I__10670 (
            .O(N__46631),
            .I(N__46625));
    LocalMux I__10669 (
            .O(N__46628),
            .I(comm_buf_6_0));
    Odrv4 I__10668 (
            .O(N__46625),
            .I(comm_buf_6_0));
    InMux I__10667 (
            .O(N__46620),
            .I(N__46617));
    LocalMux I__10666 (
            .O(N__46617),
            .I(N__46613));
    InMux I__10665 (
            .O(N__46616),
            .I(N__46610));
    Span4Mux_v I__10664 (
            .O(N__46613),
            .I(N__46607));
    LocalMux I__10663 (
            .O(N__46610),
            .I(comm_buf_6_3));
    Odrv4 I__10662 (
            .O(N__46607),
            .I(comm_buf_6_3));
    InMux I__10661 (
            .O(N__46602),
            .I(N__46599));
    LocalMux I__10660 (
            .O(N__46599),
            .I(N__46595));
    InMux I__10659 (
            .O(N__46598),
            .I(N__46591));
    Span4Mux_h I__10658 (
            .O(N__46595),
            .I(N__46588));
    InMux I__10657 (
            .O(N__46594),
            .I(N__46585));
    LocalMux I__10656 (
            .O(N__46591),
            .I(acadc_skipCount_7));
    Odrv4 I__10655 (
            .O(N__46588),
            .I(acadc_skipCount_7));
    LocalMux I__10654 (
            .O(N__46585),
            .I(acadc_skipCount_7));
    InMux I__10653 (
            .O(N__46578),
            .I(N__46575));
    LocalMux I__10652 (
            .O(N__46575),
            .I(N__46572));
    Span4Mux_v I__10651 (
            .O(N__46572),
            .I(N__46568));
    InMux I__10650 (
            .O(N__46571),
            .I(N__46564));
    Span4Mux_h I__10649 (
            .O(N__46568),
            .I(N__46561));
    InMux I__10648 (
            .O(N__46567),
            .I(N__46558));
    LocalMux I__10647 (
            .O(N__46564),
            .I(req_data_cnt_7));
    Odrv4 I__10646 (
            .O(N__46561),
            .I(req_data_cnt_7));
    LocalMux I__10645 (
            .O(N__46558),
            .I(req_data_cnt_7));
    InMux I__10644 (
            .O(N__46551),
            .I(N__46548));
    LocalMux I__10643 (
            .O(N__46548),
            .I(N__46545));
    Span4Mux_h I__10642 (
            .O(N__46545),
            .I(N__46541));
    InMux I__10641 (
            .O(N__46544),
            .I(N__46538));
    Span4Mux_h I__10640 (
            .O(N__46541),
            .I(N__46535));
    LocalMux I__10639 (
            .O(N__46538),
            .I(N__46530));
    Span4Mux_v I__10638 (
            .O(N__46535),
            .I(N__46530));
    Odrv4 I__10637 (
            .O(N__46530),
            .I(data_idxvec_7));
    InMux I__10636 (
            .O(N__46527),
            .I(N__46523));
    InMux I__10635 (
            .O(N__46526),
            .I(N__46520));
    LocalMux I__10634 (
            .O(N__46523),
            .I(N__46516));
    LocalMux I__10633 (
            .O(N__46520),
            .I(N__46513));
    InMux I__10632 (
            .O(N__46519),
            .I(N__46510));
    Span4Mux_v I__10631 (
            .O(N__46516),
            .I(N__46505));
    Span4Mux_h I__10630 (
            .O(N__46513),
            .I(N__46505));
    LocalMux I__10629 (
            .O(N__46510),
            .I(data_cntvec_7));
    Odrv4 I__10628 (
            .O(N__46505),
            .I(data_cntvec_7));
    InMux I__10627 (
            .O(N__46500),
            .I(N__46497));
    LocalMux I__10626 (
            .O(N__46497),
            .I(N__46494));
    Span4Mux_v I__10625 (
            .O(N__46494),
            .I(N__46491));
    Odrv4 I__10624 (
            .O(N__46491),
            .I(buf_data_iac_15));
    CascadeMux I__10623 (
            .O(N__46488),
            .I(n26_adj_1622_cascade_));
    InMux I__10622 (
            .O(N__46485),
            .I(N__46450));
    InMux I__10621 (
            .O(N__46484),
            .I(N__46445));
    InMux I__10620 (
            .O(N__46483),
            .I(N__46445));
    InMux I__10619 (
            .O(N__46482),
            .I(N__46438));
    InMux I__10618 (
            .O(N__46481),
            .I(N__46438));
    InMux I__10617 (
            .O(N__46480),
            .I(N__46438));
    InMux I__10616 (
            .O(N__46479),
            .I(N__46433));
    InMux I__10615 (
            .O(N__46478),
            .I(N__46433));
    InMux I__10614 (
            .O(N__46477),
            .I(N__46430));
    InMux I__10613 (
            .O(N__46476),
            .I(N__46425));
    InMux I__10612 (
            .O(N__46475),
            .I(N__46425));
    InMux I__10611 (
            .O(N__46474),
            .I(N__46418));
    InMux I__10610 (
            .O(N__46473),
            .I(N__46418));
    InMux I__10609 (
            .O(N__46472),
            .I(N__46418));
    InMux I__10608 (
            .O(N__46471),
            .I(N__46415));
    InMux I__10607 (
            .O(N__46470),
            .I(N__46412));
    CascadeMux I__10606 (
            .O(N__46469),
            .I(N__46403));
    InMux I__10605 (
            .O(N__46468),
            .I(N__46397));
    InMux I__10604 (
            .O(N__46467),
            .I(N__46397));
    InMux I__10603 (
            .O(N__46466),
            .I(N__46392));
    InMux I__10602 (
            .O(N__46465),
            .I(N__46392));
    InMux I__10601 (
            .O(N__46464),
            .I(N__46387));
    InMux I__10600 (
            .O(N__46463),
            .I(N__46387));
    InMux I__10599 (
            .O(N__46462),
            .I(N__46384));
    InMux I__10598 (
            .O(N__46461),
            .I(N__46381));
    InMux I__10597 (
            .O(N__46460),
            .I(N__46378));
    InMux I__10596 (
            .O(N__46459),
            .I(N__46360));
    InMux I__10595 (
            .O(N__46458),
            .I(N__46360));
    InMux I__10594 (
            .O(N__46457),
            .I(N__46360));
    InMux I__10593 (
            .O(N__46456),
            .I(N__46360));
    InMux I__10592 (
            .O(N__46455),
            .I(N__46357));
    InMux I__10591 (
            .O(N__46454),
            .I(N__46354));
    InMux I__10590 (
            .O(N__46453),
            .I(N__46351));
    LocalMux I__10589 (
            .O(N__46450),
            .I(N__46346));
    LocalMux I__10588 (
            .O(N__46445),
            .I(N__46346));
    LocalMux I__10587 (
            .O(N__46438),
            .I(N__46339));
    LocalMux I__10586 (
            .O(N__46433),
            .I(N__46339));
    LocalMux I__10585 (
            .O(N__46430),
            .I(N__46339));
    LocalMux I__10584 (
            .O(N__46425),
            .I(N__46336));
    LocalMux I__10583 (
            .O(N__46418),
            .I(N__46329));
    LocalMux I__10582 (
            .O(N__46415),
            .I(N__46329));
    LocalMux I__10581 (
            .O(N__46412),
            .I(N__46329));
    InMux I__10580 (
            .O(N__46411),
            .I(N__46324));
    InMux I__10579 (
            .O(N__46410),
            .I(N__46324));
    InMux I__10578 (
            .O(N__46409),
            .I(N__46319));
    InMux I__10577 (
            .O(N__46408),
            .I(N__46319));
    InMux I__10576 (
            .O(N__46407),
            .I(N__46312));
    InMux I__10575 (
            .O(N__46406),
            .I(N__46312));
    InMux I__10574 (
            .O(N__46403),
            .I(N__46303));
    InMux I__10573 (
            .O(N__46402),
            .I(N__46292));
    LocalMux I__10572 (
            .O(N__46397),
            .I(N__46287));
    LocalMux I__10571 (
            .O(N__46392),
            .I(N__46278));
    LocalMux I__10570 (
            .O(N__46387),
            .I(N__46278));
    LocalMux I__10569 (
            .O(N__46384),
            .I(N__46278));
    LocalMux I__10568 (
            .O(N__46381),
            .I(N__46278));
    LocalMux I__10567 (
            .O(N__46378),
            .I(N__46275));
    InMux I__10566 (
            .O(N__46377),
            .I(N__46272));
    InMux I__10565 (
            .O(N__46376),
            .I(N__46269));
    InMux I__10564 (
            .O(N__46375),
            .I(N__46262));
    InMux I__10563 (
            .O(N__46374),
            .I(N__46262));
    InMux I__10562 (
            .O(N__46373),
            .I(N__46262));
    InMux I__10561 (
            .O(N__46372),
            .I(N__46259));
    InMux I__10560 (
            .O(N__46371),
            .I(N__46249));
    InMux I__10559 (
            .O(N__46370),
            .I(N__46249));
    InMux I__10558 (
            .O(N__46369),
            .I(N__46249));
    LocalMux I__10557 (
            .O(N__46360),
            .I(N__46244));
    LocalMux I__10556 (
            .O(N__46357),
            .I(N__46244));
    LocalMux I__10555 (
            .O(N__46354),
            .I(N__46241));
    LocalMux I__10554 (
            .O(N__46351),
            .I(N__46238));
    Span4Mux_v I__10553 (
            .O(N__46346),
            .I(N__46225));
    Span4Mux_v I__10552 (
            .O(N__46339),
            .I(N__46225));
    Span4Mux_v I__10551 (
            .O(N__46336),
            .I(N__46225));
    Span4Mux_v I__10550 (
            .O(N__46329),
            .I(N__46225));
    LocalMux I__10549 (
            .O(N__46324),
            .I(N__46225));
    LocalMux I__10548 (
            .O(N__46319),
            .I(N__46225));
    InMux I__10547 (
            .O(N__46318),
            .I(N__46221));
    InMux I__10546 (
            .O(N__46317),
            .I(N__46218));
    LocalMux I__10545 (
            .O(N__46312),
            .I(N__46215));
    InMux I__10544 (
            .O(N__46311),
            .I(N__46210));
    InMux I__10543 (
            .O(N__46310),
            .I(N__46210));
    InMux I__10542 (
            .O(N__46309),
            .I(N__46203));
    InMux I__10541 (
            .O(N__46308),
            .I(N__46203));
    InMux I__10540 (
            .O(N__46307),
            .I(N__46203));
    InMux I__10539 (
            .O(N__46306),
            .I(N__46200));
    LocalMux I__10538 (
            .O(N__46303),
            .I(N__46197));
    InMux I__10537 (
            .O(N__46302),
            .I(N__46186));
    InMux I__10536 (
            .O(N__46301),
            .I(N__46186));
    InMux I__10535 (
            .O(N__46300),
            .I(N__46186));
    InMux I__10534 (
            .O(N__46299),
            .I(N__46186));
    InMux I__10533 (
            .O(N__46298),
            .I(N__46186));
    InMux I__10532 (
            .O(N__46297),
            .I(N__46183));
    InMux I__10531 (
            .O(N__46296),
            .I(N__46178));
    InMux I__10530 (
            .O(N__46295),
            .I(N__46178));
    LocalMux I__10529 (
            .O(N__46292),
            .I(N__46175));
    InMux I__10528 (
            .O(N__46291),
            .I(N__46172));
    InMux I__10527 (
            .O(N__46290),
            .I(N__46169));
    Span4Mux_v I__10526 (
            .O(N__46287),
            .I(N__46160));
    Span4Mux_v I__10525 (
            .O(N__46278),
            .I(N__46160));
    Span4Mux_h I__10524 (
            .O(N__46275),
            .I(N__46160));
    LocalMux I__10523 (
            .O(N__46272),
            .I(N__46160));
    LocalMux I__10522 (
            .O(N__46269),
            .I(N__46152));
    LocalMux I__10521 (
            .O(N__46262),
            .I(N__46152));
    LocalMux I__10520 (
            .O(N__46259),
            .I(N__46152));
    InMux I__10519 (
            .O(N__46258),
            .I(N__46149));
    InMux I__10518 (
            .O(N__46257),
            .I(N__46146));
    InMux I__10517 (
            .O(N__46256),
            .I(N__46143));
    LocalMux I__10516 (
            .O(N__46249),
            .I(N__46132));
    Span4Mux_v I__10515 (
            .O(N__46244),
            .I(N__46132));
    Span4Mux_v I__10514 (
            .O(N__46241),
            .I(N__46132));
    Span4Mux_v I__10513 (
            .O(N__46238),
            .I(N__46132));
    Span4Mux_h I__10512 (
            .O(N__46225),
            .I(N__46132));
    InMux I__10511 (
            .O(N__46224),
            .I(N__46129));
    LocalMux I__10510 (
            .O(N__46221),
            .I(N__46122));
    LocalMux I__10509 (
            .O(N__46218),
            .I(N__46122));
    Span4Mux_v I__10508 (
            .O(N__46215),
            .I(N__46122));
    LocalMux I__10507 (
            .O(N__46210),
            .I(N__46111));
    LocalMux I__10506 (
            .O(N__46203),
            .I(N__46111));
    LocalMux I__10505 (
            .O(N__46200),
            .I(N__46111));
    Span4Mux_v I__10504 (
            .O(N__46197),
            .I(N__46111));
    LocalMux I__10503 (
            .O(N__46186),
            .I(N__46111));
    LocalMux I__10502 (
            .O(N__46183),
            .I(N__46098));
    LocalMux I__10501 (
            .O(N__46178),
            .I(N__46098));
    Span4Mux_v I__10500 (
            .O(N__46175),
            .I(N__46098));
    LocalMux I__10499 (
            .O(N__46172),
            .I(N__46098));
    LocalMux I__10498 (
            .O(N__46169),
            .I(N__46098));
    Span4Mux_v I__10497 (
            .O(N__46160),
            .I(N__46098));
    InMux I__10496 (
            .O(N__46159),
            .I(N__46095));
    Span12Mux_h I__10495 (
            .O(N__46152),
            .I(N__46092));
    LocalMux I__10494 (
            .O(N__46149),
            .I(N__46089));
    LocalMux I__10493 (
            .O(N__46146),
            .I(N__46084));
    LocalMux I__10492 (
            .O(N__46143),
            .I(N__46084));
    Span4Mux_h I__10491 (
            .O(N__46132),
            .I(N__46081));
    LocalMux I__10490 (
            .O(N__46129),
            .I(N__46072));
    Span4Mux_v I__10489 (
            .O(N__46122),
            .I(N__46072));
    Span4Mux_v I__10488 (
            .O(N__46111),
            .I(N__46072));
    Span4Mux_h I__10487 (
            .O(N__46098),
            .I(N__46072));
    LocalMux I__10486 (
            .O(N__46095),
            .I(comm_cmd_1));
    Odrv12 I__10485 (
            .O(N__46092),
            .I(comm_cmd_1));
    Odrv4 I__10484 (
            .O(N__46089),
            .I(comm_cmd_1));
    Odrv4 I__10483 (
            .O(N__46084),
            .I(comm_cmd_1));
    Odrv4 I__10482 (
            .O(N__46081),
            .I(comm_cmd_1));
    Odrv4 I__10481 (
            .O(N__46072),
            .I(comm_cmd_1));
    SRMux I__10480 (
            .O(N__46059),
            .I(N__46056));
    LocalMux I__10479 (
            .O(N__46056),
            .I(N__46053));
    Span4Mux_v I__10478 (
            .O(N__46053),
            .I(N__46050));
    Odrv4 I__10477 (
            .O(N__46050),
            .I(n16824));
    InMux I__10476 (
            .O(N__46047),
            .I(N__46044));
    LocalMux I__10475 (
            .O(N__46044),
            .I(N__46041));
    Odrv4 I__10474 (
            .O(N__46041),
            .I(comm_length_1));
    InMux I__10473 (
            .O(N__46038),
            .I(N__46033));
    InMux I__10472 (
            .O(N__46037),
            .I(N__46030));
    InMux I__10471 (
            .O(N__46036),
            .I(N__46027));
    LocalMux I__10470 (
            .O(N__46033),
            .I(N__46024));
    LocalMux I__10469 (
            .O(N__46030),
            .I(N__46021));
    LocalMux I__10468 (
            .O(N__46027),
            .I(N__46018));
    Span4Mux_h I__10467 (
            .O(N__46024),
            .I(N__46015));
    Span12Mux_v I__10466 (
            .O(N__46021),
            .I(N__46010));
    Span12Mux_h I__10465 (
            .O(N__46018),
            .I(N__46010));
    Odrv4 I__10464 (
            .O(N__46015),
            .I(n5_adj_1524));
    Odrv12 I__10463 (
            .O(N__46010),
            .I(n5_adj_1524));
    InMux I__10462 (
            .O(N__46005),
            .I(N__46002));
    LocalMux I__10461 (
            .O(N__46002),
            .I(N__45999));
    Span4Mux_h I__10460 (
            .O(N__45999),
            .I(N__45996));
    Span4Mux_h I__10459 (
            .O(N__45996),
            .I(N__45993));
    Odrv4 I__10458 (
            .O(N__45993),
            .I(n30_adj_1605));
    InMux I__10457 (
            .O(N__45990),
            .I(N__45987));
    LocalMux I__10456 (
            .O(N__45987),
            .I(N__45984));
    Span4Mux_v I__10455 (
            .O(N__45984),
            .I(N__45981));
    Sp12to4 I__10454 (
            .O(N__45981),
            .I(N__45978));
    Odrv12 I__10453 (
            .O(N__45978),
            .I(n30_adj_1608));
    CascadeMux I__10452 (
            .O(N__45975),
            .I(N__45972));
    InMux I__10451 (
            .O(N__45972),
            .I(N__45969));
    LocalMux I__10450 (
            .O(N__45969),
            .I(N__45966));
    Odrv4 I__10449 (
            .O(N__45966),
            .I(comm_buf_2_4));
    InMux I__10448 (
            .O(N__45963),
            .I(N__45960));
    LocalMux I__10447 (
            .O(N__45960),
            .I(N__45957));
    Span4Mux_v I__10446 (
            .O(N__45957),
            .I(N__45954));
    Span4Mux_h I__10445 (
            .O(N__45954),
            .I(N__45951));
    Odrv4 I__10444 (
            .O(N__45951),
            .I(n30_adj_1611));
    InMux I__10443 (
            .O(N__45948),
            .I(N__45945));
    LocalMux I__10442 (
            .O(N__45945),
            .I(N__45942));
    Odrv4 I__10441 (
            .O(N__45942),
            .I(comm_buf_2_3));
    InMux I__10440 (
            .O(N__45939),
            .I(N__45936));
    LocalMux I__10439 (
            .O(N__45936),
            .I(N__45933));
    Span12Mux_v I__10438 (
            .O(N__45933),
            .I(N__45930));
    Odrv12 I__10437 (
            .O(N__45930),
            .I(n30_adj_1614));
    InMux I__10436 (
            .O(N__45927),
            .I(N__45924));
    LocalMux I__10435 (
            .O(N__45924),
            .I(N__45921));
    Odrv12 I__10434 (
            .O(N__45921),
            .I(comm_buf_2_2));
    InMux I__10433 (
            .O(N__45918),
            .I(N__45915));
    LocalMux I__10432 (
            .O(N__45915),
            .I(N__45912));
    Span4Mux_h I__10431 (
            .O(N__45912),
            .I(N__45909));
    Odrv4 I__10430 (
            .O(N__45909),
            .I(n30_adj_1618));
    CEMux I__10429 (
            .O(N__45906),
            .I(N__45903));
    LocalMux I__10428 (
            .O(N__45903),
            .I(N__45899));
    InMux I__10427 (
            .O(N__45902),
            .I(N__45896));
    Odrv4 I__10426 (
            .O(N__45899),
            .I(n12314));
    LocalMux I__10425 (
            .O(N__45896),
            .I(n12314));
    SRMux I__10424 (
            .O(N__45891),
            .I(N__45888));
    LocalMux I__10423 (
            .O(N__45888),
            .I(N__45885));
    Span4Mux_h I__10422 (
            .O(N__45885),
            .I(N__45882));
    Odrv4 I__10421 (
            .O(N__45882),
            .I(n14972));
    CascadeMux I__10420 (
            .O(N__45879),
            .I(N__45875));
    CascadeMux I__10419 (
            .O(N__45878),
            .I(N__45871));
    InMux I__10418 (
            .O(N__45875),
            .I(N__45865));
    CascadeMux I__10417 (
            .O(N__45874),
            .I(N__45861));
    InMux I__10416 (
            .O(N__45871),
            .I(N__45858));
    InMux I__10415 (
            .O(N__45870),
            .I(N__45855));
    CascadeMux I__10414 (
            .O(N__45869),
            .I(N__45852));
    CascadeMux I__10413 (
            .O(N__45868),
            .I(N__45849));
    LocalMux I__10412 (
            .O(N__45865),
            .I(N__45845));
    CascadeMux I__10411 (
            .O(N__45864),
            .I(N__45842));
    InMux I__10410 (
            .O(N__45861),
            .I(N__45839));
    LocalMux I__10409 (
            .O(N__45858),
            .I(N__45836));
    LocalMux I__10408 (
            .O(N__45855),
            .I(N__45833));
    InMux I__10407 (
            .O(N__45852),
            .I(N__45830));
    InMux I__10406 (
            .O(N__45849),
            .I(N__45824));
    InMux I__10405 (
            .O(N__45848),
            .I(N__45824));
    Span4Mux_h I__10404 (
            .O(N__45845),
            .I(N__45821));
    InMux I__10403 (
            .O(N__45842),
            .I(N__45818));
    LocalMux I__10402 (
            .O(N__45839),
            .I(N__45809));
    Span4Mux_v I__10401 (
            .O(N__45836),
            .I(N__45809));
    Span4Mux_h I__10400 (
            .O(N__45833),
            .I(N__45809));
    LocalMux I__10399 (
            .O(N__45830),
            .I(N__45809));
    InMux I__10398 (
            .O(N__45829),
            .I(N__45806));
    LocalMux I__10397 (
            .O(N__45824),
            .I(N__45803));
    Span4Mux_v I__10396 (
            .O(N__45821),
            .I(N__45800));
    LocalMux I__10395 (
            .O(N__45818),
            .I(N__45797));
    Span4Mux_h I__10394 (
            .O(N__45809),
            .I(N__45794));
    LocalMux I__10393 (
            .O(N__45806),
            .I(N__45791));
    Span4Mux_h I__10392 (
            .O(N__45803),
            .I(N__45788));
    Sp12to4 I__10391 (
            .O(N__45800),
            .I(N__45785));
    Span4Mux_h I__10390 (
            .O(N__45797),
            .I(N__45782));
    Span4Mux_h I__10389 (
            .O(N__45794),
            .I(N__45775));
    Span4Mux_h I__10388 (
            .O(N__45791),
            .I(N__45775));
    Span4Mux_h I__10387 (
            .O(N__45788),
            .I(N__45775));
    Odrv12 I__10386 (
            .O(N__45785),
            .I(comm_buf_0_2));
    Odrv4 I__10385 (
            .O(N__45782),
            .I(comm_buf_0_2));
    Odrv4 I__10384 (
            .O(N__45775),
            .I(comm_buf_0_2));
    InMux I__10383 (
            .O(N__45768),
            .I(N__45765));
    LocalMux I__10382 (
            .O(N__45765),
            .I(N__45762));
    Span4Mux_v I__10381 (
            .O(N__45762),
            .I(N__45759));
    Span4Mux_h I__10380 (
            .O(N__45759),
            .I(N__45756));
    Odrv4 I__10379 (
            .O(N__45756),
            .I(buf_data_iac_19));
    InMux I__10378 (
            .O(N__45753),
            .I(N__45750));
    LocalMux I__10377 (
            .O(N__45750),
            .I(N__45747));
    Span4Mux_h I__10376 (
            .O(N__45747),
            .I(N__45744));
    Span4Mux_h I__10375 (
            .O(N__45744),
            .I(N__45741));
    Odrv4 I__10374 (
            .O(N__45741),
            .I(n21543));
    IoInMux I__10373 (
            .O(N__45738),
            .I(N__45735));
    LocalMux I__10372 (
            .O(N__45735),
            .I(N__45732));
    IoSpan4Mux I__10371 (
            .O(N__45732),
            .I(N__45729));
    Span4Mux_s3_v I__10370 (
            .O(N__45729),
            .I(N__45725));
    InMux I__10369 (
            .O(N__45728),
            .I(N__45722));
    Sp12to4 I__10368 (
            .O(N__45725),
            .I(N__45719));
    LocalMux I__10367 (
            .O(N__45722),
            .I(N__45715));
    Span12Mux_s11_v I__10366 (
            .O(N__45719),
            .I(N__45712));
    InMux I__10365 (
            .O(N__45718),
            .I(N__45709));
    Span4Mux_h I__10364 (
            .O(N__45715),
            .I(N__45706));
    Odrv12 I__10363 (
            .O(N__45712),
            .I(SELIRNG0));
    LocalMux I__10362 (
            .O(N__45709),
            .I(SELIRNG0));
    Odrv4 I__10361 (
            .O(N__45706),
            .I(SELIRNG0));
    InMux I__10360 (
            .O(N__45699),
            .I(N__45696));
    LocalMux I__10359 (
            .O(N__45696),
            .I(N__45693));
    Span4Mux_h I__10358 (
            .O(N__45693),
            .I(N__45690));
    Odrv4 I__10357 (
            .O(N__45690),
            .I(n23_adj_1685));
    InMux I__10356 (
            .O(N__45687),
            .I(N__45684));
    LocalMux I__10355 (
            .O(N__45684),
            .I(n21273));
    InMux I__10354 (
            .O(N__45681),
            .I(N__45678));
    LocalMux I__10353 (
            .O(N__45678),
            .I(N__45674));
    InMux I__10352 (
            .O(N__45677),
            .I(N__45671));
    Span4Mux_h I__10351 (
            .O(N__45674),
            .I(N__45666));
    LocalMux I__10350 (
            .O(N__45671),
            .I(N__45663));
    InMux I__10349 (
            .O(N__45670),
            .I(N__45658));
    InMux I__10348 (
            .O(N__45669),
            .I(N__45658));
    Odrv4 I__10347 (
            .O(N__45666),
            .I(comm_buf_1_0));
    Odrv4 I__10346 (
            .O(N__45663),
            .I(comm_buf_1_0));
    LocalMux I__10345 (
            .O(N__45658),
            .I(comm_buf_1_0));
    CascadeMux I__10344 (
            .O(N__45651),
            .I(n22533_cascade_));
    InMux I__10343 (
            .O(N__45648),
            .I(N__45642));
    CascadeMux I__10342 (
            .O(N__45647),
            .I(N__45639));
    CascadeMux I__10341 (
            .O(N__45646),
            .I(N__45636));
    CascadeMux I__10340 (
            .O(N__45645),
            .I(N__45631));
    LocalMux I__10339 (
            .O(N__45642),
            .I(N__45628));
    InMux I__10338 (
            .O(N__45639),
            .I(N__45625));
    InMux I__10337 (
            .O(N__45636),
            .I(N__45622));
    CascadeMux I__10336 (
            .O(N__45635),
            .I(N__45617));
    InMux I__10335 (
            .O(N__45634),
            .I(N__45613));
    InMux I__10334 (
            .O(N__45631),
            .I(N__45610));
    Span4Mux_h I__10333 (
            .O(N__45628),
            .I(N__45605));
    LocalMux I__10332 (
            .O(N__45625),
            .I(N__45605));
    LocalMux I__10331 (
            .O(N__45622),
            .I(N__45602));
    InMux I__10330 (
            .O(N__45621),
            .I(N__45599));
    InMux I__10329 (
            .O(N__45620),
            .I(N__45596));
    InMux I__10328 (
            .O(N__45617),
            .I(N__45593));
    InMux I__10327 (
            .O(N__45616),
            .I(N__45590));
    LocalMux I__10326 (
            .O(N__45613),
            .I(N__45585));
    LocalMux I__10325 (
            .O(N__45610),
            .I(N__45585));
    Span4Mux_v I__10324 (
            .O(N__45605),
            .I(N__45582));
    Span4Mux_v I__10323 (
            .O(N__45602),
            .I(N__45579));
    LocalMux I__10322 (
            .O(N__45599),
            .I(N__45576));
    LocalMux I__10321 (
            .O(N__45596),
            .I(N__45573));
    LocalMux I__10320 (
            .O(N__45593),
            .I(N__45568));
    LocalMux I__10319 (
            .O(N__45590),
            .I(N__45568));
    Span4Mux_v I__10318 (
            .O(N__45585),
            .I(N__45563));
    Span4Mux_h I__10317 (
            .O(N__45582),
            .I(N__45563));
    Span4Mux_h I__10316 (
            .O(N__45579),
            .I(N__45554));
    Span4Mux_h I__10315 (
            .O(N__45576),
            .I(N__45554));
    Span4Mux_v I__10314 (
            .O(N__45573),
            .I(N__45554));
    Span4Mux_v I__10313 (
            .O(N__45568),
            .I(N__45554));
    Odrv4 I__10312 (
            .O(N__45563),
            .I(comm_buf_0_0));
    Odrv4 I__10311 (
            .O(N__45554),
            .I(comm_buf_0_0));
    InMux I__10310 (
            .O(N__45549),
            .I(N__45546));
    LocalMux I__10309 (
            .O(N__45546),
            .I(n22536));
    InMux I__10308 (
            .O(N__45543),
            .I(N__45540));
    LocalMux I__10307 (
            .O(N__45540),
            .I(n24_adj_1639));
    CascadeMux I__10306 (
            .O(N__45537),
            .I(n21497_cascade_));
    CascadeMux I__10305 (
            .O(N__45534),
            .I(n34_adj_1649_cascade_));
    InMux I__10304 (
            .O(N__45531),
            .I(N__45528));
    LocalMux I__10303 (
            .O(N__45528),
            .I(n30_adj_1531));
    InMux I__10302 (
            .O(N__45525),
            .I(N__45522));
    LocalMux I__10301 (
            .O(N__45522),
            .I(comm_buf_2_0));
    InMux I__10300 (
            .O(N__45519),
            .I(N__45516));
    LocalMux I__10299 (
            .O(N__45516),
            .I(N__45513));
    Span12Mux_h I__10298 (
            .O(N__45513),
            .I(N__45510));
    Odrv12 I__10297 (
            .O(N__45510),
            .I(n30_adj_1599));
    InMux I__10296 (
            .O(N__45507),
            .I(N__45504));
    LocalMux I__10295 (
            .O(N__45504),
            .I(comm_buf_2_7));
    InMux I__10294 (
            .O(N__45501),
            .I(N__45498));
    LocalMux I__10293 (
            .O(N__45498),
            .I(N__45495));
    Span4Mux_h I__10292 (
            .O(N__45495),
            .I(N__45492));
    Span4Mux_h I__10291 (
            .O(N__45492),
            .I(N__45489));
    Span4Mux_h I__10290 (
            .O(N__45489),
            .I(N__45486));
    Span4Mux_v I__10289 (
            .O(N__45486),
            .I(N__45483));
    Odrv4 I__10288 (
            .O(N__45483),
            .I(n30_adj_1602));
    CascadeMux I__10287 (
            .O(N__45480),
            .I(N__45476));
    InMux I__10286 (
            .O(N__45479),
            .I(N__45472));
    InMux I__10285 (
            .O(N__45476),
            .I(N__45469));
    InMux I__10284 (
            .O(N__45475),
            .I(N__45466));
    LocalMux I__10283 (
            .O(N__45472),
            .I(N__45462));
    LocalMux I__10282 (
            .O(N__45469),
            .I(N__45459));
    LocalMux I__10281 (
            .O(N__45466),
            .I(N__45456));
    InMux I__10280 (
            .O(N__45465),
            .I(N__45453));
    Span4Mux_h I__10279 (
            .O(N__45462),
            .I(N__45450));
    Span4Mux_h I__10278 (
            .O(N__45459),
            .I(N__45445));
    Span4Mux_v I__10277 (
            .O(N__45456),
            .I(N__45445));
    LocalMux I__10276 (
            .O(N__45453),
            .I(N__45442));
    Span4Mux_v I__10275 (
            .O(N__45450),
            .I(N__45439));
    Span4Mux_h I__10274 (
            .O(N__45445),
            .I(N__45434));
    Span4Mux_h I__10273 (
            .O(N__45442),
            .I(N__45434));
    Span4Mux_h I__10272 (
            .O(N__45439),
            .I(N__45431));
    Span4Mux_v I__10271 (
            .O(N__45434),
            .I(N__45428));
    Odrv4 I__10270 (
            .O(N__45431),
            .I(comm_buf_1_2));
    Odrv4 I__10269 (
            .O(N__45428),
            .I(comm_buf_1_2));
    CascadeMux I__10268 (
            .O(N__45423),
            .I(n1_cascade_));
    InMux I__10267 (
            .O(N__45420),
            .I(N__45417));
    LocalMux I__10266 (
            .O(N__45417),
            .I(n2_adj_1584));
    InMux I__10265 (
            .O(N__45414),
            .I(N__45411));
    LocalMux I__10264 (
            .O(N__45411),
            .I(N__45408));
    Odrv12 I__10263 (
            .O(N__45408),
            .I(comm_buf_4_2));
    InMux I__10262 (
            .O(N__45405),
            .I(N__45402));
    LocalMux I__10261 (
            .O(N__45402),
            .I(n21528));
    CascadeMux I__10260 (
            .O(N__45399),
            .I(n4_adj_1585_cascade_));
    InMux I__10259 (
            .O(N__45396),
            .I(N__45393));
    LocalMux I__10258 (
            .O(N__45393),
            .I(n22491));
    CascadeMux I__10257 (
            .O(N__45390),
            .I(N__45385));
    InMux I__10256 (
            .O(N__45389),
            .I(N__45382));
    InMux I__10255 (
            .O(N__45388),
            .I(N__45377));
    InMux I__10254 (
            .O(N__45385),
            .I(N__45377));
    LocalMux I__10253 (
            .O(N__45382),
            .I(N__45374));
    LocalMux I__10252 (
            .O(N__45377),
            .I(N__45371));
    Span4Mux_v I__10251 (
            .O(N__45374),
            .I(N__45366));
    Span4Mux_h I__10250 (
            .O(N__45371),
            .I(N__45366));
    Odrv4 I__10249 (
            .O(N__45366),
            .I(n21143));
    CascadeMux I__10248 (
            .O(N__45363),
            .I(n19193_cascade_));
    CascadeMux I__10247 (
            .O(N__45360),
            .I(n19188_cascade_));
    CascadeMux I__10246 (
            .O(N__45357),
            .I(N__45353));
    CascadeMux I__10245 (
            .O(N__45356),
            .I(N__45349));
    InMux I__10244 (
            .O(N__45353),
            .I(N__45345));
    InMux I__10243 (
            .O(N__45352),
            .I(N__45342));
    InMux I__10242 (
            .O(N__45349),
            .I(N__45339));
    InMux I__10241 (
            .O(N__45348),
            .I(N__45336));
    LocalMux I__10240 (
            .O(N__45345),
            .I(N__45327));
    LocalMux I__10239 (
            .O(N__45342),
            .I(N__45327));
    LocalMux I__10238 (
            .O(N__45339),
            .I(N__45327));
    LocalMux I__10237 (
            .O(N__45336),
            .I(N__45323));
    InMux I__10236 (
            .O(N__45335),
            .I(N__45320));
    InMux I__10235 (
            .O(N__45334),
            .I(N__45317));
    Span4Mux_v I__10234 (
            .O(N__45327),
            .I(N__45314));
    InMux I__10233 (
            .O(N__45326),
            .I(N__45311));
    Span4Mux_h I__10232 (
            .O(N__45323),
            .I(N__45306));
    LocalMux I__10231 (
            .O(N__45320),
            .I(N__45306));
    LocalMux I__10230 (
            .O(N__45317),
            .I(N__45303));
    Span4Mux_h I__10229 (
            .O(N__45314),
            .I(N__45293));
    LocalMux I__10228 (
            .O(N__45311),
            .I(N__45293));
    Span4Mux_h I__10227 (
            .O(N__45306),
            .I(N__45293));
    Span4Mux_h I__10226 (
            .O(N__45303),
            .I(N__45293));
    InMux I__10225 (
            .O(N__45302),
            .I(N__45290));
    Odrv4 I__10224 (
            .O(N__45293),
            .I(comm_buf_0_3));
    LocalMux I__10223 (
            .O(N__45290),
            .I(comm_buf_0_3));
    CascadeMux I__10222 (
            .O(N__45285),
            .I(n22557_cascade_));
    InMux I__10221 (
            .O(N__45282),
            .I(N__45275));
    InMux I__10220 (
            .O(N__45281),
            .I(N__45275));
    InMux I__10219 (
            .O(N__45280),
            .I(N__45272));
    LocalMux I__10218 (
            .O(N__45275),
            .I(N__45269));
    LocalMux I__10217 (
            .O(N__45272),
            .I(N__45266));
    Span4Mux_h I__10216 (
            .O(N__45269),
            .I(N__45263));
    Span4Mux_h I__10215 (
            .O(N__45266),
            .I(N__45260));
    Span4Mux_h I__10214 (
            .O(N__45263),
            .I(N__45257));
    Odrv4 I__10213 (
            .O(N__45260),
            .I(comm_buf_1_3));
    Odrv4 I__10212 (
            .O(N__45257),
            .I(comm_buf_1_3));
    InMux I__10211 (
            .O(N__45252),
            .I(N__45249));
    LocalMux I__10210 (
            .O(N__45249),
            .I(N__45246));
    Odrv12 I__10209 (
            .O(N__45246),
            .I(comm_buf_4_3));
    CascadeMux I__10208 (
            .O(N__45243),
            .I(n4_adj_1583_cascade_));
    InMux I__10207 (
            .O(N__45240),
            .I(N__45237));
    LocalMux I__10206 (
            .O(N__45237),
            .I(n22560));
    CascadeMux I__10205 (
            .O(N__45234),
            .I(n21288_cascade_));
    InMux I__10204 (
            .O(N__45231),
            .I(N__45228));
    LocalMux I__10203 (
            .O(N__45228),
            .I(N__45225));
    Span4Mux_h I__10202 (
            .O(N__45225),
            .I(N__45222));
    Odrv4 I__10201 (
            .O(N__45222),
            .I(n21479));
    CascadeMux I__10200 (
            .O(N__45219),
            .I(n21477_cascade_));
    CascadeMux I__10199 (
            .O(N__45216),
            .I(n44_cascade_));
    CEMux I__10198 (
            .O(N__45213),
            .I(N__45206));
    CEMux I__10197 (
            .O(N__45212),
            .I(N__45203));
    CEMux I__10196 (
            .O(N__45211),
            .I(N__45200));
    CEMux I__10195 (
            .O(N__45210),
            .I(N__45196));
    CEMux I__10194 (
            .O(N__45209),
            .I(N__45191));
    LocalMux I__10193 (
            .O(N__45206),
            .I(N__45186));
    LocalMux I__10192 (
            .O(N__45203),
            .I(N__45186));
    LocalMux I__10191 (
            .O(N__45200),
            .I(N__45183));
    CEMux I__10190 (
            .O(N__45199),
            .I(N__45180));
    LocalMux I__10189 (
            .O(N__45196),
            .I(N__45177));
    CEMux I__10188 (
            .O(N__45195),
            .I(N__45174));
    CEMux I__10187 (
            .O(N__45194),
            .I(N__45171));
    LocalMux I__10186 (
            .O(N__45191),
            .I(N__45167));
    Span4Mux_v I__10185 (
            .O(N__45186),
            .I(N__45164));
    Span4Mux_v I__10184 (
            .O(N__45183),
            .I(N__45157));
    LocalMux I__10183 (
            .O(N__45180),
            .I(N__45157));
    Span4Mux_v I__10182 (
            .O(N__45177),
            .I(N__45157));
    LocalMux I__10181 (
            .O(N__45174),
            .I(N__45154));
    LocalMux I__10180 (
            .O(N__45171),
            .I(N__45151));
    InMux I__10179 (
            .O(N__45170),
            .I(N__45148));
    Span4Mux_h I__10178 (
            .O(N__45167),
            .I(N__45145));
    Span4Mux_h I__10177 (
            .O(N__45164),
            .I(N__45140));
    Span4Mux_v I__10176 (
            .O(N__45157),
            .I(N__45140));
    Span4Mux_h I__10175 (
            .O(N__45154),
            .I(N__45133));
    Span4Mux_v I__10174 (
            .O(N__45151),
            .I(N__45133));
    LocalMux I__10173 (
            .O(N__45148),
            .I(N__45133));
    Odrv4 I__10172 (
            .O(N__45145),
            .I(n12260));
    Odrv4 I__10171 (
            .O(N__45140),
            .I(n12260));
    Odrv4 I__10170 (
            .O(N__45133),
            .I(n12260));
    InMux I__10169 (
            .O(N__45126),
            .I(N__45123));
    LocalMux I__10168 (
            .O(N__45123),
            .I(N__45120));
    Span4Mux_h I__10167 (
            .O(N__45120),
            .I(N__45117));
    Span4Mux_v I__10166 (
            .O(N__45117),
            .I(N__45114));
    Span4Mux_v I__10165 (
            .O(N__45114),
            .I(N__45111));
    Odrv4 I__10164 (
            .O(N__45111),
            .I(buf_data_vac_10));
    InMux I__10163 (
            .O(N__45108),
            .I(N__45105));
    LocalMux I__10162 (
            .O(N__45105),
            .I(N__45102));
    Span4Mux_h I__10161 (
            .O(N__45102),
            .I(N__45099));
    Span4Mux_v I__10160 (
            .O(N__45099),
            .I(N__45096));
    Span4Mux_v I__10159 (
            .O(N__45096),
            .I(N__45093));
    Odrv4 I__10158 (
            .O(N__45093),
            .I(buf_data_vac_9));
    SRMux I__10157 (
            .O(N__45090),
            .I(N__45087));
    LocalMux I__10156 (
            .O(N__45087),
            .I(N__45084));
    Span4Mux_h I__10155 (
            .O(N__45084),
            .I(N__45081));
    Odrv4 I__10154 (
            .O(N__45081),
            .I(n14986));
    CascadeMux I__10153 (
            .O(N__45078),
            .I(n21268_cascade_));
    InMux I__10152 (
            .O(N__45075),
            .I(N__45072));
    LocalMux I__10151 (
            .O(N__45072),
            .I(n22094));
    CascadeMux I__10150 (
            .O(N__45069),
            .I(N__45066));
    InMux I__10149 (
            .O(N__45066),
            .I(N__45063));
    LocalMux I__10148 (
            .O(N__45063),
            .I(n21266));
    CEMux I__10147 (
            .O(N__45060),
            .I(N__45056));
    InMux I__10146 (
            .O(N__45059),
            .I(N__45053));
    LocalMux I__10145 (
            .O(N__45056),
            .I(N__45050));
    LocalMux I__10144 (
            .O(N__45053),
            .I(N__45047));
    Odrv12 I__10143 (
            .O(N__45050),
            .I(n12407));
    Odrv4 I__10142 (
            .O(N__45047),
            .I(n12407));
    CascadeMux I__10141 (
            .O(N__45042),
            .I(n21085_cascade_));
    InMux I__10140 (
            .O(N__45039),
            .I(N__45036));
    LocalMux I__10139 (
            .O(N__45036),
            .I(n19188));
    InMux I__10138 (
            .O(N__45033),
            .I(N__45029));
    InMux I__10137 (
            .O(N__45032),
            .I(N__45026));
    LocalMux I__10136 (
            .O(N__45029),
            .I(N__45020));
    LocalMux I__10135 (
            .O(N__45026),
            .I(N__45020));
    InMux I__10134 (
            .O(N__45025),
            .I(N__45017));
    Span4Mux_v I__10133 (
            .O(N__45020),
            .I(N__45011));
    LocalMux I__10132 (
            .O(N__45017),
            .I(N__45011));
    InMux I__10131 (
            .O(N__45016),
            .I(N__45008));
    Span4Mux_h I__10130 (
            .O(N__45011),
            .I(N__45005));
    LocalMux I__10129 (
            .O(N__45008),
            .I(\comm_spi.n23092 ));
    Odrv4 I__10128 (
            .O(N__45005),
            .I(\comm_spi.n23092 ));
    InMux I__10127 (
            .O(N__45000),
            .I(N__44997));
    LocalMux I__10126 (
            .O(N__44997),
            .I(N__44994));
    Span4Mux_v I__10125 (
            .O(N__44994),
            .I(N__44989));
    InMux I__10124 (
            .O(N__44993),
            .I(N__44986));
    InMux I__10123 (
            .O(N__44992),
            .I(N__44983));
    Odrv4 I__10122 (
            .O(N__44989),
            .I(clk_cnt_1));
    LocalMux I__10121 (
            .O(N__44986),
            .I(clk_cnt_1));
    LocalMux I__10120 (
            .O(N__44983),
            .I(clk_cnt_1));
    InMux I__10119 (
            .O(N__44976),
            .I(N__44973));
    LocalMux I__10118 (
            .O(N__44973),
            .I(N__44970));
    Span4Mux_v I__10117 (
            .O(N__44970),
            .I(N__44964));
    InMux I__10116 (
            .O(N__44969),
            .I(N__44959));
    InMux I__10115 (
            .O(N__44968),
            .I(N__44959));
    InMux I__10114 (
            .O(N__44967),
            .I(N__44956));
    Odrv4 I__10113 (
            .O(N__44964),
            .I(clk_cnt_0));
    LocalMux I__10112 (
            .O(N__44959),
            .I(clk_cnt_0));
    LocalMux I__10111 (
            .O(N__44956),
            .I(clk_cnt_0));
    SRMux I__10110 (
            .O(N__44949),
            .I(N__44946));
    LocalMux I__10109 (
            .O(N__44946),
            .I(N__44943));
    Odrv4 I__10108 (
            .O(N__44943),
            .I(n17773));
    InMux I__10107 (
            .O(N__44940),
            .I(N__44937));
    LocalMux I__10106 (
            .O(N__44937),
            .I(N__44934));
    Span4Mux_h I__10105 (
            .O(N__44934),
            .I(N__44931));
    Span4Mux_v I__10104 (
            .O(N__44931),
            .I(N__44928));
    Sp12to4 I__10103 (
            .O(N__44928),
            .I(N__44925));
    Odrv12 I__10102 (
            .O(N__44925),
            .I(buf_data_vac_8));
    InMux I__10101 (
            .O(N__44922),
            .I(N__44919));
    LocalMux I__10100 (
            .O(N__44919),
            .I(N__44916));
    Span4Mux_h I__10099 (
            .O(N__44916),
            .I(N__44913));
    Span4Mux_v I__10098 (
            .O(N__44913),
            .I(N__44910));
    Odrv4 I__10097 (
            .O(N__44910),
            .I(buf_data_vac_15));
    InMux I__10096 (
            .O(N__44907),
            .I(N__44904));
    LocalMux I__10095 (
            .O(N__44904),
            .I(comm_buf_4_7));
    InMux I__10094 (
            .O(N__44901),
            .I(N__44898));
    LocalMux I__10093 (
            .O(N__44898),
            .I(N__44895));
    Span12Mux_h I__10092 (
            .O(N__44895),
            .I(N__44892));
    Odrv12 I__10091 (
            .O(N__44892),
            .I(buf_data_vac_14));
    InMux I__10090 (
            .O(N__44889),
            .I(N__44886));
    LocalMux I__10089 (
            .O(N__44886),
            .I(N__44883));
    Span4Mux_h I__10088 (
            .O(N__44883),
            .I(N__44880));
    Span4Mux_v I__10087 (
            .O(N__44880),
            .I(N__44877));
    Odrv4 I__10086 (
            .O(N__44877),
            .I(buf_data_vac_13));
    InMux I__10085 (
            .O(N__44874),
            .I(N__44871));
    LocalMux I__10084 (
            .O(N__44871),
            .I(N__44868));
    Span4Mux_h I__10083 (
            .O(N__44868),
            .I(N__44865));
    Span4Mux_v I__10082 (
            .O(N__44865),
            .I(N__44862));
    Span4Mux_v I__10081 (
            .O(N__44862),
            .I(N__44859));
    Odrv4 I__10080 (
            .O(N__44859),
            .I(buf_data_vac_12));
    InMux I__10079 (
            .O(N__44856),
            .I(N__44853));
    LocalMux I__10078 (
            .O(N__44853),
            .I(N__44850));
    Odrv4 I__10077 (
            .O(N__44850),
            .I(comm_buf_4_4));
    InMux I__10076 (
            .O(N__44847),
            .I(N__44844));
    LocalMux I__10075 (
            .O(N__44844),
            .I(N__44841));
    Span4Mux_v I__10074 (
            .O(N__44841),
            .I(N__44838));
    Span4Mux_v I__10073 (
            .O(N__44838),
            .I(N__44835));
    Span4Mux_h I__10072 (
            .O(N__44835),
            .I(N__44832));
    Odrv4 I__10071 (
            .O(N__44832),
            .I(buf_data_vac_11));
    InMux I__10070 (
            .O(N__44829),
            .I(N__44826));
    LocalMux I__10069 (
            .O(N__44826),
            .I(N__44823));
    Span4Mux_v I__10068 (
            .O(N__44823),
            .I(N__44819));
    InMux I__10067 (
            .O(N__44822),
            .I(N__44816));
    Span4Mux_v I__10066 (
            .O(N__44819),
            .I(N__44810));
    LocalMux I__10065 (
            .O(N__44816),
            .I(N__44810));
    InMux I__10064 (
            .O(N__44815),
            .I(N__44807));
    Span4Mux_v I__10063 (
            .O(N__44810),
            .I(N__44804));
    LocalMux I__10062 (
            .O(N__44807),
            .I(wdtick_flag));
    Odrv4 I__10061 (
            .O(N__44804),
            .I(wdtick_flag));
    InMux I__10060 (
            .O(N__44799),
            .I(N__44796));
    LocalMux I__10059 (
            .O(N__44796),
            .I(N__44793));
    Span4Mux_v I__10058 (
            .O(N__44793),
            .I(N__44788));
    InMux I__10057 (
            .O(N__44792),
            .I(N__44785));
    InMux I__10056 (
            .O(N__44791),
            .I(N__44782));
    Odrv4 I__10055 (
            .O(N__44788),
            .I(buf_control_0));
    LocalMux I__10054 (
            .O(N__44785),
            .I(buf_control_0));
    LocalMux I__10053 (
            .O(N__44782),
            .I(buf_control_0));
    IoInMux I__10052 (
            .O(N__44775),
            .I(N__44772));
    LocalMux I__10051 (
            .O(N__44772),
            .I(N__44769));
    Span4Mux_s1_v I__10050 (
            .O(N__44769),
            .I(N__44766));
    Span4Mux_h I__10049 (
            .O(N__44766),
            .I(N__44763));
    Span4Mux_v I__10048 (
            .O(N__44763),
            .I(N__44760));
    Span4Mux_v I__10047 (
            .O(N__44760),
            .I(N__44757));
    Odrv4 I__10046 (
            .O(N__44757),
            .I(CONT_SD));
    InMux I__10045 (
            .O(N__44754),
            .I(N__44749));
    CascadeMux I__10044 (
            .O(N__44753),
            .I(N__44745));
    InMux I__10043 (
            .O(N__44752),
            .I(N__44741));
    LocalMux I__10042 (
            .O(N__44749),
            .I(N__44738));
    InMux I__10041 (
            .O(N__44748),
            .I(N__44735));
    InMux I__10040 (
            .O(N__44745),
            .I(N__44730));
    InMux I__10039 (
            .O(N__44744),
            .I(N__44730));
    LocalMux I__10038 (
            .O(N__44741),
            .I(N__44727));
    Span4Mux_v I__10037 (
            .O(N__44738),
            .I(N__44719));
    LocalMux I__10036 (
            .O(N__44735),
            .I(N__44719));
    LocalMux I__10035 (
            .O(N__44730),
            .I(N__44719));
    Span4Mux_v I__10034 (
            .O(N__44727),
            .I(N__44716));
    InMux I__10033 (
            .O(N__44726),
            .I(N__44713));
    Span4Mux_h I__10032 (
            .O(N__44719),
            .I(N__44710));
    Sp12to4 I__10031 (
            .O(N__44716),
            .I(N__44703));
    LocalMux I__10030 (
            .O(N__44713),
            .I(N__44703));
    Span4Mux_h I__10029 (
            .O(N__44710),
            .I(N__44699));
    InMux I__10028 (
            .O(N__44709),
            .I(N__44696));
    InMux I__10027 (
            .O(N__44708),
            .I(N__44693));
    Span12Mux_v I__10026 (
            .O(N__44703),
            .I(N__44690));
    InMux I__10025 (
            .O(N__44702),
            .I(N__44687));
    Span4Mux_v I__10024 (
            .O(N__44699),
            .I(N__44684));
    LocalMux I__10023 (
            .O(N__44696),
            .I(N__44679));
    LocalMux I__10022 (
            .O(N__44693),
            .I(N__44679));
    Odrv12 I__10021 (
            .O(N__44690),
            .I(dds_state_0));
    LocalMux I__10020 (
            .O(N__44687),
            .I(dds_state_0));
    Odrv4 I__10019 (
            .O(N__44684),
            .I(dds_state_0));
    Odrv12 I__10018 (
            .O(N__44679),
            .I(dds_state_0));
    InMux I__10017 (
            .O(N__44670),
            .I(N__44664));
    InMux I__10016 (
            .O(N__44669),
            .I(N__44661));
    InMux I__10015 (
            .O(N__44668),
            .I(N__44658));
    InMux I__10014 (
            .O(N__44667),
            .I(N__44654));
    LocalMux I__10013 (
            .O(N__44664),
            .I(N__44633));
    LocalMux I__10012 (
            .O(N__44661),
            .I(N__44633));
    LocalMux I__10011 (
            .O(N__44658),
            .I(N__44630));
    InMux I__10010 (
            .O(N__44657),
            .I(N__44623));
    LocalMux I__10009 (
            .O(N__44654),
            .I(N__44620));
    InMux I__10008 (
            .O(N__44653),
            .I(N__44617));
    InMux I__10007 (
            .O(N__44652),
            .I(N__44602));
    InMux I__10006 (
            .O(N__44651),
            .I(N__44602));
    InMux I__10005 (
            .O(N__44650),
            .I(N__44602));
    InMux I__10004 (
            .O(N__44649),
            .I(N__44602));
    InMux I__10003 (
            .O(N__44648),
            .I(N__44602));
    InMux I__10002 (
            .O(N__44647),
            .I(N__44602));
    InMux I__10001 (
            .O(N__44646),
            .I(N__44602));
    InMux I__10000 (
            .O(N__44645),
            .I(N__44585));
    InMux I__9999 (
            .O(N__44644),
            .I(N__44585));
    InMux I__9998 (
            .O(N__44643),
            .I(N__44585));
    InMux I__9997 (
            .O(N__44642),
            .I(N__44585));
    InMux I__9996 (
            .O(N__44641),
            .I(N__44585));
    InMux I__9995 (
            .O(N__44640),
            .I(N__44585));
    InMux I__9994 (
            .O(N__44639),
            .I(N__44585));
    InMux I__9993 (
            .O(N__44638),
            .I(N__44585));
    Span4Mux_h I__9992 (
            .O(N__44633),
            .I(N__44582));
    Span4Mux_v I__9991 (
            .O(N__44630),
            .I(N__44579));
    InMux I__9990 (
            .O(N__44629),
            .I(N__44570));
    InMux I__9989 (
            .O(N__44628),
            .I(N__44570));
    InMux I__9988 (
            .O(N__44627),
            .I(N__44570));
    InMux I__9987 (
            .O(N__44626),
            .I(N__44570));
    LocalMux I__9986 (
            .O(N__44623),
            .I(N__44565));
    Span12Mux_v I__9985 (
            .O(N__44620),
            .I(N__44565));
    LocalMux I__9984 (
            .O(N__44617),
            .I(dds_state_2));
    LocalMux I__9983 (
            .O(N__44602),
            .I(dds_state_2));
    LocalMux I__9982 (
            .O(N__44585),
            .I(dds_state_2));
    Odrv4 I__9981 (
            .O(N__44582),
            .I(dds_state_2));
    Odrv4 I__9980 (
            .O(N__44579),
            .I(dds_state_2));
    LocalMux I__9979 (
            .O(N__44570),
            .I(dds_state_2));
    Odrv12 I__9978 (
            .O(N__44565),
            .I(dds_state_2));
    CEMux I__9977 (
            .O(N__44550),
            .I(N__44547));
    LocalMux I__9976 (
            .O(N__44547),
            .I(N__44544));
    Span4Mux_v I__9975 (
            .O(N__44544),
            .I(N__44540));
    CEMux I__9974 (
            .O(N__44543),
            .I(N__44537));
    Span4Mux_h I__9973 (
            .O(N__44540),
            .I(N__44534));
    LocalMux I__9972 (
            .O(N__44537),
            .I(N__44531));
    Span4Mux_h I__9971 (
            .O(N__44534),
            .I(N__44528));
    Span4Mux_v I__9970 (
            .O(N__44531),
            .I(N__44525));
    Span4Mux_v I__9969 (
            .O(N__44528),
            .I(N__44520));
    Span4Mux_h I__9968 (
            .O(N__44525),
            .I(N__44520));
    Odrv4 I__9967 (
            .O(N__44520),
            .I(\SIG_DDS.n9 ));
    CEMux I__9966 (
            .O(N__44517),
            .I(N__44512));
    InMux I__9965 (
            .O(N__44516),
            .I(N__44509));
    InMux I__9964 (
            .O(N__44515),
            .I(N__44505));
    LocalMux I__9963 (
            .O(N__44512),
            .I(N__44500));
    LocalMux I__9962 (
            .O(N__44509),
            .I(N__44488));
    InMux I__9961 (
            .O(N__44508),
            .I(N__44485));
    LocalMux I__9960 (
            .O(N__44505),
            .I(N__44482));
    InMux I__9959 (
            .O(N__44504),
            .I(N__44479));
    SRMux I__9958 (
            .O(N__44503),
            .I(N__44476));
    Span4Mux_v I__9957 (
            .O(N__44500),
            .I(N__44473));
    InMux I__9956 (
            .O(N__44499),
            .I(N__44456));
    InMux I__9955 (
            .O(N__44498),
            .I(N__44456));
    InMux I__9954 (
            .O(N__44497),
            .I(N__44456));
    InMux I__9953 (
            .O(N__44496),
            .I(N__44456));
    InMux I__9952 (
            .O(N__44495),
            .I(N__44456));
    InMux I__9951 (
            .O(N__44494),
            .I(N__44456));
    InMux I__9950 (
            .O(N__44493),
            .I(N__44456));
    InMux I__9949 (
            .O(N__44492),
            .I(N__44456));
    CascadeMux I__9948 (
            .O(N__44491),
            .I(N__44446));
    Span4Mux_h I__9947 (
            .O(N__44488),
            .I(N__44439));
    LocalMux I__9946 (
            .O(N__44485),
            .I(N__44439));
    Span4Mux_v I__9945 (
            .O(N__44482),
            .I(N__44436));
    LocalMux I__9944 (
            .O(N__44479),
            .I(N__44433));
    LocalMux I__9943 (
            .O(N__44476),
            .I(N__44430));
    Span4Mux_h I__9942 (
            .O(N__44473),
            .I(N__44425));
    LocalMux I__9941 (
            .O(N__44456),
            .I(N__44425));
    InMux I__9940 (
            .O(N__44455),
            .I(N__44410));
    InMux I__9939 (
            .O(N__44454),
            .I(N__44410));
    InMux I__9938 (
            .O(N__44453),
            .I(N__44410));
    InMux I__9937 (
            .O(N__44452),
            .I(N__44410));
    InMux I__9936 (
            .O(N__44451),
            .I(N__44410));
    InMux I__9935 (
            .O(N__44450),
            .I(N__44410));
    InMux I__9934 (
            .O(N__44449),
            .I(N__44410));
    InMux I__9933 (
            .O(N__44446),
            .I(N__44401));
    InMux I__9932 (
            .O(N__44445),
            .I(N__44401));
    InMux I__9931 (
            .O(N__44444),
            .I(N__44401));
    Span4Mux_v I__9930 (
            .O(N__44439),
            .I(N__44394));
    Span4Mux_h I__9929 (
            .O(N__44436),
            .I(N__44394));
    Span4Mux_h I__9928 (
            .O(N__44433),
            .I(N__44394));
    Span4Mux_h I__9927 (
            .O(N__44430),
            .I(N__44389));
    Span4Mux_v I__9926 (
            .O(N__44425),
            .I(N__44389));
    LocalMux I__9925 (
            .O(N__44410),
            .I(N__44385));
    InMux I__9924 (
            .O(N__44409),
            .I(N__44380));
    InMux I__9923 (
            .O(N__44408),
            .I(N__44380));
    LocalMux I__9922 (
            .O(N__44401),
            .I(N__44377));
    Span4Mux_h I__9921 (
            .O(N__44394),
            .I(N__44373));
    Span4Mux_h I__9920 (
            .O(N__44389),
            .I(N__44370));
    InMux I__9919 (
            .O(N__44388),
            .I(N__44367));
    Span4Mux_h I__9918 (
            .O(N__44385),
            .I(N__44360));
    LocalMux I__9917 (
            .O(N__44380),
            .I(N__44360));
    Span4Mux_v I__9916 (
            .O(N__44377),
            .I(N__44360));
    InMux I__9915 (
            .O(N__44376),
            .I(N__44357));
    Span4Mux_h I__9914 (
            .O(N__44373),
            .I(N__44354));
    Odrv4 I__9913 (
            .O(N__44370),
            .I(dds_state_1));
    LocalMux I__9912 (
            .O(N__44367),
            .I(dds_state_1));
    Odrv4 I__9911 (
            .O(N__44360),
            .I(dds_state_1));
    LocalMux I__9910 (
            .O(N__44357),
            .I(dds_state_1));
    Odrv4 I__9909 (
            .O(N__44354),
            .I(dds_state_1));
    InMux I__9908 (
            .O(N__44343),
            .I(N__44340));
    LocalMux I__9907 (
            .O(N__44340),
            .I(\comm_spi.n14813 ));
    InMux I__9906 (
            .O(N__44337),
            .I(N__44334));
    LocalMux I__9905 (
            .O(N__44334),
            .I(\comm_spi.n14812 ));
    InMux I__9904 (
            .O(N__44331),
            .I(N__44327));
    InMux I__9903 (
            .O(N__44330),
            .I(N__44324));
    LocalMux I__9902 (
            .O(N__44327),
            .I(N__44320));
    LocalMux I__9901 (
            .O(N__44324),
            .I(N__44317));
    InMux I__9900 (
            .O(N__44323),
            .I(N__44314));
    Span4Mux_h I__9899 (
            .O(N__44320),
            .I(N__44304));
    Span4Mux_h I__9898 (
            .O(N__44317),
            .I(N__44304));
    LocalMux I__9897 (
            .O(N__44314),
            .I(N__44304));
    InMux I__9896 (
            .O(N__44313),
            .I(N__44301));
    InMux I__9895 (
            .O(N__44312),
            .I(N__44298));
    InMux I__9894 (
            .O(N__44311),
            .I(N__44295));
    Sp12to4 I__9893 (
            .O(N__44304),
            .I(N__44288));
    LocalMux I__9892 (
            .O(N__44301),
            .I(N__44288));
    LocalMux I__9891 (
            .O(N__44298),
            .I(N__44288));
    LocalMux I__9890 (
            .O(N__44295),
            .I(\comm_spi.n14811 ));
    Odrv12 I__9889 (
            .O(N__44288),
            .I(\comm_spi.n14811 ));
    IoInMux I__9888 (
            .O(N__44283),
            .I(N__44280));
    LocalMux I__9887 (
            .O(N__44280),
            .I(N__44277));
    IoSpan4Mux I__9886 (
            .O(N__44277),
            .I(N__44274));
    IoSpan4Mux I__9885 (
            .O(N__44274),
            .I(N__44271));
    Span4Mux_s3_h I__9884 (
            .O(N__44271),
            .I(N__44268));
    Span4Mux_h I__9883 (
            .O(N__44268),
            .I(N__44265));
    Odrv4 I__9882 (
            .O(N__44265),
            .I(ICE_SPI_MISO));
    InMux I__9881 (
            .O(N__44262),
            .I(N__44259));
    LocalMux I__9880 (
            .O(N__44259),
            .I(\ADC_VDC.n11895 ));
    InMux I__9879 (
            .O(N__44256),
            .I(N__44253));
    LocalMux I__9878 (
            .O(N__44253),
            .I(\comm_spi.n23086 ));
    CascadeMux I__9877 (
            .O(N__44250),
            .I(\comm_spi.n23086_cascade_ ));
    InMux I__9876 (
            .O(N__44247),
            .I(N__44244));
    LocalMux I__9875 (
            .O(N__44244),
            .I(\comm_spi.n14804 ));
    InMux I__9874 (
            .O(N__44241),
            .I(N__44238));
    LocalMux I__9873 (
            .O(N__44238),
            .I(n80));
    CascadeMux I__9872 (
            .O(N__44235),
            .I(N__44232));
    InMux I__9871 (
            .O(N__44232),
            .I(N__44229));
    LocalMux I__9870 (
            .O(N__44229),
            .I(N__44226));
    Span4Mux_h I__9869 (
            .O(N__44226),
            .I(N__44223));
    Span4Mux_h I__9868 (
            .O(N__44223),
            .I(N__44220));
    Odrv4 I__9867 (
            .O(N__44220),
            .I(n5));
    InMux I__9866 (
            .O(N__44217),
            .I(N__44214));
    LocalMux I__9865 (
            .O(N__44214),
            .I(N__44210));
    InMux I__9864 (
            .O(N__44213),
            .I(N__44207));
    Span12Mux_v I__9863 (
            .O(N__44210),
            .I(N__44204));
    LocalMux I__9862 (
            .O(N__44207),
            .I(data_idxvec_1));
    Odrv12 I__9861 (
            .O(N__44204),
            .I(data_idxvec_1));
    InMux I__9860 (
            .O(N__44199),
            .I(N__44196));
    LocalMux I__9859 (
            .O(N__44196),
            .I(N__44191));
    InMux I__9858 (
            .O(N__44195),
            .I(N__44188));
    InMux I__9857 (
            .O(N__44194),
            .I(N__44185));
    Span4Mux_h I__9856 (
            .O(N__44191),
            .I(N__44182));
    LocalMux I__9855 (
            .O(N__44188),
            .I(data_cntvec_1));
    LocalMux I__9854 (
            .O(N__44185),
            .I(data_cntvec_1));
    Odrv4 I__9853 (
            .O(N__44182),
            .I(data_cntvec_1));
    CascadeMux I__9852 (
            .O(N__44175),
            .I(n26_adj_1653_cascade_));
    InMux I__9851 (
            .O(N__44172),
            .I(N__44169));
    LocalMux I__9850 (
            .O(N__44169),
            .I(N__44166));
    Span4Mux_v I__9849 (
            .O(N__44166),
            .I(N__44161));
    InMux I__9848 (
            .O(N__44165),
            .I(N__44156));
    InMux I__9847 (
            .O(N__44164),
            .I(N__44156));
    Odrv4 I__9846 (
            .O(N__44161),
            .I(acadc_skipCount_1));
    LocalMux I__9845 (
            .O(N__44156),
            .I(acadc_skipCount_1));
    CascadeMux I__9844 (
            .O(N__44151),
            .I(n22497_cascade_));
    InMux I__9843 (
            .O(N__44148),
            .I(N__44145));
    LocalMux I__9842 (
            .O(N__44145),
            .I(N__44142));
    Span4Mux_h I__9841 (
            .O(N__44142),
            .I(N__44137));
    InMux I__9840 (
            .O(N__44141),
            .I(N__44132));
    InMux I__9839 (
            .O(N__44140),
            .I(N__44132));
    Odrv4 I__9838 (
            .O(N__44137),
            .I(req_data_cnt_1));
    LocalMux I__9837 (
            .O(N__44132),
            .I(req_data_cnt_1));
    InMux I__9836 (
            .O(N__44127),
            .I(N__44124));
    LocalMux I__9835 (
            .O(N__44124),
            .I(n22434));
    CascadeMux I__9834 (
            .O(N__44121),
            .I(n22500_cascade_));
    CascadeMux I__9833 (
            .O(N__44118),
            .I(n30_adj_1654_cascade_));
    CascadeMux I__9832 (
            .O(N__44115),
            .I(N__44111));
    InMux I__9831 (
            .O(N__44114),
            .I(N__44108));
    InMux I__9830 (
            .O(N__44111),
            .I(N__44105));
    LocalMux I__9829 (
            .O(N__44108),
            .I(N__44102));
    LocalMux I__9828 (
            .O(N__44105),
            .I(N__44099));
    Span4Mux_h I__9827 (
            .O(N__44102),
            .I(N__44096));
    Span4Mux_v I__9826 (
            .O(N__44099),
            .I(N__44093));
    Span4Mux_v I__9825 (
            .O(N__44096),
            .I(N__44090));
    Span4Mux_h I__9824 (
            .O(N__44093),
            .I(N__44087));
    Odrv4 I__9823 (
            .O(N__44090),
            .I(n28));
    Odrv4 I__9822 (
            .O(N__44087),
            .I(n28));
    CascadeMux I__9821 (
            .O(N__44082),
            .I(N__44079));
    InMux I__9820 (
            .O(N__44079),
            .I(N__44075));
    CascadeMux I__9819 (
            .O(N__44078),
            .I(N__44072));
    LocalMux I__9818 (
            .O(N__44075),
            .I(N__44068));
    InMux I__9817 (
            .O(N__44072),
            .I(N__44065));
    InMux I__9816 (
            .O(N__44071),
            .I(N__44062));
    Span4Mux_h I__9815 (
            .O(N__44068),
            .I(N__44054));
    LocalMux I__9814 (
            .O(N__44065),
            .I(N__44054));
    LocalMux I__9813 (
            .O(N__44062),
            .I(N__44051));
    InMux I__9812 (
            .O(N__44061),
            .I(N__44048));
    InMux I__9811 (
            .O(N__44060),
            .I(N__44043));
    InMux I__9810 (
            .O(N__44059),
            .I(N__44043));
    Span4Mux_v I__9809 (
            .O(N__44054),
            .I(N__44040));
    Span4Mux_h I__9808 (
            .O(N__44051),
            .I(N__44037));
    LocalMux I__9807 (
            .O(N__44048),
            .I(N__44032));
    LocalMux I__9806 (
            .O(N__44043),
            .I(N__44032));
    Span4Mux_h I__9805 (
            .O(N__44040),
            .I(N__44029));
    Span4Mux_v I__9804 (
            .O(N__44037),
            .I(N__44026));
    Span12Mux_v I__9803 (
            .O(N__44032),
            .I(N__44023));
    Odrv4 I__9802 (
            .O(N__44029),
            .I(comm_buf_1_7));
    Odrv4 I__9801 (
            .O(N__44026),
            .I(comm_buf_1_7));
    Odrv12 I__9800 (
            .O(N__44023),
            .I(comm_buf_1_7));
    SRMux I__9799 (
            .O(N__44016),
            .I(N__44010));
    SRMux I__9798 (
            .O(N__44015),
            .I(N__44006));
    SRMux I__9797 (
            .O(N__44014),
            .I(N__44003));
    SRMux I__9796 (
            .O(N__44013),
            .I(N__43998));
    LocalMux I__9795 (
            .O(N__44010),
            .I(N__43995));
    SRMux I__9794 (
            .O(N__44009),
            .I(N__43992));
    LocalMux I__9793 (
            .O(N__44006),
            .I(N__43989));
    LocalMux I__9792 (
            .O(N__44003),
            .I(N__43986));
    SRMux I__9791 (
            .O(N__44002),
            .I(N__43983));
    SRMux I__9790 (
            .O(N__44001),
            .I(N__43980));
    LocalMux I__9789 (
            .O(N__43998),
            .I(N__43973));
    Span4Mux_h I__9788 (
            .O(N__43995),
            .I(N__43973));
    LocalMux I__9787 (
            .O(N__43992),
            .I(N__43973));
    Span4Mux_h I__9786 (
            .O(N__43989),
            .I(N__43966));
    Span4Mux_v I__9785 (
            .O(N__43986),
            .I(N__43966));
    LocalMux I__9784 (
            .O(N__43983),
            .I(N__43966));
    LocalMux I__9783 (
            .O(N__43980),
            .I(N__43963));
    Span4Mux_v I__9782 (
            .O(N__43973),
            .I(N__43957));
    Span4Mux_h I__9781 (
            .O(N__43966),
            .I(N__43957));
    Span4Mux_h I__9780 (
            .O(N__43963),
            .I(N__43954));
    SRMux I__9779 (
            .O(N__43962),
            .I(N__43951));
    Odrv4 I__9778 (
            .O(N__43957),
            .I(n14965));
    Odrv4 I__9777 (
            .O(N__43954),
            .I(n14965));
    LocalMux I__9776 (
            .O(N__43951),
            .I(n14965));
    CascadeMux I__9775 (
            .O(N__43944),
            .I(N__43940));
    CascadeMux I__9774 (
            .O(N__43943),
            .I(N__43937));
    InMux I__9773 (
            .O(N__43940),
            .I(N__43933));
    InMux I__9772 (
            .O(N__43937),
            .I(N__43930));
    CascadeMux I__9771 (
            .O(N__43936),
            .I(N__43927));
    LocalMux I__9770 (
            .O(N__43933),
            .I(N__43921));
    LocalMux I__9769 (
            .O(N__43930),
            .I(N__43921));
    InMux I__9768 (
            .O(N__43927),
            .I(N__43916));
    InMux I__9767 (
            .O(N__43926),
            .I(N__43916));
    Odrv4 I__9766 (
            .O(N__43921),
            .I(trig_dds0));
    LocalMux I__9765 (
            .O(N__43916),
            .I(trig_dds0));
    CEMux I__9764 (
            .O(N__43911),
            .I(N__43907));
    CEMux I__9763 (
            .O(N__43910),
            .I(N__43904));
    LocalMux I__9762 (
            .O(N__43907),
            .I(N__43900));
    LocalMux I__9761 (
            .O(N__43904),
            .I(N__43897));
    CEMux I__9760 (
            .O(N__43903),
            .I(N__43894));
    Span4Mux_v I__9759 (
            .O(N__43900),
            .I(N__43891));
    Span4Mux_h I__9758 (
            .O(N__43897),
            .I(N__43888));
    LocalMux I__9757 (
            .O(N__43894),
            .I(N__43885));
    Span4Mux_h I__9756 (
            .O(N__43891),
            .I(N__43882));
    Span4Mux_h I__9755 (
            .O(N__43888),
            .I(N__43879));
    Span12Mux_h I__9754 (
            .O(N__43885),
            .I(N__43876));
    Odrv4 I__9753 (
            .O(N__43882),
            .I(\SIG_DDS.n12895 ));
    Odrv4 I__9752 (
            .O(N__43879),
            .I(\SIG_DDS.n12895 ));
    Odrv12 I__9751 (
            .O(N__43876),
            .I(\SIG_DDS.n12895 ));
    InMux I__9750 (
            .O(N__43869),
            .I(N__43866));
    LocalMux I__9749 (
            .O(N__43866),
            .I(N__43862));
    CascadeMux I__9748 (
            .O(N__43865),
            .I(N__43859));
    Span4Mux_v I__9747 (
            .O(N__43862),
            .I(N__43856));
    InMux I__9746 (
            .O(N__43859),
            .I(N__43853));
    Span4Mux_h I__9745 (
            .O(N__43856),
            .I(N__43850));
    LocalMux I__9744 (
            .O(N__43853),
            .I(data_idxvec_0));
    Odrv4 I__9743 (
            .O(N__43850),
            .I(data_idxvec_0));
    InMux I__9742 (
            .O(N__43845),
            .I(N__43841));
    InMux I__9741 (
            .O(N__43844),
            .I(N__43837));
    LocalMux I__9740 (
            .O(N__43841),
            .I(N__43834));
    InMux I__9739 (
            .O(N__43840),
            .I(N__43831));
    LocalMux I__9738 (
            .O(N__43837),
            .I(N__43828));
    Span4Mux_h I__9737 (
            .O(N__43834),
            .I(N__43825));
    LocalMux I__9736 (
            .O(N__43831),
            .I(data_cntvec_0));
    Odrv12 I__9735 (
            .O(N__43828),
            .I(data_cntvec_0));
    Odrv4 I__9734 (
            .O(N__43825),
            .I(data_cntvec_0));
    InMux I__9733 (
            .O(N__43818),
            .I(N__43815));
    LocalMux I__9732 (
            .O(N__43815),
            .I(N__43812));
    Span4Mux_v I__9731 (
            .O(N__43812),
            .I(N__43809));
    Span4Mux_h I__9730 (
            .O(N__43809),
            .I(N__43806));
    Odrv4 I__9729 (
            .O(N__43806),
            .I(buf_data_iac_8));
    CascadeMux I__9728 (
            .O(N__43803),
            .I(n26_cascade_));
    CascadeMux I__9727 (
            .O(N__43800),
            .I(n21261_cascade_));
    CascadeMux I__9726 (
            .O(N__43797),
            .I(n22563_cascade_));
    InMux I__9725 (
            .O(N__43794),
            .I(N__43791));
    LocalMux I__9724 (
            .O(N__43791),
            .I(N__43788));
    Odrv4 I__9723 (
            .O(N__43788),
            .I(n21257));
    CascadeMux I__9722 (
            .O(N__43785),
            .I(n22566_cascade_));
    InMux I__9721 (
            .O(N__43782),
            .I(N__43779));
    LocalMux I__9720 (
            .O(N__43779),
            .I(N__43776));
    Span4Mux_v I__9719 (
            .O(N__43776),
            .I(N__43773));
    Sp12to4 I__9718 (
            .O(N__43773),
            .I(N__43770));
    Span12Mux_h I__9717 (
            .O(N__43770),
            .I(N__43766));
    InMux I__9716 (
            .O(N__43769),
            .I(N__43763));
    Odrv12 I__9715 (
            .O(N__43766),
            .I(buf_adcdata_vdc_8));
    LocalMux I__9714 (
            .O(N__43763),
            .I(buf_adcdata_vdc_8));
    InMux I__9713 (
            .O(N__43758),
            .I(N__43754));
    CascadeMux I__9712 (
            .O(N__43757),
            .I(N__43751));
    LocalMux I__9711 (
            .O(N__43754),
            .I(N__43748));
    InMux I__9710 (
            .O(N__43751),
            .I(N__43745));
    Span4Mux_v I__9709 (
            .O(N__43748),
            .I(N__43742));
    LocalMux I__9708 (
            .O(N__43745),
            .I(N__43738));
    Span4Mux_h I__9707 (
            .O(N__43742),
            .I(N__43735));
    CascadeMux I__9706 (
            .O(N__43741),
            .I(N__43732));
    Span4Mux_v I__9705 (
            .O(N__43738),
            .I(N__43729));
    Span4Mux_h I__9704 (
            .O(N__43735),
            .I(N__43726));
    InMux I__9703 (
            .O(N__43732),
            .I(N__43723));
    Span4Mux_h I__9702 (
            .O(N__43729),
            .I(N__43720));
    Span4Mux_h I__9701 (
            .O(N__43726),
            .I(N__43717));
    LocalMux I__9700 (
            .O(N__43723),
            .I(buf_adcdata_vac_8));
    Odrv4 I__9699 (
            .O(N__43720),
            .I(buf_adcdata_vac_8));
    Odrv4 I__9698 (
            .O(N__43717),
            .I(buf_adcdata_vac_8));
    InMux I__9697 (
            .O(N__43710),
            .I(N__43707));
    LocalMux I__9696 (
            .O(N__43707),
            .I(N__43704));
    Span4Mux_h I__9695 (
            .O(N__43704),
            .I(N__43701));
    Span4Mux_v I__9694 (
            .O(N__43701),
            .I(N__43698));
    Span4Mux_h I__9693 (
            .O(N__43698),
            .I(N__43694));
    InMux I__9692 (
            .O(N__43697),
            .I(N__43691));
    Odrv4 I__9691 (
            .O(N__43694),
            .I(buf_readRTD_0));
    LocalMux I__9690 (
            .O(N__43691),
            .I(buf_readRTD_0));
    CascadeMux I__9689 (
            .O(N__43686),
            .I(n19_cascade_));
    InMux I__9688 (
            .O(N__43683),
            .I(N__43680));
    LocalMux I__9687 (
            .O(N__43680),
            .I(n21258));
    InMux I__9686 (
            .O(N__43677),
            .I(N__43673));
    InMux I__9685 (
            .O(N__43676),
            .I(N__43669));
    LocalMux I__9684 (
            .O(N__43673),
            .I(N__43666));
    InMux I__9683 (
            .O(N__43672),
            .I(N__43663));
    LocalMux I__9682 (
            .O(N__43669),
            .I(acadc_skipCount_0));
    Odrv12 I__9681 (
            .O(N__43666),
            .I(acadc_skipCount_0));
    LocalMux I__9680 (
            .O(N__43663),
            .I(acadc_skipCount_0));
    InMux I__9679 (
            .O(N__43656),
            .I(N__43653));
    LocalMux I__9678 (
            .O(N__43653),
            .I(N__43650));
    Span4Mux_h I__9677 (
            .O(N__43650),
            .I(N__43645));
    CascadeMux I__9676 (
            .O(N__43649),
            .I(N__43642));
    InMux I__9675 (
            .O(N__43648),
            .I(N__43639));
    Span4Mux_h I__9674 (
            .O(N__43645),
            .I(N__43636));
    InMux I__9673 (
            .O(N__43642),
            .I(N__43633));
    LocalMux I__9672 (
            .O(N__43639),
            .I(req_data_cnt_0));
    Odrv4 I__9671 (
            .O(N__43636),
            .I(req_data_cnt_0));
    LocalMux I__9670 (
            .O(N__43633),
            .I(req_data_cnt_0));
    InMux I__9669 (
            .O(N__43626),
            .I(N__43623));
    LocalMux I__9668 (
            .O(N__43623),
            .I(n21260));
    InMux I__9667 (
            .O(N__43620),
            .I(N__43617));
    LocalMux I__9666 (
            .O(N__43617),
            .I(N__43614));
    Span4Mux_h I__9665 (
            .O(N__43614),
            .I(N__43610));
    InMux I__9664 (
            .O(N__43613),
            .I(N__43607));
    Span4Mux_v I__9663 (
            .O(N__43610),
            .I(N__43602));
    LocalMux I__9662 (
            .O(N__43607),
            .I(N__43602));
    Span4Mux_h I__9661 (
            .O(N__43602),
            .I(N__43598));
    InMux I__9660 (
            .O(N__43601),
            .I(N__43595));
    Span4Mux_h I__9659 (
            .O(N__43598),
            .I(N__43592));
    LocalMux I__9658 (
            .O(N__43595),
            .I(buf_adcdata_iac_9));
    Odrv4 I__9657 (
            .O(N__43592),
            .I(buf_adcdata_iac_9));
    CascadeMux I__9656 (
            .O(N__43587),
            .I(N__43584));
    InMux I__9655 (
            .O(N__43584),
            .I(N__43581));
    LocalMux I__9654 (
            .O(N__43581),
            .I(N__43578));
    Odrv12 I__9653 (
            .O(N__43578),
            .I(n16_adj_1651));
    InMux I__9652 (
            .O(N__43575),
            .I(N__43572));
    LocalMux I__9651 (
            .O(N__43572),
            .I(N__43569));
    Span4Mux_v I__9650 (
            .O(N__43569),
            .I(N__43566));
    Span4Mux_h I__9649 (
            .O(N__43566),
            .I(N__43563));
    Odrv4 I__9648 (
            .O(N__43563),
            .I(n22431));
    CascadeMux I__9647 (
            .O(N__43560),
            .I(N__43556));
    InMux I__9646 (
            .O(N__43559),
            .I(N__43553));
    InMux I__9645 (
            .O(N__43556),
            .I(N__43550));
    LocalMux I__9644 (
            .O(N__43553),
            .I(N__43547));
    LocalMux I__9643 (
            .O(N__43550),
            .I(comm_buf_6_7));
    Odrv4 I__9642 (
            .O(N__43547),
            .I(comm_buf_6_7));
    InMux I__9641 (
            .O(N__43542),
            .I(N__43539));
    LocalMux I__9640 (
            .O(N__43539),
            .I(N__43535));
    InMux I__9639 (
            .O(N__43538),
            .I(N__43531));
    Span4Mux_h I__9638 (
            .O(N__43535),
            .I(N__43528));
    InMux I__9637 (
            .O(N__43534),
            .I(N__43525));
    LocalMux I__9636 (
            .O(N__43531),
            .I(acadc_skipCount_6));
    Odrv4 I__9635 (
            .O(N__43528),
            .I(acadc_skipCount_6));
    LocalMux I__9634 (
            .O(N__43525),
            .I(acadc_skipCount_6));
    InMux I__9633 (
            .O(N__43518),
            .I(N__43514));
    InMux I__9632 (
            .O(N__43517),
            .I(N__43510));
    LocalMux I__9631 (
            .O(N__43514),
            .I(N__43507));
    InMux I__9630 (
            .O(N__43513),
            .I(N__43504));
    LocalMux I__9629 (
            .O(N__43510),
            .I(req_data_cnt_6));
    Odrv12 I__9628 (
            .O(N__43507),
            .I(req_data_cnt_6));
    LocalMux I__9627 (
            .O(N__43504),
            .I(req_data_cnt_6));
    InMux I__9626 (
            .O(N__43497),
            .I(N__43494));
    LocalMux I__9625 (
            .O(N__43494),
            .I(N__43491));
    Odrv12 I__9624 (
            .O(N__43491),
            .I(n19_adj_1625));
    CascadeMux I__9623 (
            .O(N__43488),
            .I(N__43485));
    InMux I__9622 (
            .O(N__43485),
            .I(N__43482));
    LocalMux I__9621 (
            .O(N__43482),
            .I(N__43479));
    Span4Mux_v I__9620 (
            .O(N__43479),
            .I(N__43476));
    Span4Mux_h I__9619 (
            .O(N__43476),
            .I(N__43473));
    Sp12to4 I__9618 (
            .O(N__43473),
            .I(N__43469));
    InMux I__9617 (
            .O(N__43472),
            .I(N__43466));
    Odrv12 I__9616 (
            .O(N__43469),
            .I(buf_readRTD_6));
    LocalMux I__9615 (
            .O(N__43466),
            .I(buf_readRTD_6));
    InMux I__9614 (
            .O(N__43461),
            .I(N__43458));
    LocalMux I__9613 (
            .O(N__43458),
            .I(N__43454));
    CascadeMux I__9612 (
            .O(N__43457),
            .I(N__43451));
    Span4Mux_h I__9611 (
            .O(N__43454),
            .I(N__43448));
    InMux I__9610 (
            .O(N__43451),
            .I(N__43445));
    Span4Mux_h I__9609 (
            .O(N__43448),
            .I(N__43442));
    LocalMux I__9608 (
            .O(N__43445),
            .I(data_idxvec_6));
    Odrv4 I__9607 (
            .O(N__43442),
            .I(data_idxvec_6));
    InMux I__9606 (
            .O(N__43437),
            .I(N__43433));
    InMux I__9605 (
            .O(N__43436),
            .I(N__43429));
    LocalMux I__9604 (
            .O(N__43433),
            .I(N__43426));
    InMux I__9603 (
            .O(N__43432),
            .I(N__43423));
    LocalMux I__9602 (
            .O(N__43429),
            .I(N__43416));
    Span4Mux_h I__9601 (
            .O(N__43426),
            .I(N__43416));
    LocalMux I__9600 (
            .O(N__43423),
            .I(N__43416));
    Odrv4 I__9599 (
            .O(N__43416),
            .I(data_cntvec_6));
    CascadeMux I__9598 (
            .O(N__43413),
            .I(n26_adj_1626_cascade_));
    InMux I__9597 (
            .O(N__43410),
            .I(N__43407));
    LocalMux I__9596 (
            .O(N__43407),
            .I(n22515));
    InMux I__9595 (
            .O(N__43404),
            .I(N__43401));
    LocalMux I__9594 (
            .O(N__43401),
            .I(N__43398));
    Span4Mux_h I__9593 (
            .O(N__43398),
            .I(N__43395));
    Odrv4 I__9592 (
            .O(N__43395),
            .I(n16_adj_1624));
    InMux I__9591 (
            .O(N__43392),
            .I(N__43389));
    LocalMux I__9590 (
            .O(N__43389),
            .I(N__43385));
    CascadeMux I__9589 (
            .O(N__43388),
            .I(N__43382));
    Span4Mux_v I__9588 (
            .O(N__43385),
            .I(N__43379));
    InMux I__9587 (
            .O(N__43382),
            .I(N__43375));
    Sp12to4 I__9586 (
            .O(N__43379),
            .I(N__43372));
    InMux I__9585 (
            .O(N__43378),
            .I(N__43369));
    LocalMux I__9584 (
            .O(N__43375),
            .I(N__43364));
    Span12Mux_s10_h I__9583 (
            .O(N__43372),
            .I(N__43364));
    LocalMux I__9582 (
            .O(N__43369),
            .I(buf_adcdata_iac_14));
    Odrv12 I__9581 (
            .O(N__43364),
            .I(buf_adcdata_iac_14));
    InMux I__9580 (
            .O(N__43359),
            .I(N__43356));
    LocalMux I__9579 (
            .O(N__43356),
            .I(n22527));
    CascadeMux I__9578 (
            .O(N__43353),
            .I(n22530_cascade_));
    InMux I__9577 (
            .O(N__43350),
            .I(N__43347));
    LocalMux I__9576 (
            .O(N__43347),
            .I(n22518));
    CascadeMux I__9575 (
            .O(N__43344),
            .I(n30_adj_1627_cascade_));
    CascadeMux I__9574 (
            .O(N__43341),
            .I(n30_adj_1695_cascade_));
    CEMux I__9573 (
            .O(N__43338),
            .I(N__43333));
    CEMux I__9572 (
            .O(N__43337),
            .I(N__43330));
    CEMux I__9571 (
            .O(N__43336),
            .I(N__43327));
    LocalMux I__9570 (
            .O(N__43333),
            .I(N__43321));
    LocalMux I__9569 (
            .O(N__43330),
            .I(N__43318));
    LocalMux I__9568 (
            .O(N__43327),
            .I(N__43315));
    CEMux I__9567 (
            .O(N__43326),
            .I(N__43312));
    CEMux I__9566 (
            .O(N__43325),
            .I(N__43309));
    CEMux I__9565 (
            .O(N__43324),
            .I(N__43306));
    Span4Mux_h I__9564 (
            .O(N__43321),
            .I(N__43302));
    Span4Mux_v I__9563 (
            .O(N__43318),
            .I(N__43295));
    Span4Mux_h I__9562 (
            .O(N__43315),
            .I(N__43295));
    LocalMux I__9561 (
            .O(N__43312),
            .I(N__43295));
    LocalMux I__9560 (
            .O(N__43309),
            .I(N__43292));
    LocalMux I__9559 (
            .O(N__43306),
            .I(N__43289));
    InMux I__9558 (
            .O(N__43305),
            .I(N__43286));
    Odrv4 I__9557 (
            .O(N__43302),
            .I(n12184));
    Odrv4 I__9556 (
            .O(N__43295),
            .I(n12184));
    Odrv12 I__9555 (
            .O(N__43292),
            .I(n12184));
    Odrv4 I__9554 (
            .O(N__43289),
            .I(n12184));
    LocalMux I__9553 (
            .O(N__43286),
            .I(n12184));
    SRMux I__9552 (
            .O(N__43275),
            .I(N__43271));
    SRMux I__9551 (
            .O(N__43274),
            .I(N__43268));
    LocalMux I__9550 (
            .O(N__43271),
            .I(N__43265));
    LocalMux I__9549 (
            .O(N__43268),
            .I(N__43260));
    Span4Mux_h I__9548 (
            .O(N__43265),
            .I(N__43257));
    SRMux I__9547 (
            .O(N__43264),
            .I(N__43254));
    SRMux I__9546 (
            .O(N__43263),
            .I(N__43251));
    Span4Mux_v I__9545 (
            .O(N__43260),
            .I(N__43242));
    Span4Mux_h I__9544 (
            .O(N__43257),
            .I(N__43242));
    LocalMux I__9543 (
            .O(N__43254),
            .I(N__43242));
    LocalMux I__9542 (
            .O(N__43251),
            .I(N__43239));
    SRMux I__9541 (
            .O(N__43250),
            .I(N__43236));
    SRMux I__9540 (
            .O(N__43249),
            .I(N__43233));
    Span4Mux_v I__9539 (
            .O(N__43242),
            .I(N__43230));
    Sp12to4 I__9538 (
            .O(N__43239),
            .I(N__43225));
    LocalMux I__9537 (
            .O(N__43236),
            .I(N__43225));
    LocalMux I__9536 (
            .O(N__43233),
            .I(N__43222));
    Odrv4 I__9535 (
            .O(N__43230),
            .I(n14958));
    Odrv12 I__9534 (
            .O(N__43225),
            .I(n14958));
    Odrv12 I__9533 (
            .O(N__43222),
            .I(n14958));
    InMux I__9532 (
            .O(N__43215),
            .I(N__43212));
    LocalMux I__9531 (
            .O(N__43212),
            .I(N__43209));
    Odrv12 I__9530 (
            .O(N__43209),
            .I(n22539));
    InMux I__9529 (
            .O(N__43206),
            .I(N__43203));
    LocalMux I__9528 (
            .O(N__43203),
            .I(N__43200));
    Span4Mux_v I__9527 (
            .O(N__43200),
            .I(N__43195));
    InMux I__9526 (
            .O(N__43199),
            .I(N__43191));
    InMux I__9525 (
            .O(N__43198),
            .I(N__43188));
    Span4Mux_h I__9524 (
            .O(N__43195),
            .I(N__43185));
    InMux I__9523 (
            .O(N__43194),
            .I(N__43182));
    LocalMux I__9522 (
            .O(N__43191),
            .I(N__43179));
    LocalMux I__9521 (
            .O(N__43188),
            .I(N__43176));
    Span4Mux_h I__9520 (
            .O(N__43185),
            .I(N__43173));
    LocalMux I__9519 (
            .O(N__43182),
            .I(N__43170));
    Span4Mux_v I__9518 (
            .O(N__43179),
            .I(N__43165));
    Span4Mux_v I__9517 (
            .O(N__43176),
            .I(N__43165));
    Span4Mux_h I__9516 (
            .O(N__43173),
            .I(N__43162));
    Span4Mux_v I__9515 (
            .O(N__43170),
            .I(N__43157));
    Span4Mux_h I__9514 (
            .O(N__43165),
            .I(N__43157));
    Odrv4 I__9513 (
            .O(N__43162),
            .I(n14_adj_1541));
    Odrv4 I__9512 (
            .O(N__43157),
            .I(n14_adj_1541));
    InMux I__9511 (
            .O(N__43152),
            .I(N__43149));
    LocalMux I__9510 (
            .O(N__43149),
            .I(N__43146));
    Span4Mux_h I__9509 (
            .O(N__43146),
            .I(N__43143));
    Span4Mux_v I__9508 (
            .O(N__43143),
            .I(N__43140));
    Odrv4 I__9507 (
            .O(N__43140),
            .I(buf_data_iac_0));
    InMux I__9506 (
            .O(N__43137),
            .I(N__43134));
    LocalMux I__9505 (
            .O(N__43134),
            .I(N__43131));
    Span12Mux_v I__9504 (
            .O(N__43131),
            .I(N__43128));
    Odrv12 I__9503 (
            .O(N__43128),
            .I(n22_adj_1532));
    CascadeMux I__9502 (
            .O(N__43125),
            .I(N__43122));
    InMux I__9501 (
            .O(N__43122),
            .I(N__43119));
    LocalMux I__9500 (
            .O(N__43119),
            .I(N__43116));
    Odrv4 I__9499 (
            .O(N__43116),
            .I(n21586));
    CascadeMux I__9498 (
            .O(N__43113),
            .I(n21474_cascade_));
    CascadeMux I__9497 (
            .O(N__43110),
            .I(n12_adj_1596_cascade_));
    InMux I__9496 (
            .O(N__43107),
            .I(N__43103));
    CascadeMux I__9495 (
            .O(N__43106),
            .I(N__43100));
    LocalMux I__9494 (
            .O(N__43103),
            .I(N__43097));
    InMux I__9493 (
            .O(N__43100),
            .I(N__43094));
    Span12Mux_v I__9492 (
            .O(N__43097),
            .I(N__43091));
    LocalMux I__9491 (
            .O(N__43094),
            .I(data_idxvec_9));
    Odrv12 I__9490 (
            .O(N__43091),
            .I(data_idxvec_9));
    InMux I__9489 (
            .O(N__43086),
            .I(N__43082));
    InMux I__9488 (
            .O(N__43085),
            .I(N__43079));
    LocalMux I__9487 (
            .O(N__43082),
            .I(N__43075));
    LocalMux I__9486 (
            .O(N__43079),
            .I(N__43072));
    InMux I__9485 (
            .O(N__43078),
            .I(N__43069));
    Span4Mux_v I__9484 (
            .O(N__43075),
            .I(N__43064));
    Span4Mux_h I__9483 (
            .O(N__43072),
            .I(N__43064));
    LocalMux I__9482 (
            .O(N__43069),
            .I(data_cntvec_9));
    Odrv4 I__9481 (
            .O(N__43064),
            .I(data_cntvec_9));
    InMux I__9480 (
            .O(N__43059),
            .I(N__43056));
    LocalMux I__9479 (
            .O(N__43056),
            .I(N__43053));
    Odrv12 I__9478 (
            .O(N__43053),
            .I(buf_data_iac_17));
    CascadeMux I__9477 (
            .O(N__43050),
            .I(n26_adj_1694_cascade_));
    InMux I__9476 (
            .O(N__43047),
            .I(N__43044));
    LocalMux I__9475 (
            .O(N__43044),
            .I(N__43038));
    InMux I__9474 (
            .O(N__43043),
            .I(N__43035));
    InMux I__9473 (
            .O(N__43042),
            .I(N__43032));
    InMux I__9472 (
            .O(N__43041),
            .I(N__43029));
    Span4Mux_h I__9471 (
            .O(N__43038),
            .I(N__43025));
    LocalMux I__9470 (
            .O(N__43035),
            .I(N__43018));
    LocalMux I__9469 (
            .O(N__43032),
            .I(N__43018));
    LocalMux I__9468 (
            .O(N__43029),
            .I(N__43018));
    InMux I__9467 (
            .O(N__43028),
            .I(N__43015));
    Span4Mux_h I__9466 (
            .O(N__43025),
            .I(N__43012));
    Span4Mux_v I__9465 (
            .O(N__43018),
            .I(N__43009));
    LocalMux I__9464 (
            .O(N__43015),
            .I(eis_stop));
    Odrv4 I__9463 (
            .O(N__43012),
            .I(eis_stop));
    Odrv4 I__9462 (
            .O(N__43009),
            .I(eis_stop));
    InMux I__9461 (
            .O(N__43002),
            .I(N__42999));
    LocalMux I__9460 (
            .O(N__42999),
            .I(N__42996));
    Span4Mux_h I__9459 (
            .O(N__42996),
            .I(N__42991));
    InMux I__9458 (
            .O(N__42995),
            .I(N__42986));
    InMux I__9457 (
            .O(N__42994),
            .I(N__42986));
    Odrv4 I__9456 (
            .O(N__42991),
            .I(req_data_cnt_9));
    LocalMux I__9455 (
            .O(N__42986),
            .I(req_data_cnt_9));
    InMux I__9454 (
            .O(N__42981),
            .I(N__42978));
    LocalMux I__9453 (
            .O(N__42978),
            .I(N__42974));
    InMux I__9452 (
            .O(N__42977),
            .I(N__42970));
    Span12Mux_v I__9451 (
            .O(N__42974),
            .I(N__42967));
    InMux I__9450 (
            .O(N__42973),
            .I(N__42964));
    LocalMux I__9449 (
            .O(N__42970),
            .I(acadc_skipCount_9));
    Odrv12 I__9448 (
            .O(N__42967),
            .I(acadc_skipCount_9));
    LocalMux I__9447 (
            .O(N__42964),
            .I(acadc_skipCount_9));
    IoInMux I__9446 (
            .O(N__42957),
            .I(N__42954));
    LocalMux I__9445 (
            .O(N__42954),
            .I(N__42950));
    InMux I__9444 (
            .O(N__42953),
            .I(N__42947));
    Span12Mux_s0_v I__9443 (
            .O(N__42950),
            .I(N__42944));
    LocalMux I__9442 (
            .O(N__42947),
            .I(N__42941));
    Span12Mux_v I__9441 (
            .O(N__42944),
            .I(N__42938));
    Span4Mux_v I__9440 (
            .O(N__42941),
            .I(N__42934));
    Span12Mux_h I__9439 (
            .O(N__42938),
            .I(N__42931));
    InMux I__9438 (
            .O(N__42937),
            .I(N__42928));
    Span4Mux_h I__9437 (
            .O(N__42934),
            .I(N__42925));
    Odrv12 I__9436 (
            .O(N__42931),
            .I(DDS_RNG_0));
    LocalMux I__9435 (
            .O(N__42928),
            .I(DDS_RNG_0));
    Odrv4 I__9434 (
            .O(N__42925),
            .I(DDS_RNG_0));
    CascadeMux I__9433 (
            .O(N__42918),
            .I(n22617_cascade_));
    CascadeMux I__9432 (
            .O(N__42915),
            .I(n22620_cascade_));
    InMux I__9431 (
            .O(N__42912),
            .I(N__42909));
    LocalMux I__9430 (
            .O(N__42909),
            .I(n21360));
    InMux I__9429 (
            .O(N__42906),
            .I(N__42903));
    LocalMux I__9428 (
            .O(N__42903),
            .I(N__42900));
    Span4Mux_v I__9427 (
            .O(N__42900),
            .I(N__42897));
    Sp12to4 I__9426 (
            .O(N__42897),
            .I(N__42894));
    Odrv12 I__9425 (
            .O(N__42894),
            .I(n22410));
    CascadeMux I__9424 (
            .O(N__42891),
            .I(n21361_cascade_));
    SRMux I__9423 (
            .O(N__42888),
            .I(N__42884));
    SRMux I__9422 (
            .O(N__42887),
            .I(N__42881));
    LocalMux I__9421 (
            .O(N__42884),
            .I(N__42877));
    LocalMux I__9420 (
            .O(N__42881),
            .I(N__42874));
    SRMux I__9419 (
            .O(N__42880),
            .I(N__42871));
    Span4Mux_v I__9418 (
            .O(N__42877),
            .I(N__42866));
    Span4Mux_v I__9417 (
            .O(N__42874),
            .I(N__42866));
    LocalMux I__9416 (
            .O(N__42871),
            .I(N__42863));
    Span4Mux_v I__9415 (
            .O(N__42866),
            .I(N__42860));
    Span4Mux_v I__9414 (
            .O(N__42863),
            .I(N__42857));
    Odrv4 I__9413 (
            .O(N__42860),
            .I(\comm_spi.data_tx_7__N_814 ));
    Odrv4 I__9412 (
            .O(N__42857),
            .I(\comm_spi.data_tx_7__N_814 ));
    CascadeMux I__9411 (
            .O(N__42852),
            .I(N__42848));
    InMux I__9410 (
            .O(N__42851),
            .I(N__42840));
    InMux I__9409 (
            .O(N__42848),
            .I(N__42840));
    InMux I__9408 (
            .O(N__42847),
            .I(N__42840));
    LocalMux I__9407 (
            .O(N__42840),
            .I(comm_tx_buf_7));
    SRMux I__9406 (
            .O(N__42837),
            .I(N__42833));
    SRMux I__9405 (
            .O(N__42836),
            .I(N__42830));
    LocalMux I__9404 (
            .O(N__42833),
            .I(N__42826));
    LocalMux I__9403 (
            .O(N__42830),
            .I(N__42823));
    SRMux I__9402 (
            .O(N__42829),
            .I(N__42820));
    Span4Mux_v I__9401 (
            .O(N__42826),
            .I(N__42815));
    Span4Mux_h I__9400 (
            .O(N__42823),
            .I(N__42815));
    LocalMux I__9399 (
            .O(N__42820),
            .I(N__42812));
    Span4Mux_v I__9398 (
            .O(N__42815),
            .I(N__42809));
    Span4Mux_v I__9397 (
            .O(N__42812),
            .I(N__42806));
    Odrv4 I__9396 (
            .O(N__42809),
            .I(\comm_spi.data_tx_7__N_806 ));
    Odrv4 I__9395 (
            .O(N__42806),
            .I(\comm_spi.data_tx_7__N_806 ));
    InMux I__9394 (
            .O(N__42801),
            .I(N__42798));
    LocalMux I__9393 (
            .O(N__42798),
            .I(N__42792));
    CascadeMux I__9392 (
            .O(N__42797),
            .I(N__42788));
    CascadeMux I__9391 (
            .O(N__42796),
            .I(N__42785));
    CascadeMux I__9390 (
            .O(N__42795),
            .I(N__42782));
    Span4Mux_v I__9389 (
            .O(N__42792),
            .I(N__42775));
    InMux I__9388 (
            .O(N__42791),
            .I(N__42772));
    InMux I__9387 (
            .O(N__42788),
            .I(N__42757));
    InMux I__9386 (
            .O(N__42785),
            .I(N__42757));
    InMux I__9385 (
            .O(N__42782),
            .I(N__42757));
    InMux I__9384 (
            .O(N__42781),
            .I(N__42757));
    InMux I__9383 (
            .O(N__42780),
            .I(N__42757));
    InMux I__9382 (
            .O(N__42779),
            .I(N__42757));
    InMux I__9381 (
            .O(N__42778),
            .I(N__42757));
    Odrv4 I__9380 (
            .O(N__42775),
            .I(\comm_spi.bit_cnt_3 ));
    LocalMux I__9379 (
            .O(N__42772),
            .I(\comm_spi.bit_cnt_3 ));
    LocalMux I__9378 (
            .O(N__42757),
            .I(\comm_spi.bit_cnt_3 ));
    InMux I__9377 (
            .O(N__42750),
            .I(N__42747));
    LocalMux I__9376 (
            .O(N__42747),
            .I(N__42737));
    InMux I__9375 (
            .O(N__42746),
            .I(N__42722));
    InMux I__9374 (
            .O(N__42745),
            .I(N__42722));
    InMux I__9373 (
            .O(N__42744),
            .I(N__42722));
    InMux I__9372 (
            .O(N__42743),
            .I(N__42722));
    InMux I__9371 (
            .O(N__42742),
            .I(N__42722));
    InMux I__9370 (
            .O(N__42741),
            .I(N__42722));
    InMux I__9369 (
            .O(N__42740),
            .I(N__42722));
    Odrv4 I__9368 (
            .O(N__42737),
            .I(\comm_spi.n17254 ));
    LocalMux I__9367 (
            .O(N__42722),
            .I(\comm_spi.n17254 ));
    CascadeMux I__9366 (
            .O(N__42717),
            .I(n22551_cascade_));
    CascadeMux I__9365 (
            .O(N__42714),
            .I(N__42711));
    InMux I__9364 (
            .O(N__42711),
            .I(N__42704));
    InMux I__9363 (
            .O(N__42710),
            .I(N__42701));
    InMux I__9362 (
            .O(N__42709),
            .I(N__42698));
    InMux I__9361 (
            .O(N__42708),
            .I(N__42695));
    CascadeMux I__9360 (
            .O(N__42707),
            .I(N__42692));
    LocalMux I__9359 (
            .O(N__42704),
            .I(N__42689));
    LocalMux I__9358 (
            .O(N__42701),
            .I(N__42686));
    LocalMux I__9357 (
            .O(N__42698),
            .I(N__42683));
    LocalMux I__9356 (
            .O(N__42695),
            .I(N__42680));
    InMux I__9355 (
            .O(N__42692),
            .I(N__42677));
    Span4Mux_h I__9354 (
            .O(N__42689),
            .I(N__42672));
    Span4Mux_h I__9353 (
            .O(N__42686),
            .I(N__42672));
    Span4Mux_v I__9352 (
            .O(N__42683),
            .I(N__42669));
    Span4Mux_h I__9351 (
            .O(N__42680),
            .I(N__42666));
    LocalMux I__9350 (
            .O(N__42677),
            .I(N__42663));
    Span4Mux_h I__9349 (
            .O(N__42672),
            .I(N__42660));
    Span4Mux_h I__9348 (
            .O(N__42669),
            .I(N__42655));
    Span4Mux_v I__9347 (
            .O(N__42666),
            .I(N__42655));
    Odrv4 I__9346 (
            .O(N__42663),
            .I(comm_buf_1_4));
    Odrv4 I__9345 (
            .O(N__42660),
            .I(comm_buf_1_4));
    Odrv4 I__9344 (
            .O(N__42655),
            .I(comm_buf_1_4));
    CascadeMux I__9343 (
            .O(N__42648),
            .I(n4_adj_1582_cascade_));
    CascadeMux I__9342 (
            .O(N__42645),
            .I(n21285_cascade_));
    InMux I__9341 (
            .O(N__42642),
            .I(N__42639));
    LocalMux I__9340 (
            .O(N__42639),
            .I(n22554));
    CEMux I__9339 (
            .O(N__42636),
            .I(N__42632));
    CEMux I__9338 (
            .O(N__42635),
            .I(N__42627));
    LocalMux I__9337 (
            .O(N__42632),
            .I(N__42624));
    CEMux I__9336 (
            .O(N__42631),
            .I(N__42621));
    CEMux I__9335 (
            .O(N__42630),
            .I(N__42618));
    LocalMux I__9334 (
            .O(N__42627),
            .I(N__42615));
    Span4Mux_v I__9333 (
            .O(N__42624),
            .I(N__42612));
    LocalMux I__9332 (
            .O(N__42621),
            .I(N__42609));
    LocalMux I__9331 (
            .O(N__42618),
            .I(N__42606));
    Span4Mux_h I__9330 (
            .O(N__42615),
            .I(N__42601));
    Span4Mux_h I__9329 (
            .O(N__42612),
            .I(N__42601));
    Span4Mux_h I__9328 (
            .O(N__42609),
            .I(N__42598));
    Span4Mux_h I__9327 (
            .O(N__42606),
            .I(N__42595));
    Odrv4 I__9326 (
            .O(N__42601),
            .I(n11910));
    Odrv4 I__9325 (
            .O(N__42598),
            .I(n11910));
    Odrv4 I__9324 (
            .O(N__42595),
            .I(n11910));
    InMux I__9323 (
            .O(N__42588),
            .I(N__42585));
    LocalMux I__9322 (
            .O(N__42585),
            .I(N__42582));
    Span4Mux_v I__9321 (
            .O(N__42582),
            .I(N__42579));
    Span4Mux_v I__9320 (
            .O(N__42579),
            .I(N__42576));
    Span4Mux_h I__9319 (
            .O(N__42576),
            .I(N__42573));
    Odrv4 I__9318 (
            .O(N__42573),
            .I(buf_data_iac_10));
    InMux I__9317 (
            .O(N__42570),
            .I(N__42567));
    LocalMux I__9316 (
            .O(N__42567),
            .I(N__42564));
    Span4Mux_v I__9315 (
            .O(N__42564),
            .I(N__42561));
    Span4Mux_h I__9314 (
            .O(N__42561),
            .I(N__42558));
    Odrv4 I__9313 (
            .O(N__42558),
            .I(n21385));
    InMux I__9312 (
            .O(N__42555),
            .I(N__42551));
    CascadeMux I__9311 (
            .O(N__42554),
            .I(N__42547));
    LocalMux I__9310 (
            .O(N__42551),
            .I(N__42544));
    CascadeMux I__9309 (
            .O(N__42550),
            .I(N__42539));
    InMux I__9308 (
            .O(N__42547),
            .I(N__42536));
    Span4Mux_h I__9307 (
            .O(N__42544),
            .I(N__42532));
    InMux I__9306 (
            .O(N__42543),
            .I(N__42527));
    InMux I__9305 (
            .O(N__42542),
            .I(N__42527));
    InMux I__9304 (
            .O(N__42539),
            .I(N__42524));
    LocalMux I__9303 (
            .O(N__42536),
            .I(N__42521));
    InMux I__9302 (
            .O(N__42535),
            .I(N__42518));
    Sp12to4 I__9301 (
            .O(N__42532),
            .I(N__42512));
    LocalMux I__9300 (
            .O(N__42527),
            .I(N__42512));
    LocalMux I__9299 (
            .O(N__42524),
            .I(N__42509));
    Span4Mux_v I__9298 (
            .O(N__42521),
            .I(N__42504));
    LocalMux I__9297 (
            .O(N__42518),
            .I(N__42504));
    InMux I__9296 (
            .O(N__42517),
            .I(N__42501));
    Span12Mux_v I__9295 (
            .O(N__42512),
            .I(N__42498));
    Span4Mux_v I__9294 (
            .O(N__42509),
            .I(N__42495));
    Span4Mux_h I__9293 (
            .O(N__42504),
            .I(N__42490));
    LocalMux I__9292 (
            .O(N__42501),
            .I(N__42490));
    Odrv12 I__9291 (
            .O(N__42498),
            .I(comm_buf_0_7));
    Odrv4 I__9290 (
            .O(N__42495),
            .I(comm_buf_0_7));
    Odrv4 I__9289 (
            .O(N__42490),
            .I(comm_buf_0_7));
    InMux I__9288 (
            .O(N__42483),
            .I(N__42480));
    LocalMux I__9287 (
            .O(N__42480),
            .I(N__42477));
    Odrv4 I__9286 (
            .O(N__42477),
            .I(n21276));
    CascadeMux I__9285 (
            .O(N__42474),
            .I(n22542_cascade_));
    InMux I__9284 (
            .O(N__42471),
            .I(N__42468));
    LocalMux I__9283 (
            .O(N__42468),
            .I(N__42465));
    Odrv4 I__9282 (
            .O(N__42465),
            .I(n4_adj_1580));
    IoInMux I__9281 (
            .O(N__42462),
            .I(N__42459));
    LocalMux I__9280 (
            .O(N__42459),
            .I(N__42456));
    IoSpan4Mux I__9279 (
            .O(N__42456),
            .I(N__42453));
    Span4Mux_s0_h I__9278 (
            .O(N__42453),
            .I(N__42450));
    Sp12to4 I__9277 (
            .O(N__42450),
            .I(N__42447));
    Span12Mux_h I__9276 (
            .O(N__42447),
            .I(N__42443));
    InMux I__9275 (
            .O(N__42446),
            .I(N__42440));
    Odrv12 I__9274 (
            .O(N__42443),
            .I(VDC_SCLK));
    LocalMux I__9273 (
            .O(N__42440),
            .I(VDC_SCLK));
    IoInMux I__9272 (
            .O(N__42435),
            .I(N__42431));
    ClkMux I__9271 (
            .O(N__42434),
            .I(N__42426));
    LocalMux I__9270 (
            .O(N__42431),
            .I(N__42421));
    ClkMux I__9269 (
            .O(N__42430),
            .I(N__42418));
    ClkMux I__9268 (
            .O(N__42429),
            .I(N__42415));
    LocalMux I__9267 (
            .O(N__42426),
            .I(N__42406));
    ClkMux I__9266 (
            .O(N__42425),
            .I(N__42403));
    ClkMux I__9265 (
            .O(N__42424),
            .I(N__42400));
    Span4Mux_s1_h I__9264 (
            .O(N__42421),
            .I(N__42395));
    LocalMux I__9263 (
            .O(N__42418),
            .I(N__42391));
    LocalMux I__9262 (
            .O(N__42415),
            .I(N__42388));
    ClkMux I__9261 (
            .O(N__42414),
            .I(N__42385));
    ClkMux I__9260 (
            .O(N__42413),
            .I(N__42380));
    ClkMux I__9259 (
            .O(N__42412),
            .I(N__42377));
    ClkMux I__9258 (
            .O(N__42411),
            .I(N__42374));
    ClkMux I__9257 (
            .O(N__42410),
            .I(N__42369));
    ClkMux I__9256 (
            .O(N__42409),
            .I(N__42366));
    Span4Mux_h I__9255 (
            .O(N__42406),
            .I(N__42357));
    LocalMux I__9254 (
            .O(N__42403),
            .I(N__42357));
    LocalMux I__9253 (
            .O(N__42400),
            .I(N__42354));
    ClkMux I__9252 (
            .O(N__42399),
            .I(N__42351));
    ClkMux I__9251 (
            .O(N__42398),
            .I(N__42348));
    Span4Mux_h I__9250 (
            .O(N__42395),
            .I(N__42345));
    ClkMux I__9249 (
            .O(N__42394),
            .I(N__42342));
    Span4Mux_v I__9248 (
            .O(N__42391),
            .I(N__42335));
    Span4Mux_v I__9247 (
            .O(N__42388),
            .I(N__42335));
    LocalMux I__9246 (
            .O(N__42385),
            .I(N__42335));
    ClkMux I__9245 (
            .O(N__42384),
            .I(N__42331));
    ClkMux I__9244 (
            .O(N__42383),
            .I(N__42328));
    LocalMux I__9243 (
            .O(N__42380),
            .I(N__42325));
    LocalMux I__9242 (
            .O(N__42377),
            .I(N__42320));
    LocalMux I__9241 (
            .O(N__42374),
            .I(N__42320));
    ClkMux I__9240 (
            .O(N__42373),
            .I(N__42317));
    ClkMux I__9239 (
            .O(N__42372),
            .I(N__42314));
    LocalMux I__9238 (
            .O(N__42369),
            .I(N__42309));
    LocalMux I__9237 (
            .O(N__42366),
            .I(N__42309));
    ClkMux I__9236 (
            .O(N__42365),
            .I(N__42306));
    ClkMux I__9235 (
            .O(N__42364),
            .I(N__42302));
    ClkMux I__9234 (
            .O(N__42363),
            .I(N__42298));
    ClkMux I__9233 (
            .O(N__42362),
            .I(N__42295));
    Span4Mux_v I__9232 (
            .O(N__42357),
            .I(N__42286));
    Span4Mux_h I__9231 (
            .O(N__42354),
            .I(N__42286));
    LocalMux I__9230 (
            .O(N__42351),
            .I(N__42286));
    LocalMux I__9229 (
            .O(N__42348),
            .I(N__42286));
    Span4Mux_h I__9228 (
            .O(N__42345),
            .I(N__42279));
    LocalMux I__9227 (
            .O(N__42342),
            .I(N__42279));
    Span4Mux_h I__9226 (
            .O(N__42335),
            .I(N__42279));
    ClkMux I__9225 (
            .O(N__42334),
            .I(N__42276));
    LocalMux I__9224 (
            .O(N__42331),
            .I(N__42269));
    LocalMux I__9223 (
            .O(N__42328),
            .I(N__42269));
    Span4Mux_v I__9222 (
            .O(N__42325),
            .I(N__42269));
    Span4Mux_v I__9221 (
            .O(N__42320),
            .I(N__42264));
    LocalMux I__9220 (
            .O(N__42317),
            .I(N__42264));
    LocalMux I__9219 (
            .O(N__42314),
            .I(N__42261));
    Span4Mux_v I__9218 (
            .O(N__42309),
            .I(N__42256));
    LocalMux I__9217 (
            .O(N__42306),
            .I(N__42256));
    ClkMux I__9216 (
            .O(N__42305),
            .I(N__42253));
    LocalMux I__9215 (
            .O(N__42302),
            .I(N__42250));
    ClkMux I__9214 (
            .O(N__42301),
            .I(N__42247));
    LocalMux I__9213 (
            .O(N__42298),
            .I(N__42244));
    LocalMux I__9212 (
            .O(N__42295),
            .I(N__42235));
    Span4Mux_v I__9211 (
            .O(N__42286),
            .I(N__42235));
    Span4Mux_h I__9210 (
            .O(N__42279),
            .I(N__42235));
    LocalMux I__9209 (
            .O(N__42276),
            .I(N__42235));
    Span4Mux_v I__9208 (
            .O(N__42269),
            .I(N__42230));
    Span4Mux_h I__9207 (
            .O(N__42264),
            .I(N__42230));
    Span4Mux_v I__9206 (
            .O(N__42261),
            .I(N__42227));
    Span4Mux_h I__9205 (
            .O(N__42256),
            .I(N__42222));
    LocalMux I__9204 (
            .O(N__42253),
            .I(N__42222));
    Span4Mux_h I__9203 (
            .O(N__42250),
            .I(N__42218));
    LocalMux I__9202 (
            .O(N__42247),
            .I(N__42215));
    Span4Mux_v I__9201 (
            .O(N__42244),
            .I(N__42212));
    Span4Mux_h I__9200 (
            .O(N__42235),
            .I(N__42209));
    Span4Mux_h I__9199 (
            .O(N__42230),
            .I(N__42204));
    Span4Mux_v I__9198 (
            .O(N__42227),
            .I(N__42204));
    Span4Mux_h I__9197 (
            .O(N__42222),
            .I(N__42201));
    ClkMux I__9196 (
            .O(N__42221),
            .I(N__42198));
    Odrv4 I__9195 (
            .O(N__42218),
            .I(VDC_CLK));
    Odrv12 I__9194 (
            .O(N__42215),
            .I(VDC_CLK));
    Odrv4 I__9193 (
            .O(N__42212),
            .I(VDC_CLK));
    Odrv4 I__9192 (
            .O(N__42209),
            .I(VDC_CLK));
    Odrv4 I__9191 (
            .O(N__42204),
            .I(VDC_CLK));
    Odrv4 I__9190 (
            .O(N__42201),
            .I(VDC_CLK));
    LocalMux I__9189 (
            .O(N__42198),
            .I(VDC_CLK));
    InMux I__9188 (
            .O(N__42183),
            .I(N__42180));
    LocalMux I__9187 (
            .O(N__42180),
            .I(N__42177));
    Span4Mux_h I__9186 (
            .O(N__42177),
            .I(N__42174));
    Span4Mux_h I__9185 (
            .O(N__42174),
            .I(N__42171));
    Odrv4 I__9184 (
            .O(N__42171),
            .I(buf_data_iac_20));
    InMux I__9183 (
            .O(N__42168),
            .I(N__42165));
    LocalMux I__9182 (
            .O(N__42165),
            .I(N__42162));
    Span4Mux_h I__9181 (
            .O(N__42162),
            .I(N__42159));
    Span4Mux_v I__9180 (
            .O(N__42159),
            .I(N__42156));
    Odrv4 I__9179 (
            .O(N__42156),
            .I(n21557));
    SRMux I__9178 (
            .O(N__42153),
            .I(N__42148));
    SRMux I__9177 (
            .O(N__42152),
            .I(N__42144));
    SRMux I__9176 (
            .O(N__42151),
            .I(N__42140));
    LocalMux I__9175 (
            .O(N__42148),
            .I(N__42137));
    SRMux I__9174 (
            .O(N__42147),
            .I(N__42134));
    LocalMux I__9173 (
            .O(N__42144),
            .I(N__42131));
    SRMux I__9172 (
            .O(N__42143),
            .I(N__42128));
    LocalMux I__9171 (
            .O(N__42140),
            .I(N__42125));
    Span4Mux_v I__9170 (
            .O(N__42137),
            .I(N__42120));
    LocalMux I__9169 (
            .O(N__42134),
            .I(N__42120));
    Span4Mux_h I__9168 (
            .O(N__42131),
            .I(N__42115));
    LocalMux I__9167 (
            .O(N__42128),
            .I(N__42115));
    Span4Mux_h I__9166 (
            .O(N__42125),
            .I(N__42112));
    Span4Mux_h I__9165 (
            .O(N__42120),
            .I(N__42109));
    Odrv4 I__9164 (
            .O(N__42115),
            .I(flagcntwd));
    Odrv4 I__9163 (
            .O(N__42112),
            .I(flagcntwd));
    Odrv4 I__9162 (
            .O(N__42109),
            .I(flagcntwd));
    CascadeMux I__9161 (
            .O(N__42102),
            .I(n21187_cascade_));
    CEMux I__9160 (
            .O(N__42099),
            .I(N__42096));
    LocalMux I__9159 (
            .O(N__42096),
            .I(n11605));
    SRMux I__9158 (
            .O(N__42093),
            .I(N__42090));
    LocalMux I__9157 (
            .O(N__42090),
            .I(N__42087));
    Span4Mux_h I__9156 (
            .O(N__42087),
            .I(N__42084));
    Span4Mux_h I__9155 (
            .O(N__42084),
            .I(N__42080));
    SRMux I__9154 (
            .O(N__42083),
            .I(N__42077));
    Odrv4 I__9153 (
            .O(N__42080),
            .I(n20578));
    LocalMux I__9152 (
            .O(N__42077),
            .I(n20578));
    CascadeMux I__9151 (
            .O(N__42072),
            .I(n11576_cascade_));
    CEMux I__9150 (
            .O(N__42069),
            .I(N__42066));
    LocalMux I__9149 (
            .O(N__42066),
            .I(N__42063));
    Span4Mux_h I__9148 (
            .O(N__42063),
            .I(N__42060));
    Span4Mux_h I__9147 (
            .O(N__42060),
            .I(N__42057));
    Odrv4 I__9146 (
            .O(N__42057),
            .I(n12148));
    InMux I__9145 (
            .O(N__42054),
            .I(N__42051));
    LocalMux I__9144 (
            .O(N__42051),
            .I(N__42047));
    InMux I__9143 (
            .O(N__42050),
            .I(N__42043));
    Span4Mux_v I__9142 (
            .O(N__42047),
            .I(N__42040));
    CascadeMux I__9141 (
            .O(N__42046),
            .I(N__42037));
    LocalMux I__9140 (
            .O(N__42043),
            .I(N__42032));
    Span4Mux_h I__9139 (
            .O(N__42040),
            .I(N__42032));
    InMux I__9138 (
            .O(N__42037),
            .I(N__42029));
    Span4Mux_h I__9137 (
            .O(N__42032),
            .I(N__42026));
    LocalMux I__9136 (
            .O(N__42029),
            .I(buf_adcdata_iac_15));
    Odrv4 I__9135 (
            .O(N__42026),
            .I(buf_adcdata_iac_15));
    InMux I__9134 (
            .O(N__42021),
            .I(N__42018));
    LocalMux I__9133 (
            .O(N__42018),
            .I(N__42015));
    Span4Mux_h I__9132 (
            .O(N__42015),
            .I(N__42012));
    Odrv4 I__9131 (
            .O(N__42012),
            .I(n16_adj_1620));
    CascadeMux I__9130 (
            .O(N__42009),
            .I(N__42005));
    InMux I__9129 (
            .O(N__42008),
            .I(N__42002));
    InMux I__9128 (
            .O(N__42005),
            .I(N__41998));
    LocalMux I__9127 (
            .O(N__42002),
            .I(N__41995));
    InMux I__9126 (
            .O(N__42001),
            .I(N__41992));
    LocalMux I__9125 (
            .O(N__41998),
            .I(N__41985));
    Span4Mux_h I__9124 (
            .O(N__41995),
            .I(N__41982));
    LocalMux I__9123 (
            .O(N__41992),
            .I(N__41979));
    InMux I__9122 (
            .O(N__41991),
            .I(N__41974));
    InMux I__9121 (
            .O(N__41990),
            .I(N__41974));
    InMux I__9120 (
            .O(N__41989),
            .I(N__41969));
    InMux I__9119 (
            .O(N__41988),
            .I(N__41969));
    Span4Mux_h I__9118 (
            .O(N__41985),
            .I(N__41966));
    Sp12to4 I__9117 (
            .O(N__41982),
            .I(N__41963));
    Sp12to4 I__9116 (
            .O(N__41979),
            .I(N__41960));
    LocalMux I__9115 (
            .O(N__41974),
            .I(n12144));
    LocalMux I__9114 (
            .O(N__41969),
            .I(n12144));
    Odrv4 I__9113 (
            .O(N__41966),
            .I(n12144));
    Odrv12 I__9112 (
            .O(N__41963),
            .I(n12144));
    Odrv12 I__9111 (
            .O(N__41960),
            .I(n12144));
    IoInMux I__9110 (
            .O(N__41949),
            .I(N__41946));
    LocalMux I__9109 (
            .O(N__41946),
            .I(N__41943));
    Span12Mux_s0_v I__9108 (
            .O(N__41943),
            .I(N__41940));
    Span12Mux_h I__9107 (
            .O(N__41940),
            .I(N__41937));
    Odrv12 I__9106 (
            .O(N__41937),
            .I(DDS_CS));
    CEMux I__9105 (
            .O(N__41934),
            .I(N__41931));
    LocalMux I__9104 (
            .O(N__41931),
            .I(N__41928));
    Span4Mux_h I__9103 (
            .O(N__41928),
            .I(N__41925));
    Odrv4 I__9102 (
            .O(N__41925),
            .I(\SIG_DDS.n9_adj_1434 ));
    CascadeMux I__9101 (
            .O(N__41922),
            .I(N__41919));
    InMux I__9100 (
            .O(N__41919),
            .I(N__41916));
    LocalMux I__9099 (
            .O(N__41916),
            .I(N__41912));
    InMux I__9098 (
            .O(N__41915),
            .I(N__41909));
    Odrv4 I__9097 (
            .O(N__41912),
            .I(n8_adj_1556));
    LocalMux I__9096 (
            .O(N__41909),
            .I(n8_adj_1556));
    InMux I__9095 (
            .O(N__41904),
            .I(N__41901));
    LocalMux I__9094 (
            .O(N__41901),
            .I(N__41897));
    InMux I__9093 (
            .O(N__41900),
            .I(N__41894));
    Span4Mux_v I__9092 (
            .O(N__41897),
            .I(N__41891));
    LocalMux I__9091 (
            .O(N__41894),
            .I(n7_adj_1555));
    Odrv4 I__9090 (
            .O(N__41891),
            .I(n7_adj_1555));
    CascadeMux I__9089 (
            .O(N__41886),
            .I(N__41883));
    CascadeBuf I__9088 (
            .O(N__41883),
            .I(N__41880));
    CascadeMux I__9087 (
            .O(N__41880),
            .I(N__41877));
    CascadeBuf I__9086 (
            .O(N__41877),
            .I(N__41874));
    CascadeMux I__9085 (
            .O(N__41874),
            .I(N__41871));
    CascadeBuf I__9084 (
            .O(N__41871),
            .I(N__41868));
    CascadeMux I__9083 (
            .O(N__41868),
            .I(N__41865));
    CascadeBuf I__9082 (
            .O(N__41865),
            .I(N__41862));
    CascadeMux I__9081 (
            .O(N__41862),
            .I(N__41859));
    CascadeBuf I__9080 (
            .O(N__41859),
            .I(N__41856));
    CascadeMux I__9079 (
            .O(N__41856),
            .I(N__41853));
    CascadeBuf I__9078 (
            .O(N__41853),
            .I(N__41850));
    CascadeMux I__9077 (
            .O(N__41850),
            .I(N__41847));
    CascadeBuf I__9076 (
            .O(N__41847),
            .I(N__41844));
    CascadeMux I__9075 (
            .O(N__41844),
            .I(N__41840));
    CascadeMux I__9074 (
            .O(N__41843),
            .I(N__41837));
    CascadeBuf I__9073 (
            .O(N__41840),
            .I(N__41834));
    CascadeBuf I__9072 (
            .O(N__41837),
            .I(N__41831));
    CascadeMux I__9071 (
            .O(N__41834),
            .I(N__41828));
    CascadeMux I__9070 (
            .O(N__41831),
            .I(N__41825));
    CascadeBuf I__9069 (
            .O(N__41828),
            .I(N__41822));
    InMux I__9068 (
            .O(N__41825),
            .I(N__41819));
    CascadeMux I__9067 (
            .O(N__41822),
            .I(N__41816));
    LocalMux I__9066 (
            .O(N__41819),
            .I(N__41813));
    InMux I__9065 (
            .O(N__41816),
            .I(N__41810));
    Span12Mux_h I__9064 (
            .O(N__41813),
            .I(N__41807));
    LocalMux I__9063 (
            .O(N__41810),
            .I(N__41804));
    Odrv12 I__9062 (
            .O(N__41807),
            .I(data_index_9_N_212_9));
    Odrv12 I__9061 (
            .O(N__41804),
            .I(data_index_9_N_212_9));
    InMux I__9060 (
            .O(N__41799),
            .I(N__41795));
    InMux I__9059 (
            .O(N__41798),
            .I(N__41792));
    LocalMux I__9058 (
            .O(N__41795),
            .I(\comm_spi.n14818 ));
    LocalMux I__9057 (
            .O(N__41792),
            .I(\comm_spi.n14818 ));
    InMux I__9056 (
            .O(N__41787),
            .I(N__41784));
    LocalMux I__9055 (
            .O(N__41784),
            .I(N__41780));
    InMux I__9054 (
            .O(N__41783),
            .I(N__41777));
    Span4Mux_v I__9053 (
            .O(N__41780),
            .I(N__41772));
    LocalMux I__9052 (
            .O(N__41777),
            .I(N__41772));
    Odrv4 I__9051 (
            .O(N__41772),
            .I(\comm_spi.n14819 ));
    InMux I__9050 (
            .O(N__41769),
            .I(N__41766));
    LocalMux I__9049 (
            .O(N__41766),
            .I(N__41763));
    Span4Mux_h I__9048 (
            .O(N__41763),
            .I(N__41760));
    Span4Mux_h I__9047 (
            .O(N__41760),
            .I(N__41757));
    Odrv4 I__9046 (
            .O(N__41757),
            .I(buf_data_iac_21));
    InMux I__9045 (
            .O(N__41754),
            .I(N__41751));
    LocalMux I__9044 (
            .O(N__41751),
            .I(N__41748));
    Span4Mux_h I__9043 (
            .O(N__41748),
            .I(N__41745));
    Span4Mux_v I__9042 (
            .O(N__41745),
            .I(N__41742));
    Odrv4 I__9041 (
            .O(N__41742),
            .I(n21672));
    CascadeMux I__9040 (
            .O(N__41739),
            .I(\ADC_VDC.n22124_cascade_ ));
    CascadeMux I__9039 (
            .O(N__41736),
            .I(N__41733));
    InMux I__9038 (
            .O(N__41733),
            .I(N__41730));
    LocalMux I__9037 (
            .O(N__41730),
            .I(N__41727));
    Span4Mux_h I__9036 (
            .O(N__41727),
            .I(N__41724));
    Span4Mux_h I__9035 (
            .O(N__41724),
            .I(N__41719));
    InMux I__9034 (
            .O(N__41723),
            .I(N__41714));
    InMux I__9033 (
            .O(N__41722),
            .I(N__41714));
    Odrv4 I__9032 (
            .O(N__41719),
            .I(buf_dds1_0));
    LocalMux I__9031 (
            .O(N__41714),
            .I(buf_dds1_0));
    CascadeMux I__9030 (
            .O(N__41709),
            .I(n16_cascade_));
    InMux I__9029 (
            .O(N__41706),
            .I(N__41702));
    InMux I__9028 (
            .O(N__41705),
            .I(N__41698));
    LocalMux I__9027 (
            .O(N__41702),
            .I(N__41695));
    CascadeMux I__9026 (
            .O(N__41701),
            .I(N__41692));
    LocalMux I__9025 (
            .O(N__41698),
            .I(N__41689));
    Span4Mux_v I__9024 (
            .O(N__41695),
            .I(N__41686));
    InMux I__9023 (
            .O(N__41692),
            .I(N__41683));
    Span4Mux_v I__9022 (
            .O(N__41689),
            .I(N__41680));
    Sp12to4 I__9021 (
            .O(N__41686),
            .I(N__41677));
    LocalMux I__9020 (
            .O(N__41683),
            .I(buf_adcdata_iac_8));
    Odrv4 I__9019 (
            .O(N__41680),
            .I(buf_adcdata_iac_8));
    Odrv12 I__9018 (
            .O(N__41677),
            .I(buf_adcdata_iac_8));
    CascadeMux I__9017 (
            .O(N__41670),
            .I(N__41659));
    InMux I__9016 (
            .O(N__41669),
            .I(N__41654));
    InMux I__9015 (
            .O(N__41668),
            .I(N__41651));
    InMux I__9014 (
            .O(N__41667),
            .I(N__41648));
    InMux I__9013 (
            .O(N__41666),
            .I(N__41645));
    InMux I__9012 (
            .O(N__41665),
            .I(N__41641));
    InMux I__9011 (
            .O(N__41664),
            .I(N__41638));
    InMux I__9010 (
            .O(N__41663),
            .I(N__41634));
    InMux I__9009 (
            .O(N__41662),
            .I(N__41631));
    InMux I__9008 (
            .O(N__41659),
            .I(N__41628));
    InMux I__9007 (
            .O(N__41658),
            .I(N__41625));
    InMux I__9006 (
            .O(N__41657),
            .I(N__41622));
    LocalMux I__9005 (
            .O(N__41654),
            .I(N__41619));
    LocalMux I__9004 (
            .O(N__41651),
            .I(N__41616));
    LocalMux I__9003 (
            .O(N__41648),
            .I(N__41610));
    LocalMux I__9002 (
            .O(N__41645),
            .I(N__41607));
    InMux I__9001 (
            .O(N__41644),
            .I(N__41604));
    LocalMux I__9000 (
            .O(N__41641),
            .I(N__41599));
    LocalMux I__8999 (
            .O(N__41638),
            .I(N__41599));
    InMux I__8998 (
            .O(N__41637),
            .I(N__41596));
    LocalMux I__8997 (
            .O(N__41634),
            .I(N__41591));
    LocalMux I__8996 (
            .O(N__41631),
            .I(N__41591));
    LocalMux I__8995 (
            .O(N__41628),
            .I(N__41584));
    LocalMux I__8994 (
            .O(N__41625),
            .I(N__41584));
    LocalMux I__8993 (
            .O(N__41622),
            .I(N__41584));
    Span4Mux_v I__8992 (
            .O(N__41619),
            .I(N__41579));
    Span4Mux_h I__8991 (
            .O(N__41616),
            .I(N__41579));
    InMux I__8990 (
            .O(N__41615),
            .I(N__41574));
    InMux I__8989 (
            .O(N__41614),
            .I(N__41574));
    InMux I__8988 (
            .O(N__41613),
            .I(N__41571));
    Span4Mux_h I__8987 (
            .O(N__41610),
            .I(N__41568));
    Span4Mux_h I__8986 (
            .O(N__41607),
            .I(N__41565));
    LocalMux I__8985 (
            .O(N__41604),
            .I(N__41560));
    Span4Mux_h I__8984 (
            .O(N__41599),
            .I(N__41560));
    LocalMux I__8983 (
            .O(N__41596),
            .I(N__41551));
    Span4Mux_h I__8982 (
            .O(N__41591),
            .I(N__41551));
    Span4Mux_v I__8981 (
            .O(N__41584),
            .I(N__41551));
    Span4Mux_v I__8980 (
            .O(N__41579),
            .I(N__41551));
    LocalMux I__8979 (
            .O(N__41574),
            .I(n12596));
    LocalMux I__8978 (
            .O(N__41571),
            .I(n12596));
    Odrv4 I__8977 (
            .O(N__41568),
            .I(n12596));
    Odrv4 I__8976 (
            .O(N__41565),
            .I(n12596));
    Odrv4 I__8975 (
            .O(N__41560),
            .I(n12596));
    Odrv4 I__8974 (
            .O(N__41551),
            .I(n12596));
    InMux I__8973 (
            .O(N__41538),
            .I(N__41535));
    LocalMux I__8972 (
            .O(N__41535),
            .I(N__41532));
    Span4Mux_v I__8971 (
            .O(N__41532),
            .I(N__41527));
    InMux I__8970 (
            .O(N__41531),
            .I(N__41522));
    InMux I__8969 (
            .O(N__41530),
            .I(N__41522));
    Odrv4 I__8968 (
            .O(N__41527),
            .I(buf_dds0_0));
    LocalMux I__8967 (
            .O(N__41522),
            .I(buf_dds0_0));
    IoInMux I__8966 (
            .O(N__41517),
            .I(N__41514));
    LocalMux I__8965 (
            .O(N__41514),
            .I(N__41511));
    Span4Mux_s2_h I__8964 (
            .O(N__41511),
            .I(N__41508));
    Span4Mux_h I__8963 (
            .O(N__41508),
            .I(N__41505));
    Sp12to4 I__8962 (
            .O(N__41505),
            .I(N__41502));
    Span12Mux_v I__8961 (
            .O(N__41502),
            .I(N__41498));
    CascadeMux I__8960 (
            .O(N__41501),
            .I(N__41494));
    Span12Mux_h I__8959 (
            .O(N__41498),
            .I(N__41491));
    InMux I__8958 (
            .O(N__41497),
            .I(N__41488));
    InMux I__8957 (
            .O(N__41494),
            .I(N__41485));
    Odrv12 I__8956 (
            .O(N__41491),
            .I(VDC_RNG0));
    LocalMux I__8955 (
            .O(N__41488),
            .I(VDC_RNG0));
    LocalMux I__8954 (
            .O(N__41485),
            .I(VDC_RNG0));
    CascadeMux I__8953 (
            .O(N__41478),
            .I(N__41475));
    InMux I__8952 (
            .O(N__41475),
            .I(N__41472));
    LocalMux I__8951 (
            .O(N__41472),
            .I(N__41469));
    Span4Mux_v I__8950 (
            .O(N__41469),
            .I(N__41466));
    Odrv4 I__8949 (
            .O(N__41466),
            .I(n23_adj_1675));
    InMux I__8948 (
            .O(N__41463),
            .I(N__41460));
    LocalMux I__8947 (
            .O(N__41460),
            .I(N__41457));
    Span4Mux_v I__8946 (
            .O(N__41457),
            .I(N__41452));
    InMux I__8945 (
            .O(N__41456),
            .I(N__41449));
    InMux I__8944 (
            .O(N__41455),
            .I(N__41446));
    Odrv4 I__8943 (
            .O(N__41452),
            .I(buf_dds0_6));
    LocalMux I__8942 (
            .O(N__41449),
            .I(buf_dds0_6));
    LocalMux I__8941 (
            .O(N__41446),
            .I(buf_dds0_6));
    InMux I__8940 (
            .O(N__41439),
            .I(N__41435));
    InMux I__8939 (
            .O(N__41438),
            .I(N__41432));
    LocalMux I__8938 (
            .O(N__41435),
            .I(n17705));
    LocalMux I__8937 (
            .O(N__41432),
            .I(n17705));
    CascadeMux I__8936 (
            .O(N__41427),
            .I(n9342_cascade_));
    CascadeMux I__8935 (
            .O(N__41424),
            .I(N__41421));
    InMux I__8934 (
            .O(N__41421),
            .I(N__41418));
    LocalMux I__8933 (
            .O(N__41418),
            .I(N__41414));
    InMux I__8932 (
            .O(N__41417),
            .I(N__41411));
    Odrv4 I__8931 (
            .O(N__41414),
            .I(n17703));
    LocalMux I__8930 (
            .O(N__41411),
            .I(n17703));
    CascadeMux I__8929 (
            .O(N__41406),
            .I(N__41403));
    CascadeBuf I__8928 (
            .O(N__41403),
            .I(N__41400));
    CascadeMux I__8927 (
            .O(N__41400),
            .I(N__41397));
    CascadeBuf I__8926 (
            .O(N__41397),
            .I(N__41394));
    CascadeMux I__8925 (
            .O(N__41394),
            .I(N__41391));
    CascadeBuf I__8924 (
            .O(N__41391),
            .I(N__41388));
    CascadeMux I__8923 (
            .O(N__41388),
            .I(N__41385));
    CascadeBuf I__8922 (
            .O(N__41385),
            .I(N__41382));
    CascadeMux I__8921 (
            .O(N__41382),
            .I(N__41379));
    CascadeBuf I__8920 (
            .O(N__41379),
            .I(N__41376));
    CascadeMux I__8919 (
            .O(N__41376),
            .I(N__41373));
    CascadeBuf I__8918 (
            .O(N__41373),
            .I(N__41370));
    CascadeMux I__8917 (
            .O(N__41370),
            .I(N__41366));
    CascadeMux I__8916 (
            .O(N__41369),
            .I(N__41363));
    CascadeBuf I__8915 (
            .O(N__41366),
            .I(N__41360));
    CascadeBuf I__8914 (
            .O(N__41363),
            .I(N__41357));
    CascadeMux I__8913 (
            .O(N__41360),
            .I(N__41354));
    CascadeMux I__8912 (
            .O(N__41357),
            .I(N__41351));
    CascadeBuf I__8911 (
            .O(N__41354),
            .I(N__41348));
    InMux I__8910 (
            .O(N__41351),
            .I(N__41345));
    CascadeMux I__8909 (
            .O(N__41348),
            .I(N__41342));
    LocalMux I__8908 (
            .O(N__41345),
            .I(N__41339));
    CascadeBuf I__8907 (
            .O(N__41342),
            .I(N__41336));
    Span4Mux_h I__8906 (
            .O(N__41339),
            .I(N__41333));
    CascadeMux I__8905 (
            .O(N__41336),
            .I(N__41330));
    Span4Mux_v I__8904 (
            .O(N__41333),
            .I(N__41327));
    InMux I__8903 (
            .O(N__41330),
            .I(N__41324));
    Span4Mux_v I__8902 (
            .O(N__41327),
            .I(N__41321));
    LocalMux I__8901 (
            .O(N__41324),
            .I(N__41318));
    Span4Mux_h I__8900 (
            .O(N__41321),
            .I(N__41315));
    Span4Mux_h I__8899 (
            .O(N__41318),
            .I(N__41312));
    Span4Mux_h I__8898 (
            .O(N__41315),
            .I(N__41307));
    Span4Mux_h I__8897 (
            .O(N__41312),
            .I(N__41307));
    Odrv4 I__8896 (
            .O(N__41307),
            .I(data_index_9_N_212_5));
    InMux I__8895 (
            .O(N__41304),
            .I(N__41300));
    InMux I__8894 (
            .O(N__41303),
            .I(N__41297));
    LocalMux I__8893 (
            .O(N__41300),
            .I(N__41293));
    LocalMux I__8892 (
            .O(N__41297),
            .I(N__41290));
    CascadeMux I__8891 (
            .O(N__41296),
            .I(N__41287));
    Span4Mux_h I__8890 (
            .O(N__41293),
            .I(N__41284));
    Span12Mux_s11_v I__8889 (
            .O(N__41290),
            .I(N__41281));
    InMux I__8888 (
            .O(N__41287),
            .I(N__41278));
    Span4Mux_h I__8887 (
            .O(N__41284),
            .I(N__41275));
    Span12Mux_h I__8886 (
            .O(N__41281),
            .I(N__41272));
    LocalMux I__8885 (
            .O(N__41278),
            .I(buf_adcdata_iac_11));
    Odrv4 I__8884 (
            .O(N__41275),
            .I(buf_adcdata_iac_11));
    Odrv12 I__8883 (
            .O(N__41272),
            .I(buf_adcdata_iac_11));
    InMux I__8882 (
            .O(N__41265),
            .I(N__41262));
    LocalMux I__8881 (
            .O(N__41262),
            .I(N__41259));
    Odrv12 I__8880 (
            .O(N__41259),
            .I(n16_adj_1640));
    CascadeMux I__8879 (
            .O(N__41256),
            .I(n22623_cascade_));
    CascadeMux I__8878 (
            .O(N__41253),
            .I(n22626_cascade_));
    InMux I__8877 (
            .O(N__41250),
            .I(N__41247));
    LocalMux I__8876 (
            .O(N__41247),
            .I(n30_adj_1643));
    InMux I__8875 (
            .O(N__41244),
            .I(N__41241));
    LocalMux I__8874 (
            .O(N__41241),
            .I(N__41238));
    Span4Mux_h I__8873 (
            .O(N__41238),
            .I(N__41234));
    InMux I__8872 (
            .O(N__41237),
            .I(N__41231));
    Span4Mux_h I__8871 (
            .O(N__41234),
            .I(N__41228));
    LocalMux I__8870 (
            .O(N__41231),
            .I(data_idxvec_3));
    Odrv4 I__8869 (
            .O(N__41228),
            .I(data_idxvec_3));
    InMux I__8868 (
            .O(N__41223),
            .I(N__41220));
    LocalMux I__8867 (
            .O(N__41220),
            .I(N__41216));
    InMux I__8866 (
            .O(N__41219),
            .I(N__41212));
    Span4Mux_v I__8865 (
            .O(N__41216),
            .I(N__41209));
    InMux I__8864 (
            .O(N__41215),
            .I(N__41206));
    LocalMux I__8863 (
            .O(N__41212),
            .I(data_cntvec_3));
    Odrv4 I__8862 (
            .O(N__41209),
            .I(data_cntvec_3));
    LocalMux I__8861 (
            .O(N__41206),
            .I(data_cntvec_3));
    CascadeMux I__8860 (
            .O(N__41199),
            .I(n26_adj_1642_cascade_));
    InMux I__8859 (
            .O(N__41196),
            .I(N__41193));
    LocalMux I__8858 (
            .O(N__41193),
            .I(N__41189));
    InMux I__8857 (
            .O(N__41192),
            .I(N__41185));
    Span4Mux_v I__8856 (
            .O(N__41189),
            .I(N__41182));
    InMux I__8855 (
            .O(N__41188),
            .I(N__41179));
    LocalMux I__8854 (
            .O(N__41185),
            .I(req_data_cnt_3));
    Odrv4 I__8853 (
            .O(N__41182),
            .I(req_data_cnt_3));
    LocalMux I__8852 (
            .O(N__41179),
            .I(req_data_cnt_3));
    CascadeMux I__8851 (
            .O(N__41172),
            .I(n22425_cascade_));
    InMux I__8850 (
            .O(N__41169),
            .I(N__41166));
    LocalMux I__8849 (
            .O(N__41166),
            .I(N__41163));
    Span4Mux_h I__8848 (
            .O(N__41163),
            .I(N__41158));
    InMux I__8847 (
            .O(N__41162),
            .I(N__41153));
    InMux I__8846 (
            .O(N__41161),
            .I(N__41153));
    Odrv4 I__8845 (
            .O(N__41158),
            .I(acadc_skipCount_3));
    LocalMux I__8844 (
            .O(N__41153),
            .I(acadc_skipCount_3));
    InMux I__8843 (
            .O(N__41148),
            .I(N__41145));
    LocalMux I__8842 (
            .O(N__41145),
            .I(n22428));
    InMux I__8841 (
            .O(N__41142),
            .I(N__41137));
    InMux I__8840 (
            .O(N__41141),
            .I(N__41134));
    InMux I__8839 (
            .O(N__41140),
            .I(N__41131));
    LocalMux I__8838 (
            .O(N__41137),
            .I(data_index_0));
    LocalMux I__8837 (
            .O(N__41134),
            .I(data_index_0));
    LocalMux I__8836 (
            .O(N__41131),
            .I(data_index_0));
    InMux I__8835 (
            .O(N__41124),
            .I(N__41116));
    InMux I__8834 (
            .O(N__41123),
            .I(N__41113));
    InMux I__8833 (
            .O(N__41122),
            .I(N__41108));
    InMux I__8832 (
            .O(N__41121),
            .I(N__41108));
    InMux I__8831 (
            .O(N__41120),
            .I(N__41103));
    InMux I__8830 (
            .O(N__41119),
            .I(N__41103));
    LocalMux I__8829 (
            .O(N__41116),
            .I(N__41097));
    LocalMux I__8828 (
            .O(N__41113),
            .I(N__41093));
    LocalMux I__8827 (
            .O(N__41108),
            .I(N__41088));
    LocalMux I__8826 (
            .O(N__41103),
            .I(N__41088));
    InMux I__8825 (
            .O(N__41102),
            .I(N__41085));
    InMux I__8824 (
            .O(N__41101),
            .I(N__41080));
    InMux I__8823 (
            .O(N__41100),
            .I(N__41080));
    Span4Mux_v I__8822 (
            .O(N__41097),
            .I(N__41076));
    InMux I__8821 (
            .O(N__41096),
            .I(N__41073));
    Span4Mux_v I__8820 (
            .O(N__41093),
            .I(N__41064));
    Span4Mux_v I__8819 (
            .O(N__41088),
            .I(N__41064));
    LocalMux I__8818 (
            .O(N__41085),
            .I(N__41064));
    LocalMux I__8817 (
            .O(N__41080),
            .I(N__41064));
    InMux I__8816 (
            .O(N__41079),
            .I(N__41061));
    Odrv4 I__8815 (
            .O(N__41076),
            .I(n8841));
    LocalMux I__8814 (
            .O(N__41073),
            .I(n8841));
    Odrv4 I__8813 (
            .O(N__41064),
            .I(n8841));
    LocalMux I__8812 (
            .O(N__41061),
            .I(n8841));
    InMux I__8811 (
            .O(N__41052),
            .I(N__41049));
    LocalMux I__8810 (
            .O(N__41049),
            .I(n8_adj_1540));
    InMux I__8809 (
            .O(N__41046),
            .I(N__41040));
    InMux I__8808 (
            .O(N__41045),
            .I(N__41040));
    LocalMux I__8807 (
            .O(N__41040),
            .I(n7_adj_1539));
    CascadeMux I__8806 (
            .O(N__41037),
            .I(n8_adj_1540_cascade_));
    CascadeMux I__8805 (
            .O(N__41034),
            .I(N__41031));
    CascadeBuf I__8804 (
            .O(N__41031),
            .I(N__41028));
    CascadeMux I__8803 (
            .O(N__41028),
            .I(N__41025));
    CascadeBuf I__8802 (
            .O(N__41025),
            .I(N__41022));
    CascadeMux I__8801 (
            .O(N__41022),
            .I(N__41019));
    CascadeBuf I__8800 (
            .O(N__41019),
            .I(N__41016));
    CascadeMux I__8799 (
            .O(N__41016),
            .I(N__41013));
    CascadeBuf I__8798 (
            .O(N__41013),
            .I(N__41010));
    CascadeMux I__8797 (
            .O(N__41010),
            .I(N__41007));
    CascadeBuf I__8796 (
            .O(N__41007),
            .I(N__41004));
    CascadeMux I__8795 (
            .O(N__41004),
            .I(N__41001));
    CascadeBuf I__8794 (
            .O(N__41001),
            .I(N__40998));
    CascadeMux I__8793 (
            .O(N__40998),
            .I(N__40995));
    CascadeBuf I__8792 (
            .O(N__40995),
            .I(N__40991));
    CascadeMux I__8791 (
            .O(N__40994),
            .I(N__40988));
    CascadeMux I__8790 (
            .O(N__40991),
            .I(N__40985));
    CascadeBuf I__8789 (
            .O(N__40988),
            .I(N__40982));
    CascadeBuf I__8788 (
            .O(N__40985),
            .I(N__40979));
    CascadeMux I__8787 (
            .O(N__40982),
            .I(N__40976));
    CascadeMux I__8786 (
            .O(N__40979),
            .I(N__40973));
    InMux I__8785 (
            .O(N__40976),
            .I(N__40970));
    CascadeBuf I__8784 (
            .O(N__40973),
            .I(N__40967));
    LocalMux I__8783 (
            .O(N__40970),
            .I(N__40964));
    CascadeMux I__8782 (
            .O(N__40967),
            .I(N__40961));
    Span4Mux_h I__8781 (
            .O(N__40964),
            .I(N__40958));
    InMux I__8780 (
            .O(N__40961),
            .I(N__40955));
    Span4Mux_v I__8779 (
            .O(N__40958),
            .I(N__40952));
    LocalMux I__8778 (
            .O(N__40955),
            .I(N__40949));
    Span4Mux_h I__8777 (
            .O(N__40952),
            .I(N__40946));
    Span4Mux_h I__8776 (
            .O(N__40949),
            .I(N__40943));
    Span4Mux_h I__8775 (
            .O(N__40946),
            .I(N__40940));
    Span4Mux_v I__8774 (
            .O(N__40943),
            .I(N__40937));
    Odrv4 I__8773 (
            .O(N__40940),
            .I(data_index_9_N_212_0));
    Odrv4 I__8772 (
            .O(N__40937),
            .I(data_index_9_N_212_0));
    CascadeMux I__8771 (
            .O(N__40932),
            .I(n30_adj_1688_cascade_));
    InMux I__8770 (
            .O(N__40929),
            .I(N__40926));
    LocalMux I__8769 (
            .O(N__40926),
            .I(N__40922));
    CascadeMux I__8768 (
            .O(N__40925),
            .I(N__40919));
    Span4Mux_h I__8767 (
            .O(N__40922),
            .I(N__40916));
    InMux I__8766 (
            .O(N__40919),
            .I(N__40913));
    Span4Mux_h I__8765 (
            .O(N__40916),
            .I(N__40910));
    LocalMux I__8764 (
            .O(N__40913),
            .I(data_idxvec_8));
    Odrv4 I__8763 (
            .O(N__40910),
            .I(data_idxvec_8));
    InMux I__8762 (
            .O(N__40905),
            .I(N__40902));
    LocalMux I__8761 (
            .O(N__40902),
            .I(N__40898));
    InMux I__8760 (
            .O(N__40901),
            .I(N__40894));
    Span4Mux_v I__8759 (
            .O(N__40898),
            .I(N__40891));
    InMux I__8758 (
            .O(N__40897),
            .I(N__40888));
    LocalMux I__8757 (
            .O(N__40894),
            .I(data_cntvec_8));
    Odrv4 I__8756 (
            .O(N__40891),
            .I(data_cntvec_8));
    LocalMux I__8755 (
            .O(N__40888),
            .I(data_cntvec_8));
    InMux I__8754 (
            .O(N__40881),
            .I(N__40878));
    LocalMux I__8753 (
            .O(N__40878),
            .I(N__40875));
    Span4Mux_h I__8752 (
            .O(N__40875),
            .I(N__40872));
    Span4Mux_h I__8751 (
            .O(N__40872),
            .I(N__40869));
    Odrv4 I__8750 (
            .O(N__40869),
            .I(buf_data_iac_16));
    CascadeMux I__8749 (
            .O(N__40866),
            .I(n26_adj_1533_cascade_));
    InMux I__8748 (
            .O(N__40863),
            .I(N__40860));
    LocalMux I__8747 (
            .O(N__40860),
            .I(N__40857));
    Odrv12 I__8746 (
            .O(N__40857),
            .I(n22398));
    CascadeMux I__8745 (
            .O(N__40854),
            .I(n21246_cascade_));
    InMux I__8744 (
            .O(N__40851),
            .I(N__40848));
    LocalMux I__8743 (
            .O(N__40848),
            .I(N__40845));
    Span4Mux_h I__8742 (
            .O(N__40845),
            .I(N__40842));
    Odrv4 I__8741 (
            .O(N__40842),
            .I(n22392));
    InMux I__8740 (
            .O(N__40839),
            .I(N__40836));
    LocalMux I__8739 (
            .O(N__40836),
            .I(N__40833));
    Span4Mux_v I__8738 (
            .O(N__40833),
            .I(N__40830));
    Span4Mux_h I__8737 (
            .O(N__40830),
            .I(N__40827));
    Odrv4 I__8736 (
            .O(N__40827),
            .I(n22578));
    CascadeMux I__8735 (
            .O(N__40824),
            .I(n22581_cascade_));
    CascadeMux I__8734 (
            .O(N__40821),
            .I(n22584_cascade_));
    InMux I__8733 (
            .O(N__40818),
            .I(N__40815));
    LocalMux I__8732 (
            .O(N__40815),
            .I(N__40812));
    Span4Mux_h I__8731 (
            .O(N__40812),
            .I(N__40809));
    Span4Mux_h I__8730 (
            .O(N__40809),
            .I(N__40806));
    Span4Mux_h I__8729 (
            .O(N__40806),
            .I(N__40802));
    InMux I__8728 (
            .O(N__40805),
            .I(N__40799));
    Odrv4 I__8727 (
            .O(N__40802),
            .I(buf_readRTD_3));
    LocalMux I__8726 (
            .O(N__40799),
            .I(buf_readRTD_3));
    CascadeMux I__8725 (
            .O(N__40794),
            .I(N__40791));
    InMux I__8724 (
            .O(N__40791),
            .I(N__40788));
    LocalMux I__8723 (
            .O(N__40788),
            .I(N__40785));
    Span4Mux_v I__8722 (
            .O(N__40785),
            .I(N__40782));
    Odrv4 I__8721 (
            .O(N__40782),
            .I(n19_adj_1641));
    CascadeMux I__8720 (
            .O(N__40779),
            .I(n21556_cascade_));
    InMux I__8719 (
            .O(N__40776),
            .I(N__40773));
    LocalMux I__8718 (
            .O(N__40773),
            .I(N__40770));
    Span4Mux_v I__8717 (
            .O(N__40770),
            .I(N__40767));
    Odrv4 I__8716 (
            .O(N__40767),
            .I(n21703));
    InMux I__8715 (
            .O(N__40764),
            .I(N__40761));
    LocalMux I__8714 (
            .O(N__40761),
            .I(n22521));
    InMux I__8713 (
            .O(N__40758),
            .I(N__40755));
    LocalMux I__8712 (
            .O(N__40755),
            .I(n22464));
    CascadeMux I__8711 (
            .O(N__40752),
            .I(n22524_cascade_));
    CascadeMux I__8710 (
            .O(N__40749),
            .I(n30_adj_1676_cascade_));
    InMux I__8709 (
            .O(N__40746),
            .I(N__40743));
    LocalMux I__8708 (
            .O(N__40743),
            .I(N__40740));
    Span4Mux_h I__8707 (
            .O(N__40740),
            .I(N__40737));
    Span4Mux_h I__8706 (
            .O(N__40737),
            .I(N__40734));
    Odrv4 I__8705 (
            .O(N__40734),
            .I(n17_adj_1682));
    CascadeMux I__8704 (
            .O(N__40731),
            .I(N__40728));
    InMux I__8703 (
            .O(N__40728),
            .I(N__40725));
    LocalMux I__8702 (
            .O(N__40725),
            .I(N__40722));
    Span4Mux_v I__8701 (
            .O(N__40722),
            .I(N__40719));
    Odrv4 I__8700 (
            .O(N__40719),
            .I(n16_adj_1681));
    InMux I__8699 (
            .O(N__40716),
            .I(N__40713));
    LocalMux I__8698 (
            .O(N__40713),
            .I(N__40710));
    Span4Mux_h I__8697 (
            .O(N__40710),
            .I(N__40707));
    Odrv4 I__8696 (
            .O(N__40707),
            .I(n22485));
    InMux I__8695 (
            .O(N__40704),
            .I(N__40700));
    CascadeMux I__8694 (
            .O(N__40703),
            .I(N__40697));
    LocalMux I__8693 (
            .O(N__40700),
            .I(N__40694));
    InMux I__8692 (
            .O(N__40697),
            .I(N__40691));
    Span12Mux_v I__8691 (
            .O(N__40694),
            .I(N__40688));
    LocalMux I__8690 (
            .O(N__40691),
            .I(data_idxvec_10));
    Odrv12 I__8689 (
            .O(N__40688),
            .I(data_idxvec_10));
    InMux I__8688 (
            .O(N__40683),
            .I(N__40679));
    InMux I__8687 (
            .O(N__40682),
            .I(N__40675));
    LocalMux I__8686 (
            .O(N__40679),
            .I(N__40672));
    InMux I__8685 (
            .O(N__40678),
            .I(N__40669));
    LocalMux I__8684 (
            .O(N__40675),
            .I(N__40666));
    Span4Mux_v I__8683 (
            .O(N__40672),
            .I(N__40663));
    LocalMux I__8682 (
            .O(N__40669),
            .I(data_cntvec_10));
    Odrv4 I__8681 (
            .O(N__40666),
            .I(data_cntvec_10));
    Odrv4 I__8680 (
            .O(N__40663),
            .I(data_cntvec_10));
    CascadeMux I__8679 (
            .O(N__40656),
            .I(n26_adj_1687_cascade_));
    CascadeMux I__8678 (
            .O(N__40653),
            .I(n22455_cascade_));
    InMux I__8677 (
            .O(N__40650),
            .I(N__40647));
    LocalMux I__8676 (
            .O(N__40647),
            .I(N__40644));
    Span4Mux_v I__8675 (
            .O(N__40644),
            .I(N__40641));
    Span4Mux_h I__8674 (
            .O(N__40641),
            .I(N__40638));
    Sp12to4 I__8673 (
            .O(N__40638),
            .I(N__40635));
    Odrv12 I__8672 (
            .O(N__40635),
            .I(n24_adj_1686));
    InMux I__8671 (
            .O(N__40632),
            .I(N__40629));
    LocalMux I__8670 (
            .O(N__40629),
            .I(n22488));
    CascadeMux I__8669 (
            .O(N__40626),
            .I(n22458_cascade_));
    ClkMux I__8668 (
            .O(N__40623),
            .I(N__40618));
    ClkMux I__8667 (
            .O(N__40622),
            .I(N__40604));
    ClkMux I__8666 (
            .O(N__40621),
            .I(N__40601));
    LocalMux I__8665 (
            .O(N__40618),
            .I(N__40598));
    ClkMux I__8664 (
            .O(N__40617),
            .I(N__40595));
    ClkMux I__8663 (
            .O(N__40616),
            .I(N__40592));
    ClkMux I__8662 (
            .O(N__40615),
            .I(N__40589));
    ClkMux I__8661 (
            .O(N__40614),
            .I(N__40586));
    ClkMux I__8660 (
            .O(N__40613),
            .I(N__40583));
    ClkMux I__8659 (
            .O(N__40612),
            .I(N__40579));
    ClkMux I__8658 (
            .O(N__40611),
            .I(N__40576));
    ClkMux I__8657 (
            .O(N__40610),
            .I(N__40573));
    ClkMux I__8656 (
            .O(N__40609),
            .I(N__40570));
    ClkMux I__8655 (
            .O(N__40608),
            .I(N__40566));
    ClkMux I__8654 (
            .O(N__40607),
            .I(N__40563));
    LocalMux I__8653 (
            .O(N__40604),
            .I(N__40558));
    LocalMux I__8652 (
            .O(N__40601),
            .I(N__40558));
    Span4Mux_v I__8651 (
            .O(N__40598),
            .I(N__40555));
    LocalMux I__8650 (
            .O(N__40595),
            .I(N__40550));
    LocalMux I__8649 (
            .O(N__40592),
            .I(N__40550));
    LocalMux I__8648 (
            .O(N__40589),
            .I(N__40547));
    LocalMux I__8647 (
            .O(N__40586),
            .I(N__40542));
    LocalMux I__8646 (
            .O(N__40583),
            .I(N__40542));
    ClkMux I__8645 (
            .O(N__40582),
            .I(N__40539));
    LocalMux I__8644 (
            .O(N__40579),
            .I(N__40535));
    LocalMux I__8643 (
            .O(N__40576),
            .I(N__40530));
    LocalMux I__8642 (
            .O(N__40573),
            .I(N__40530));
    LocalMux I__8641 (
            .O(N__40570),
            .I(N__40527));
    ClkMux I__8640 (
            .O(N__40569),
            .I(N__40524));
    LocalMux I__8639 (
            .O(N__40566),
            .I(N__40519));
    LocalMux I__8638 (
            .O(N__40563),
            .I(N__40519));
    Span4Mux_v I__8637 (
            .O(N__40558),
            .I(N__40516));
    Span4Mux_v I__8636 (
            .O(N__40555),
            .I(N__40505));
    Span4Mux_v I__8635 (
            .O(N__40550),
            .I(N__40505));
    Span4Mux_h I__8634 (
            .O(N__40547),
            .I(N__40505));
    Span4Mux_v I__8633 (
            .O(N__40542),
            .I(N__40505));
    LocalMux I__8632 (
            .O(N__40539),
            .I(N__40505));
    ClkMux I__8631 (
            .O(N__40538),
            .I(N__40502));
    Span4Mux_v I__8630 (
            .O(N__40535),
            .I(N__40497));
    Span4Mux_v I__8629 (
            .O(N__40530),
            .I(N__40497));
    Span4Mux_v I__8628 (
            .O(N__40527),
            .I(N__40492));
    LocalMux I__8627 (
            .O(N__40524),
            .I(N__40492));
    Span4Mux_v I__8626 (
            .O(N__40519),
            .I(N__40485));
    Span4Mux_h I__8625 (
            .O(N__40516),
            .I(N__40485));
    Span4Mux_h I__8624 (
            .O(N__40505),
            .I(N__40485));
    LocalMux I__8623 (
            .O(N__40502),
            .I(N__40482));
    Span4Mux_h I__8622 (
            .O(N__40497),
            .I(N__40477));
    Span4Mux_h I__8621 (
            .O(N__40492),
            .I(N__40477));
    Span4Mux_h I__8620 (
            .O(N__40485),
            .I(N__40474));
    Span12Mux_h I__8619 (
            .O(N__40482),
            .I(N__40470));
    Span4Mux_h I__8618 (
            .O(N__40477),
            .I(N__40467));
    Span4Mux_h I__8617 (
            .O(N__40474),
            .I(N__40464));
    InMux I__8616 (
            .O(N__40473),
            .I(N__40461));
    Odrv12 I__8615 (
            .O(N__40470),
            .I(clk_RTD));
    Odrv4 I__8614 (
            .O(N__40467),
            .I(clk_RTD));
    Odrv4 I__8613 (
            .O(N__40464),
            .I(clk_RTD));
    LocalMux I__8612 (
            .O(N__40461),
            .I(clk_RTD));
    InMux I__8611 (
            .O(N__40452),
            .I(N__40449));
    LocalMux I__8610 (
            .O(N__40449),
            .I(N__40444));
    InMux I__8609 (
            .O(N__40448),
            .I(N__40441));
    InMux I__8608 (
            .O(N__40447),
            .I(N__40438));
    Span4Mux_h I__8607 (
            .O(N__40444),
            .I(N__40435));
    LocalMux I__8606 (
            .O(N__40441),
            .I(N__40430));
    LocalMux I__8605 (
            .O(N__40438),
            .I(N__40430));
    Span4Mux_h I__8604 (
            .O(N__40435),
            .I(N__40427));
    Odrv12 I__8603 (
            .O(N__40430),
            .I(n14_adj_1550));
    Odrv4 I__8602 (
            .O(N__40427),
            .I(n14_adj_1550));
    InMux I__8601 (
            .O(N__40422),
            .I(N__40419));
    LocalMux I__8600 (
            .O(N__40419),
            .I(N__40416));
    Odrv12 I__8599 (
            .O(N__40416),
            .I(n17_adj_1672));
    InMux I__8598 (
            .O(N__40413),
            .I(N__40410));
    LocalMux I__8597 (
            .O(N__40410),
            .I(N__40407));
    Span4Mux_h I__8596 (
            .O(N__40407),
            .I(N__40404));
    Odrv4 I__8595 (
            .O(N__40404),
            .I(n22461));
    CascadeMux I__8594 (
            .O(N__40401),
            .I(N__40398));
    InMux I__8593 (
            .O(N__40398),
            .I(N__40395));
    LocalMux I__8592 (
            .O(N__40395),
            .I(N__40392));
    Span4Mux_v I__8591 (
            .O(N__40392),
            .I(N__40389));
    Span4Mux_v I__8590 (
            .O(N__40389),
            .I(N__40386));
    Odrv4 I__8589 (
            .O(N__40386),
            .I(n16_adj_1671));
    InMux I__8588 (
            .O(N__40383),
            .I(N__40380));
    LocalMux I__8587 (
            .O(N__40380),
            .I(N__40376));
    CascadeMux I__8586 (
            .O(N__40379),
            .I(N__40373));
    Span4Mux_h I__8585 (
            .O(N__40376),
            .I(N__40370));
    InMux I__8584 (
            .O(N__40373),
            .I(N__40367));
    Span4Mux_h I__8583 (
            .O(N__40370),
            .I(N__40364));
    LocalMux I__8582 (
            .O(N__40367),
            .I(data_idxvec_12));
    Odrv4 I__8581 (
            .O(N__40364),
            .I(data_idxvec_12));
    InMux I__8580 (
            .O(N__40359),
            .I(N__40355));
    InMux I__8579 (
            .O(N__40358),
            .I(N__40352));
    LocalMux I__8578 (
            .O(N__40355),
            .I(wdtick_cnt_22));
    LocalMux I__8577 (
            .O(N__40352),
            .I(wdtick_cnt_22));
    InMux I__8576 (
            .O(N__40347),
            .I(n19953));
    InMux I__8575 (
            .O(N__40344),
            .I(N__40340));
    InMux I__8574 (
            .O(N__40343),
            .I(N__40337));
    LocalMux I__8573 (
            .O(N__40340),
            .I(wdtick_cnt_23));
    LocalMux I__8572 (
            .O(N__40337),
            .I(wdtick_cnt_23));
    InMux I__8571 (
            .O(N__40332),
            .I(n19954));
    InMux I__8570 (
            .O(N__40329),
            .I(N__40296));
    InMux I__8569 (
            .O(N__40328),
            .I(N__40296));
    InMux I__8568 (
            .O(N__40327),
            .I(N__40296));
    InMux I__8567 (
            .O(N__40326),
            .I(N__40296));
    InMux I__8566 (
            .O(N__40325),
            .I(N__40293));
    InMux I__8565 (
            .O(N__40324),
            .I(N__40284));
    InMux I__8564 (
            .O(N__40323),
            .I(N__40284));
    InMux I__8563 (
            .O(N__40322),
            .I(N__40284));
    InMux I__8562 (
            .O(N__40321),
            .I(N__40284));
    InMux I__8561 (
            .O(N__40320),
            .I(N__40275));
    InMux I__8560 (
            .O(N__40319),
            .I(N__40275));
    InMux I__8559 (
            .O(N__40318),
            .I(N__40275));
    InMux I__8558 (
            .O(N__40317),
            .I(N__40275));
    InMux I__8557 (
            .O(N__40316),
            .I(N__40266));
    InMux I__8556 (
            .O(N__40315),
            .I(N__40266));
    InMux I__8555 (
            .O(N__40314),
            .I(N__40266));
    InMux I__8554 (
            .O(N__40313),
            .I(N__40266));
    InMux I__8553 (
            .O(N__40312),
            .I(N__40257));
    InMux I__8552 (
            .O(N__40311),
            .I(N__40257));
    InMux I__8551 (
            .O(N__40310),
            .I(N__40257));
    InMux I__8550 (
            .O(N__40309),
            .I(N__40257));
    InMux I__8549 (
            .O(N__40308),
            .I(N__40248));
    InMux I__8548 (
            .O(N__40307),
            .I(N__40248));
    InMux I__8547 (
            .O(N__40306),
            .I(N__40248));
    InMux I__8546 (
            .O(N__40305),
            .I(N__40248));
    LocalMux I__8545 (
            .O(N__40296),
            .I(N__40243));
    LocalMux I__8544 (
            .O(N__40293),
            .I(N__40243));
    LocalMux I__8543 (
            .O(N__40284),
            .I(n49));
    LocalMux I__8542 (
            .O(N__40275),
            .I(n49));
    LocalMux I__8541 (
            .O(N__40266),
            .I(n49));
    LocalMux I__8540 (
            .O(N__40257),
            .I(n49));
    LocalMux I__8539 (
            .O(N__40248),
            .I(n49));
    Odrv4 I__8538 (
            .O(N__40243),
            .I(n49));
    InMux I__8537 (
            .O(N__40230),
            .I(bfn_15_8_0_));
    InMux I__8536 (
            .O(N__40227),
            .I(N__40223));
    InMux I__8535 (
            .O(N__40226),
            .I(N__40220));
    LocalMux I__8534 (
            .O(N__40223),
            .I(N__40217));
    LocalMux I__8533 (
            .O(N__40220),
            .I(wdtick_cnt_24));
    Odrv4 I__8532 (
            .O(N__40217),
            .I(wdtick_cnt_24));
    InMux I__8531 (
            .O(N__40212),
            .I(N__40208));
    InMux I__8530 (
            .O(N__40211),
            .I(N__40205));
    LocalMux I__8529 (
            .O(N__40208),
            .I(N__40200));
    LocalMux I__8528 (
            .O(N__40205),
            .I(N__40200));
    Odrv4 I__8527 (
            .O(N__40200),
            .I(wdtick_cnt_14));
    InMux I__8526 (
            .O(N__40197),
            .I(n19945));
    InMux I__8525 (
            .O(N__40194),
            .I(N__40190));
    InMux I__8524 (
            .O(N__40193),
            .I(N__40187));
    LocalMux I__8523 (
            .O(N__40190),
            .I(wdtick_cnt_15));
    LocalMux I__8522 (
            .O(N__40187),
            .I(wdtick_cnt_15));
    InMux I__8521 (
            .O(N__40182),
            .I(n19946));
    InMux I__8520 (
            .O(N__40179),
            .I(N__40175));
    InMux I__8519 (
            .O(N__40178),
            .I(N__40172));
    LocalMux I__8518 (
            .O(N__40175),
            .I(wdtick_cnt_16));
    LocalMux I__8517 (
            .O(N__40172),
            .I(wdtick_cnt_16));
    InMux I__8516 (
            .O(N__40167),
            .I(bfn_15_7_0_));
    InMux I__8515 (
            .O(N__40164),
            .I(N__40160));
    InMux I__8514 (
            .O(N__40163),
            .I(N__40157));
    LocalMux I__8513 (
            .O(N__40160),
            .I(wdtick_cnt_17));
    LocalMux I__8512 (
            .O(N__40157),
            .I(wdtick_cnt_17));
    InMux I__8511 (
            .O(N__40152),
            .I(n19948));
    CascadeMux I__8510 (
            .O(N__40149),
            .I(N__40145));
    InMux I__8509 (
            .O(N__40148),
            .I(N__40142));
    InMux I__8508 (
            .O(N__40145),
            .I(N__40139));
    LocalMux I__8507 (
            .O(N__40142),
            .I(wdtick_cnt_18));
    LocalMux I__8506 (
            .O(N__40139),
            .I(wdtick_cnt_18));
    InMux I__8505 (
            .O(N__40134),
            .I(n19949));
    CascadeMux I__8504 (
            .O(N__40131),
            .I(N__40127));
    InMux I__8503 (
            .O(N__40130),
            .I(N__40124));
    InMux I__8502 (
            .O(N__40127),
            .I(N__40121));
    LocalMux I__8501 (
            .O(N__40124),
            .I(wdtick_cnt_19));
    LocalMux I__8500 (
            .O(N__40121),
            .I(wdtick_cnt_19));
    InMux I__8499 (
            .O(N__40116),
            .I(n19950));
    CascadeMux I__8498 (
            .O(N__40113),
            .I(N__40109));
    InMux I__8497 (
            .O(N__40112),
            .I(N__40106));
    InMux I__8496 (
            .O(N__40109),
            .I(N__40103));
    LocalMux I__8495 (
            .O(N__40106),
            .I(wdtick_cnt_20));
    LocalMux I__8494 (
            .O(N__40103),
            .I(wdtick_cnt_20));
    InMux I__8493 (
            .O(N__40098),
            .I(n19951));
    InMux I__8492 (
            .O(N__40095),
            .I(N__40091));
    InMux I__8491 (
            .O(N__40094),
            .I(N__40088));
    LocalMux I__8490 (
            .O(N__40091),
            .I(wdtick_cnt_21));
    LocalMux I__8489 (
            .O(N__40088),
            .I(wdtick_cnt_21));
    InMux I__8488 (
            .O(N__40083),
            .I(n19952));
    CascadeMux I__8487 (
            .O(N__40080),
            .I(N__40077));
    InMux I__8486 (
            .O(N__40077),
            .I(N__40074));
    LocalMux I__8485 (
            .O(N__40074),
            .I(N__40070));
    InMux I__8484 (
            .O(N__40073),
            .I(N__40067));
    Span4Mux_h I__8483 (
            .O(N__40070),
            .I(N__40064));
    LocalMux I__8482 (
            .O(N__40067),
            .I(wdtick_cnt_6));
    Odrv4 I__8481 (
            .O(N__40064),
            .I(wdtick_cnt_6));
    InMux I__8480 (
            .O(N__40059),
            .I(n19937));
    InMux I__8479 (
            .O(N__40056),
            .I(N__40052));
    InMux I__8478 (
            .O(N__40055),
            .I(N__40049));
    LocalMux I__8477 (
            .O(N__40052),
            .I(N__40046));
    LocalMux I__8476 (
            .O(N__40049),
            .I(wdtick_cnt_7));
    Odrv4 I__8475 (
            .O(N__40046),
            .I(wdtick_cnt_7));
    InMux I__8474 (
            .O(N__40041),
            .I(n19938));
    CascadeMux I__8473 (
            .O(N__40038),
            .I(N__40035));
    InMux I__8472 (
            .O(N__40035),
            .I(N__40031));
    InMux I__8471 (
            .O(N__40034),
            .I(N__40028));
    LocalMux I__8470 (
            .O(N__40031),
            .I(N__40025));
    LocalMux I__8469 (
            .O(N__40028),
            .I(wdtick_cnt_8));
    Odrv4 I__8468 (
            .O(N__40025),
            .I(wdtick_cnt_8));
    InMux I__8467 (
            .O(N__40020),
            .I(bfn_15_6_0_));
    InMux I__8466 (
            .O(N__40017),
            .I(N__40013));
    InMux I__8465 (
            .O(N__40016),
            .I(N__40010));
    LocalMux I__8464 (
            .O(N__40013),
            .I(wdtick_cnt_9));
    LocalMux I__8463 (
            .O(N__40010),
            .I(wdtick_cnt_9));
    InMux I__8462 (
            .O(N__40005),
            .I(n19940));
    InMux I__8461 (
            .O(N__40002),
            .I(N__39999));
    LocalMux I__8460 (
            .O(N__39999),
            .I(N__39995));
    InMux I__8459 (
            .O(N__39998),
            .I(N__39992));
    Span4Mux_h I__8458 (
            .O(N__39995),
            .I(N__39989));
    LocalMux I__8457 (
            .O(N__39992),
            .I(wdtick_cnt_10));
    Odrv4 I__8456 (
            .O(N__39989),
            .I(wdtick_cnt_10));
    InMux I__8455 (
            .O(N__39984),
            .I(n19941));
    InMux I__8454 (
            .O(N__39981),
            .I(N__39977));
    InMux I__8453 (
            .O(N__39980),
            .I(N__39974));
    LocalMux I__8452 (
            .O(N__39977),
            .I(wdtick_cnt_11));
    LocalMux I__8451 (
            .O(N__39974),
            .I(wdtick_cnt_11));
    InMux I__8450 (
            .O(N__39969),
            .I(n19942));
    InMux I__8449 (
            .O(N__39966),
            .I(N__39963));
    LocalMux I__8448 (
            .O(N__39963),
            .I(N__39959));
    InMux I__8447 (
            .O(N__39962),
            .I(N__39956));
    Span4Mux_v I__8446 (
            .O(N__39959),
            .I(N__39953));
    LocalMux I__8445 (
            .O(N__39956),
            .I(wdtick_cnt_12));
    Odrv4 I__8444 (
            .O(N__39953),
            .I(wdtick_cnt_12));
    InMux I__8443 (
            .O(N__39948),
            .I(n19943));
    InMux I__8442 (
            .O(N__39945),
            .I(N__39941));
    InMux I__8441 (
            .O(N__39944),
            .I(N__39938));
    LocalMux I__8440 (
            .O(N__39941),
            .I(wdtick_cnt_13));
    LocalMux I__8439 (
            .O(N__39938),
            .I(wdtick_cnt_13));
    InMux I__8438 (
            .O(N__39933),
            .I(n19944));
    CascadeMux I__8437 (
            .O(N__39930),
            .I(N__39926));
    CascadeMux I__8436 (
            .O(N__39929),
            .I(N__39923));
    InMux I__8435 (
            .O(N__39926),
            .I(N__39918));
    InMux I__8434 (
            .O(N__39923),
            .I(N__39918));
    LocalMux I__8433 (
            .O(N__39918),
            .I(n8_adj_1568));
    InMux I__8432 (
            .O(N__39915),
            .I(N__39909));
    InMux I__8431 (
            .O(N__39914),
            .I(N__39909));
    LocalMux I__8430 (
            .O(N__39909),
            .I(N__39906));
    Odrv12 I__8429 (
            .O(N__39906),
            .I(n7_adj_1567));
    CascadeMux I__8428 (
            .O(N__39903),
            .I(N__39900));
    CascadeBuf I__8427 (
            .O(N__39900),
            .I(N__39897));
    CascadeMux I__8426 (
            .O(N__39897),
            .I(N__39894));
    CascadeBuf I__8425 (
            .O(N__39894),
            .I(N__39891));
    CascadeMux I__8424 (
            .O(N__39891),
            .I(N__39888));
    CascadeBuf I__8423 (
            .O(N__39888),
            .I(N__39885));
    CascadeMux I__8422 (
            .O(N__39885),
            .I(N__39882));
    CascadeBuf I__8421 (
            .O(N__39882),
            .I(N__39879));
    CascadeMux I__8420 (
            .O(N__39879),
            .I(N__39876));
    CascadeBuf I__8419 (
            .O(N__39876),
            .I(N__39873));
    CascadeMux I__8418 (
            .O(N__39873),
            .I(N__39870));
    CascadeBuf I__8417 (
            .O(N__39870),
            .I(N__39867));
    CascadeMux I__8416 (
            .O(N__39867),
            .I(N__39864));
    CascadeBuf I__8415 (
            .O(N__39864),
            .I(N__39860));
    CascadeMux I__8414 (
            .O(N__39863),
            .I(N__39857));
    CascadeMux I__8413 (
            .O(N__39860),
            .I(N__39854));
    CascadeBuf I__8412 (
            .O(N__39857),
            .I(N__39851));
    CascadeBuf I__8411 (
            .O(N__39854),
            .I(N__39848));
    CascadeMux I__8410 (
            .O(N__39851),
            .I(N__39845));
    CascadeMux I__8409 (
            .O(N__39848),
            .I(N__39842));
    InMux I__8408 (
            .O(N__39845),
            .I(N__39839));
    CascadeBuf I__8407 (
            .O(N__39842),
            .I(N__39836));
    LocalMux I__8406 (
            .O(N__39839),
            .I(N__39833));
    CascadeMux I__8405 (
            .O(N__39836),
            .I(N__39830));
    Span12Mux_h I__8404 (
            .O(N__39833),
            .I(N__39827));
    InMux I__8403 (
            .O(N__39830),
            .I(N__39824));
    Span12Mux_v I__8402 (
            .O(N__39827),
            .I(N__39821));
    LocalMux I__8401 (
            .O(N__39824),
            .I(N__39818));
    Odrv12 I__8400 (
            .O(N__39821),
            .I(data_index_9_N_212_2));
    Odrv12 I__8399 (
            .O(N__39818),
            .I(data_index_9_N_212_2));
    InMux I__8398 (
            .O(N__39813),
            .I(N__39809));
    InMux I__8397 (
            .O(N__39812),
            .I(N__39806));
    LocalMux I__8396 (
            .O(N__39809),
            .I(N__39803));
    LocalMux I__8395 (
            .O(N__39806),
            .I(\comm_spi.n14815 ));
    Odrv4 I__8394 (
            .O(N__39803),
            .I(\comm_spi.n14815 ));
    InMux I__8393 (
            .O(N__39798),
            .I(N__39794));
    InMux I__8392 (
            .O(N__39797),
            .I(N__39791));
    LocalMux I__8391 (
            .O(N__39794),
            .I(\comm_spi.n14816 ));
    LocalMux I__8390 (
            .O(N__39791),
            .I(\comm_spi.n14816 ));
    InMux I__8389 (
            .O(N__39786),
            .I(N__39782));
    InMux I__8388 (
            .O(N__39785),
            .I(N__39779));
    LocalMux I__8387 (
            .O(N__39782),
            .I(\comm_spi.imosi ));
    LocalMux I__8386 (
            .O(N__39779),
            .I(\comm_spi.imosi ));
    SRMux I__8385 (
            .O(N__39774),
            .I(N__39771));
    LocalMux I__8384 (
            .O(N__39771),
            .I(N__39768));
    Span4Mux_v I__8383 (
            .O(N__39768),
            .I(N__39765));
    Span4Mux_v I__8382 (
            .O(N__39765),
            .I(N__39762));
    Odrv4 I__8381 (
            .O(N__39762),
            .I(\comm_spi.DOUT_7__N_787 ));
    InMux I__8380 (
            .O(N__39759),
            .I(N__39755));
    InMux I__8379 (
            .O(N__39758),
            .I(N__39752));
    LocalMux I__8378 (
            .O(N__39755),
            .I(wdtick_cnt_0));
    LocalMux I__8377 (
            .O(N__39752),
            .I(wdtick_cnt_0));
    InMux I__8376 (
            .O(N__39747),
            .I(bfn_15_5_0_));
    InMux I__8375 (
            .O(N__39744),
            .I(N__39741));
    LocalMux I__8374 (
            .O(N__39741),
            .I(N__39737));
    InMux I__8373 (
            .O(N__39740),
            .I(N__39734));
    Span4Mux_h I__8372 (
            .O(N__39737),
            .I(N__39731));
    LocalMux I__8371 (
            .O(N__39734),
            .I(wdtick_cnt_1));
    Odrv4 I__8370 (
            .O(N__39731),
            .I(wdtick_cnt_1));
    InMux I__8369 (
            .O(N__39726),
            .I(n19932));
    InMux I__8368 (
            .O(N__39723),
            .I(N__39719));
    InMux I__8367 (
            .O(N__39722),
            .I(N__39716));
    LocalMux I__8366 (
            .O(N__39719),
            .I(wdtick_cnt_2));
    LocalMux I__8365 (
            .O(N__39716),
            .I(wdtick_cnt_2));
    InMux I__8364 (
            .O(N__39711),
            .I(n19933));
    InMux I__8363 (
            .O(N__39708),
            .I(N__39704));
    InMux I__8362 (
            .O(N__39707),
            .I(N__39701));
    LocalMux I__8361 (
            .O(N__39704),
            .I(wdtick_cnt_3));
    LocalMux I__8360 (
            .O(N__39701),
            .I(wdtick_cnt_3));
    InMux I__8359 (
            .O(N__39696),
            .I(n19934));
    InMux I__8358 (
            .O(N__39693),
            .I(N__39689));
    InMux I__8357 (
            .O(N__39692),
            .I(N__39686));
    LocalMux I__8356 (
            .O(N__39689),
            .I(wdtick_cnt_4));
    LocalMux I__8355 (
            .O(N__39686),
            .I(wdtick_cnt_4));
    InMux I__8354 (
            .O(N__39681),
            .I(n19935));
    InMux I__8353 (
            .O(N__39678),
            .I(N__39674));
    InMux I__8352 (
            .O(N__39677),
            .I(N__39671));
    LocalMux I__8351 (
            .O(N__39674),
            .I(wdtick_cnt_5));
    LocalMux I__8350 (
            .O(N__39671),
            .I(wdtick_cnt_5));
    InMux I__8349 (
            .O(N__39666),
            .I(n19936));
    InMux I__8348 (
            .O(N__39663),
            .I(N__39659));
    InMux I__8347 (
            .O(N__39662),
            .I(N__39656));
    LocalMux I__8346 (
            .O(N__39659),
            .I(N__39653));
    LocalMux I__8345 (
            .O(N__39656),
            .I(N__39650));
    Span4Mux_v I__8344 (
            .O(N__39653),
            .I(N__39646));
    Span4Mux_h I__8343 (
            .O(N__39650),
            .I(N__39643));
    InMux I__8342 (
            .O(N__39649),
            .I(N__39636));
    Span4Mux_h I__8341 (
            .O(N__39646),
            .I(N__39631));
    Span4Mux_v I__8340 (
            .O(N__39643),
            .I(N__39631));
    InMux I__8339 (
            .O(N__39642),
            .I(N__39628));
    InMux I__8338 (
            .O(N__39641),
            .I(N__39625));
    InMux I__8337 (
            .O(N__39640),
            .I(N__39622));
    InMux I__8336 (
            .O(N__39639),
            .I(N__39619));
    LocalMux I__8335 (
            .O(N__39636),
            .I(N__39616));
    Span4Mux_v I__8334 (
            .O(N__39631),
            .I(N__39613));
    LocalMux I__8333 (
            .O(N__39628),
            .I(n12624));
    LocalMux I__8332 (
            .O(N__39625),
            .I(n12624));
    LocalMux I__8331 (
            .O(N__39622),
            .I(n12624));
    LocalMux I__8330 (
            .O(N__39619),
            .I(n12624));
    Odrv12 I__8329 (
            .O(N__39616),
            .I(n12624));
    Odrv4 I__8328 (
            .O(N__39613),
            .I(n12624));
    CascadeMux I__8327 (
            .O(N__39600),
            .I(N__39597));
    InMux I__8326 (
            .O(N__39597),
            .I(N__39592));
    InMux I__8325 (
            .O(N__39596),
            .I(N__39589));
    CascadeMux I__8324 (
            .O(N__39595),
            .I(N__39586));
    LocalMux I__8323 (
            .O(N__39592),
            .I(N__39582));
    LocalMux I__8322 (
            .O(N__39589),
            .I(N__39579));
    InMux I__8321 (
            .O(N__39586),
            .I(N__39574));
    InMux I__8320 (
            .O(N__39585),
            .I(N__39574));
    Span4Mux_v I__8319 (
            .O(N__39582),
            .I(N__39567));
    Span4Mux_v I__8318 (
            .O(N__39579),
            .I(N__39567));
    LocalMux I__8317 (
            .O(N__39574),
            .I(N__39567));
    Span4Mux_h I__8316 (
            .O(N__39567),
            .I(N__39564));
    Span4Mux_v I__8315 (
            .O(N__39564),
            .I(N__39560));
    CascadeMux I__8314 (
            .O(N__39563),
            .I(N__39557));
    Span4Mux_v I__8313 (
            .O(N__39560),
            .I(N__39554));
    InMux I__8312 (
            .O(N__39557),
            .I(N__39551));
    Span4Mux_h I__8311 (
            .O(N__39554),
            .I(N__39548));
    LocalMux I__8310 (
            .O(N__39551),
            .I(buf_cfgRTD_1));
    Odrv4 I__8309 (
            .O(N__39548),
            .I(buf_cfgRTD_1));
    InMux I__8308 (
            .O(N__39543),
            .I(N__39540));
    LocalMux I__8307 (
            .O(N__39540),
            .I(N__39535));
    InMux I__8306 (
            .O(N__39539),
            .I(N__39532));
    InMux I__8305 (
            .O(N__39538),
            .I(N__39529));
    Span4Mux_v I__8304 (
            .O(N__39535),
            .I(N__39525));
    LocalMux I__8303 (
            .O(N__39532),
            .I(N__39520));
    LocalMux I__8302 (
            .O(N__39529),
            .I(N__39520));
    InMux I__8301 (
            .O(N__39528),
            .I(N__39517));
    Span4Mux_h I__8300 (
            .O(N__39525),
            .I(N__39509));
    Span4Mux_v I__8299 (
            .O(N__39520),
            .I(N__39509));
    LocalMux I__8298 (
            .O(N__39517),
            .I(N__39506));
    InMux I__8297 (
            .O(N__39516),
            .I(N__39503));
    InMux I__8296 (
            .O(N__39515),
            .I(N__39498));
    InMux I__8295 (
            .O(N__39514),
            .I(N__39498));
    Span4Mux_v I__8294 (
            .O(N__39509),
            .I(N__39495));
    Span4Mux_h I__8293 (
            .O(N__39506),
            .I(N__39490));
    LocalMux I__8292 (
            .O(N__39503),
            .I(N__39490));
    LocalMux I__8291 (
            .O(N__39498),
            .I(N__39487));
    Sp12to4 I__8290 (
            .O(N__39495),
            .I(N__39484));
    Span4Mux_v I__8289 (
            .O(N__39490),
            .I(N__39479));
    Span4Mux_h I__8288 (
            .O(N__39487),
            .I(N__39479));
    Odrv12 I__8287 (
            .O(N__39484),
            .I(n12610));
    Odrv4 I__8286 (
            .O(N__39479),
            .I(n12610));
    IoInMux I__8285 (
            .O(N__39474),
            .I(N__39471));
    LocalMux I__8284 (
            .O(N__39471),
            .I(N__39468));
    Span4Mux_s0_v I__8283 (
            .O(N__39468),
            .I(N__39465));
    Span4Mux_v I__8282 (
            .O(N__39465),
            .I(N__39462));
    Span4Mux_v I__8281 (
            .O(N__39462),
            .I(N__39457));
    InMux I__8280 (
            .O(N__39461),
            .I(N__39454));
    InMux I__8279 (
            .O(N__39460),
            .I(N__39451));
    Odrv4 I__8278 (
            .O(N__39457),
            .I(IAC_OSR0));
    LocalMux I__8277 (
            .O(N__39454),
            .I(IAC_OSR0));
    LocalMux I__8276 (
            .O(N__39451),
            .I(IAC_OSR0));
    CascadeMux I__8275 (
            .O(N__39444),
            .I(N__39441));
    CascadeBuf I__8274 (
            .O(N__39441),
            .I(N__39438));
    CascadeMux I__8273 (
            .O(N__39438),
            .I(N__39435));
    CascadeBuf I__8272 (
            .O(N__39435),
            .I(N__39432));
    CascadeMux I__8271 (
            .O(N__39432),
            .I(N__39429));
    CascadeBuf I__8270 (
            .O(N__39429),
            .I(N__39426));
    CascadeMux I__8269 (
            .O(N__39426),
            .I(N__39423));
    CascadeBuf I__8268 (
            .O(N__39423),
            .I(N__39420));
    CascadeMux I__8267 (
            .O(N__39420),
            .I(N__39417));
    CascadeBuf I__8266 (
            .O(N__39417),
            .I(N__39414));
    CascadeMux I__8265 (
            .O(N__39414),
            .I(N__39411));
    CascadeBuf I__8264 (
            .O(N__39411),
            .I(N__39408));
    CascadeMux I__8263 (
            .O(N__39408),
            .I(N__39405));
    CascadeBuf I__8262 (
            .O(N__39405),
            .I(N__39402));
    CascadeMux I__8261 (
            .O(N__39402),
            .I(N__39398));
    CascadeMux I__8260 (
            .O(N__39401),
            .I(N__39395));
    CascadeBuf I__8259 (
            .O(N__39398),
            .I(N__39392));
    CascadeBuf I__8258 (
            .O(N__39395),
            .I(N__39389));
    CascadeMux I__8257 (
            .O(N__39392),
            .I(N__39386));
    CascadeMux I__8256 (
            .O(N__39389),
            .I(N__39383));
    CascadeBuf I__8255 (
            .O(N__39386),
            .I(N__39380));
    InMux I__8254 (
            .O(N__39383),
            .I(N__39377));
    CascadeMux I__8253 (
            .O(N__39380),
            .I(N__39374));
    LocalMux I__8252 (
            .O(N__39377),
            .I(N__39371));
    InMux I__8251 (
            .O(N__39374),
            .I(N__39368));
    Span12Mux_h I__8250 (
            .O(N__39371),
            .I(N__39365));
    LocalMux I__8249 (
            .O(N__39368),
            .I(N__39362));
    Odrv12 I__8248 (
            .O(N__39365),
            .I(data_index_9_N_212_8));
    Odrv12 I__8247 (
            .O(N__39362),
            .I(data_index_9_N_212_8));
    InMux I__8246 (
            .O(N__39357),
            .I(N__39352));
    InMux I__8245 (
            .O(N__39356),
            .I(N__39349));
    InMux I__8244 (
            .O(N__39355),
            .I(N__39346));
    LocalMux I__8243 (
            .O(N__39352),
            .I(N__39341));
    LocalMux I__8242 (
            .O(N__39349),
            .I(N__39341));
    LocalMux I__8241 (
            .O(N__39346),
            .I(data_index_1));
    Odrv4 I__8240 (
            .O(N__39341),
            .I(data_index_1));
    InMux I__8239 (
            .O(N__39336),
            .I(N__39333));
    LocalMux I__8238 (
            .O(N__39333),
            .I(n8_adj_1570));
    CascadeMux I__8237 (
            .O(N__39330),
            .I(n8_adj_1570_cascade_));
    InMux I__8236 (
            .O(N__39327),
            .I(N__39323));
    InMux I__8235 (
            .O(N__39326),
            .I(N__39320));
    LocalMux I__8234 (
            .O(N__39323),
            .I(N__39315));
    LocalMux I__8233 (
            .O(N__39320),
            .I(N__39315));
    Odrv12 I__8232 (
            .O(N__39315),
            .I(n7_adj_1569));
    CascadeMux I__8231 (
            .O(N__39312),
            .I(N__39309));
    CascadeBuf I__8230 (
            .O(N__39309),
            .I(N__39306));
    CascadeMux I__8229 (
            .O(N__39306),
            .I(N__39303));
    CascadeBuf I__8228 (
            .O(N__39303),
            .I(N__39300));
    CascadeMux I__8227 (
            .O(N__39300),
            .I(N__39297));
    CascadeBuf I__8226 (
            .O(N__39297),
            .I(N__39294));
    CascadeMux I__8225 (
            .O(N__39294),
            .I(N__39291));
    CascadeBuf I__8224 (
            .O(N__39291),
            .I(N__39288));
    CascadeMux I__8223 (
            .O(N__39288),
            .I(N__39285));
    CascadeBuf I__8222 (
            .O(N__39285),
            .I(N__39282));
    CascadeMux I__8221 (
            .O(N__39282),
            .I(N__39279));
    CascadeBuf I__8220 (
            .O(N__39279),
            .I(N__39276));
    CascadeMux I__8219 (
            .O(N__39276),
            .I(N__39273));
    CascadeBuf I__8218 (
            .O(N__39273),
            .I(N__39269));
    CascadeMux I__8217 (
            .O(N__39272),
            .I(N__39266));
    CascadeMux I__8216 (
            .O(N__39269),
            .I(N__39263));
    CascadeBuf I__8215 (
            .O(N__39266),
            .I(N__39260));
    CascadeBuf I__8214 (
            .O(N__39263),
            .I(N__39257));
    CascadeMux I__8213 (
            .O(N__39260),
            .I(N__39254));
    CascadeMux I__8212 (
            .O(N__39257),
            .I(N__39251));
    InMux I__8211 (
            .O(N__39254),
            .I(N__39248));
    CascadeBuf I__8210 (
            .O(N__39251),
            .I(N__39245));
    LocalMux I__8209 (
            .O(N__39248),
            .I(N__39242));
    CascadeMux I__8208 (
            .O(N__39245),
            .I(N__39239));
    Span12Mux_s9_h I__8207 (
            .O(N__39242),
            .I(N__39236));
    InMux I__8206 (
            .O(N__39239),
            .I(N__39233));
    Span12Mux_v I__8205 (
            .O(N__39236),
            .I(N__39230));
    LocalMux I__8204 (
            .O(N__39233),
            .I(N__39227));
    Odrv12 I__8203 (
            .O(N__39230),
            .I(data_index_9_N_212_1));
    Odrv12 I__8202 (
            .O(N__39227),
            .I(data_index_9_N_212_1));
    InMux I__8201 (
            .O(N__39222),
            .I(N__39218));
    InMux I__8200 (
            .O(N__39221),
            .I(N__39215));
    LocalMux I__8199 (
            .O(N__39218),
            .I(N__39209));
    LocalMux I__8198 (
            .O(N__39215),
            .I(N__39209));
    InMux I__8197 (
            .O(N__39214),
            .I(N__39206));
    Span4Mux_h I__8196 (
            .O(N__39209),
            .I(N__39203));
    LocalMux I__8195 (
            .O(N__39206),
            .I(data_index_2));
    Odrv4 I__8194 (
            .O(N__39203),
            .I(data_index_2));
    InMux I__8193 (
            .O(N__39198),
            .I(N__39192));
    InMux I__8192 (
            .O(N__39197),
            .I(N__39192));
    LocalMux I__8191 (
            .O(N__39192),
            .I(n8_adj_1558));
    InMux I__8190 (
            .O(N__39189),
            .I(N__39183));
    InMux I__8189 (
            .O(N__39188),
            .I(N__39183));
    LocalMux I__8188 (
            .O(N__39183),
            .I(N__39180));
    Odrv12 I__8187 (
            .O(N__39180),
            .I(n7_adj_1557));
    InMux I__8186 (
            .O(N__39177),
            .I(N__39173));
    InMux I__8185 (
            .O(N__39176),
            .I(N__39170));
    LocalMux I__8184 (
            .O(N__39173),
            .I(N__39166));
    LocalMux I__8183 (
            .O(N__39170),
            .I(N__39163));
    InMux I__8182 (
            .O(N__39169),
            .I(N__39160));
    Span4Mux_v I__8181 (
            .O(N__39166),
            .I(N__39155));
    Span4Mux_h I__8180 (
            .O(N__39163),
            .I(N__39155));
    LocalMux I__8179 (
            .O(N__39160),
            .I(data_index_8));
    Odrv4 I__8178 (
            .O(N__39155),
            .I(data_index_8));
    CascadeMux I__8177 (
            .O(N__39150),
            .I(N__39147));
    InMux I__8176 (
            .O(N__39147),
            .I(N__39144));
    LocalMux I__8175 (
            .O(N__39144),
            .I(N__39139));
    InMux I__8174 (
            .O(N__39143),
            .I(N__39136));
    CascadeMux I__8173 (
            .O(N__39142),
            .I(N__39133));
    Span4Mux_h I__8172 (
            .O(N__39139),
            .I(N__39130));
    LocalMux I__8171 (
            .O(N__39136),
            .I(N__39127));
    InMux I__8170 (
            .O(N__39133),
            .I(N__39124));
    Span4Mux_h I__8169 (
            .O(N__39130),
            .I(N__39121));
    Span12Mux_v I__8168 (
            .O(N__39127),
            .I(N__39118));
    LocalMux I__8167 (
            .O(N__39124),
            .I(buf_adcdata_iac_16));
    Odrv4 I__8166 (
            .O(N__39121),
            .I(buf_adcdata_iac_16));
    Odrv12 I__8165 (
            .O(N__39118),
            .I(buf_adcdata_iac_16));
    InMux I__8164 (
            .O(N__39111),
            .I(N__39108));
    LocalMux I__8163 (
            .O(N__39108),
            .I(N__39105));
    Span4Mux_v I__8162 (
            .O(N__39105),
            .I(N__39100));
    InMux I__8161 (
            .O(N__39104),
            .I(N__39097));
    InMux I__8160 (
            .O(N__39103),
            .I(N__39094));
    Span4Mux_h I__8159 (
            .O(N__39100),
            .I(N__39091));
    LocalMux I__8158 (
            .O(N__39097),
            .I(buf_dds1_8));
    LocalMux I__8157 (
            .O(N__39094),
            .I(buf_dds1_8));
    Odrv4 I__8156 (
            .O(N__39091),
            .I(buf_dds1_8));
    CascadeMux I__8155 (
            .O(N__39084),
            .I(n22389_cascade_));
    CascadeMux I__8154 (
            .O(N__39081),
            .I(N__39078));
    InMux I__8153 (
            .O(N__39078),
            .I(N__39073));
    InMux I__8152 (
            .O(N__39077),
            .I(N__39070));
    InMux I__8151 (
            .O(N__39076),
            .I(N__39067));
    LocalMux I__8150 (
            .O(N__39073),
            .I(N__39062));
    LocalMux I__8149 (
            .O(N__39070),
            .I(N__39062));
    LocalMux I__8148 (
            .O(N__39067),
            .I(buf_dds0_8));
    Odrv4 I__8147 (
            .O(N__39062),
            .I(buf_dds0_8));
    InMux I__8146 (
            .O(N__39057),
            .I(N__39052));
    InMux I__8145 (
            .O(N__39056),
            .I(N__39049));
    InMux I__8144 (
            .O(N__39055),
            .I(N__39046));
    LocalMux I__8143 (
            .O(N__39052),
            .I(N__39041));
    LocalMux I__8142 (
            .O(N__39049),
            .I(N__39041));
    LocalMux I__8141 (
            .O(N__39046),
            .I(data_index_5));
    Odrv4 I__8140 (
            .O(N__39041),
            .I(data_index_5));
    IoInMux I__8139 (
            .O(N__39036),
            .I(N__39033));
    LocalMux I__8138 (
            .O(N__39033),
            .I(N__39030));
    Span4Mux_s0_v I__8137 (
            .O(N__39030),
            .I(N__39027));
    Sp12to4 I__8136 (
            .O(N__39027),
            .I(N__39023));
    CascadeMux I__8135 (
            .O(N__39026),
            .I(N__39020));
    Span12Mux_h I__8134 (
            .O(N__39023),
            .I(N__39017));
    InMux I__8133 (
            .O(N__39020),
            .I(N__39014));
    Odrv12 I__8132 (
            .O(N__39017),
            .I(DDS_SCK));
    LocalMux I__8131 (
            .O(N__39014),
            .I(DDS_SCK));
    InMux I__8130 (
            .O(N__39009),
            .I(N__39006));
    LocalMux I__8129 (
            .O(N__39006),
            .I(N__39002));
    CascadeMux I__8128 (
            .O(N__39005),
            .I(N__38999));
    Span4Mux_v I__8127 (
            .O(N__39002),
            .I(N__38996));
    InMux I__8126 (
            .O(N__38999),
            .I(N__38993));
    Span4Mux_h I__8125 (
            .O(N__38996),
            .I(N__38988));
    LocalMux I__8124 (
            .O(N__38993),
            .I(N__38988));
    Odrv4 I__8123 (
            .O(N__38988),
            .I(tmp_buf_15));
    IoInMux I__8122 (
            .O(N__38985),
            .I(N__38982));
    LocalMux I__8121 (
            .O(N__38982),
            .I(N__38979));
    Span12Mux_s11_v I__8120 (
            .O(N__38979),
            .I(N__38976));
    Span12Mux_h I__8119 (
            .O(N__38976),
            .I(N__38972));
    InMux I__8118 (
            .O(N__38975),
            .I(N__38969));
    Odrv12 I__8117 (
            .O(N__38972),
            .I(DDS_MOSI));
    LocalMux I__8116 (
            .O(N__38969),
            .I(DDS_MOSI));
    InMux I__8115 (
            .O(N__38964),
            .I(N__38959));
    InMux I__8114 (
            .O(N__38963),
            .I(N__38956));
    InMux I__8113 (
            .O(N__38962),
            .I(N__38953));
    LocalMux I__8112 (
            .O(N__38959),
            .I(data_index_9));
    LocalMux I__8111 (
            .O(N__38956),
            .I(data_index_9));
    LocalMux I__8110 (
            .O(N__38953),
            .I(data_index_9));
    InMux I__8109 (
            .O(N__38946),
            .I(N__38941));
    CascadeMux I__8108 (
            .O(N__38945),
            .I(N__38938));
    CascadeMux I__8107 (
            .O(N__38944),
            .I(N__38935));
    LocalMux I__8106 (
            .O(N__38941),
            .I(N__38924));
    InMux I__8105 (
            .O(N__38938),
            .I(N__38921));
    InMux I__8104 (
            .O(N__38935),
            .I(N__38918));
    CascadeMux I__8103 (
            .O(N__38934),
            .I(N__38915));
    CascadeMux I__8102 (
            .O(N__38933),
            .I(N__38912));
    CascadeMux I__8101 (
            .O(N__38932),
            .I(N__38909));
    CascadeMux I__8100 (
            .O(N__38931),
            .I(N__38906));
    CascadeMux I__8099 (
            .O(N__38930),
            .I(N__38903));
    CascadeMux I__8098 (
            .O(N__38929),
            .I(N__38900));
    CascadeMux I__8097 (
            .O(N__38928),
            .I(N__38897));
    CascadeMux I__8096 (
            .O(N__38927),
            .I(N__38894));
    Span4Mux_h I__8095 (
            .O(N__38924),
            .I(N__38891));
    LocalMux I__8094 (
            .O(N__38921),
            .I(N__38886));
    LocalMux I__8093 (
            .O(N__38918),
            .I(N__38886));
    InMux I__8092 (
            .O(N__38915),
            .I(N__38877));
    InMux I__8091 (
            .O(N__38912),
            .I(N__38877));
    InMux I__8090 (
            .O(N__38909),
            .I(N__38877));
    InMux I__8089 (
            .O(N__38906),
            .I(N__38877));
    InMux I__8088 (
            .O(N__38903),
            .I(N__38868));
    InMux I__8087 (
            .O(N__38900),
            .I(N__38868));
    InMux I__8086 (
            .O(N__38897),
            .I(N__38868));
    InMux I__8085 (
            .O(N__38894),
            .I(N__38868));
    Odrv4 I__8084 (
            .O(N__38891),
            .I(n10756));
    Odrv4 I__8083 (
            .O(N__38886),
            .I(n10756));
    LocalMux I__8082 (
            .O(N__38877),
            .I(n10756));
    LocalMux I__8081 (
            .O(N__38868),
            .I(n10756));
    InMux I__8080 (
            .O(N__38859),
            .I(n19812));
    InMux I__8079 (
            .O(N__38856),
            .I(N__38853));
    LocalMux I__8078 (
            .O(N__38853),
            .I(N__38850));
    Span4Mux_v I__8077 (
            .O(N__38850),
            .I(N__38847));
    Span4Mux_h I__8076 (
            .O(N__38847),
            .I(N__38844));
    Span4Mux_h I__8075 (
            .O(N__38844),
            .I(N__38841));
    Span4Mux_v I__8074 (
            .O(N__38841),
            .I(N__38838));
    Odrv4 I__8073 (
            .O(N__38838),
            .I(buf_data_iac_1));
    InMux I__8072 (
            .O(N__38835),
            .I(N__38832));
    LocalMux I__8071 (
            .O(N__38832),
            .I(n22_adj_1617));
    CascadeMux I__8070 (
            .O(N__38829),
            .I(N__38825));
    CascadeMux I__8069 (
            .O(N__38828),
            .I(N__38821));
    InMux I__8068 (
            .O(N__38825),
            .I(N__38814));
    InMux I__8067 (
            .O(N__38824),
            .I(N__38814));
    InMux I__8066 (
            .O(N__38821),
            .I(N__38814));
    LocalMux I__8065 (
            .O(N__38814),
            .I(N__38811));
    Span4Mux_h I__8064 (
            .O(N__38811),
            .I(N__38807));
    CascadeMux I__8063 (
            .O(N__38810),
            .I(N__38804));
    Span4Mux_v I__8062 (
            .O(N__38807),
            .I(N__38801));
    InMux I__8061 (
            .O(N__38804),
            .I(N__38798));
    Sp12to4 I__8060 (
            .O(N__38801),
            .I(N__38795));
    LocalMux I__8059 (
            .O(N__38798),
            .I(trig_dds1));
    Odrv12 I__8058 (
            .O(N__38795),
            .I(trig_dds1));
    InMux I__8057 (
            .O(N__38790),
            .I(N__38785));
    InMux I__8056 (
            .O(N__38789),
            .I(N__38780));
    InMux I__8055 (
            .O(N__38788),
            .I(N__38780));
    LocalMux I__8054 (
            .O(N__38785),
            .I(buf_dds0_7));
    LocalMux I__8053 (
            .O(N__38780),
            .I(buf_dds0_7));
    InMux I__8052 (
            .O(N__38775),
            .I(N__38765));
    InMux I__8051 (
            .O(N__38774),
            .I(N__38765));
    InMux I__8050 (
            .O(N__38773),
            .I(N__38759));
    InMux I__8049 (
            .O(N__38772),
            .I(N__38754));
    InMux I__8048 (
            .O(N__38771),
            .I(N__38754));
    CascadeMux I__8047 (
            .O(N__38770),
            .I(N__38739));
    LocalMux I__8046 (
            .O(N__38765),
            .I(N__38734));
    InMux I__8045 (
            .O(N__38764),
            .I(N__38731));
    InMux I__8044 (
            .O(N__38763),
            .I(N__38728));
    InMux I__8043 (
            .O(N__38762),
            .I(N__38725));
    LocalMux I__8042 (
            .O(N__38759),
            .I(N__38722));
    LocalMux I__8041 (
            .O(N__38754),
            .I(N__38719));
    InMux I__8040 (
            .O(N__38753),
            .I(N__38712));
    InMux I__8039 (
            .O(N__38752),
            .I(N__38712));
    InMux I__8038 (
            .O(N__38751),
            .I(N__38712));
    InMux I__8037 (
            .O(N__38750),
            .I(N__38709));
    InMux I__8036 (
            .O(N__38749),
            .I(N__38706));
    InMux I__8035 (
            .O(N__38748),
            .I(N__38701));
    InMux I__8034 (
            .O(N__38747),
            .I(N__38701));
    InMux I__8033 (
            .O(N__38746),
            .I(N__38696));
    InMux I__8032 (
            .O(N__38745),
            .I(N__38696));
    InMux I__8031 (
            .O(N__38744),
            .I(N__38693));
    InMux I__8030 (
            .O(N__38743),
            .I(N__38688));
    InMux I__8029 (
            .O(N__38742),
            .I(N__38688));
    InMux I__8028 (
            .O(N__38739),
            .I(N__38685));
    InMux I__8027 (
            .O(N__38738),
            .I(N__38680));
    InMux I__8026 (
            .O(N__38737),
            .I(N__38680));
    Span4Mux_h I__8025 (
            .O(N__38734),
            .I(N__38673));
    LocalMux I__8024 (
            .O(N__38731),
            .I(N__38673));
    LocalMux I__8023 (
            .O(N__38728),
            .I(N__38673));
    LocalMux I__8022 (
            .O(N__38725),
            .I(N__38670));
    Span4Mux_h I__8021 (
            .O(N__38722),
            .I(N__38665));
    Span4Mux_h I__8020 (
            .O(N__38719),
            .I(N__38665));
    LocalMux I__8019 (
            .O(N__38712),
            .I(N__38662));
    LocalMux I__8018 (
            .O(N__38709),
            .I(N__38659));
    LocalMux I__8017 (
            .O(N__38706),
            .I(N__38654));
    LocalMux I__8016 (
            .O(N__38701),
            .I(N__38654));
    LocalMux I__8015 (
            .O(N__38696),
            .I(N__38651));
    LocalMux I__8014 (
            .O(N__38693),
            .I(N__38644));
    LocalMux I__8013 (
            .O(N__38688),
            .I(N__38644));
    LocalMux I__8012 (
            .O(N__38685),
            .I(N__38644));
    LocalMux I__8011 (
            .O(N__38680),
            .I(N__38641));
    Span4Mux_v I__8010 (
            .O(N__38673),
            .I(N__38635));
    Span4Mux_h I__8009 (
            .O(N__38670),
            .I(N__38635));
    Span4Mux_h I__8008 (
            .O(N__38665),
            .I(N__38628));
    Span4Mux_v I__8007 (
            .O(N__38662),
            .I(N__38628));
    Span4Mux_h I__8006 (
            .O(N__38659),
            .I(N__38628));
    Span4Mux_h I__8005 (
            .O(N__38654),
            .I(N__38619));
    Span4Mux_v I__8004 (
            .O(N__38651),
            .I(N__38619));
    Span4Mux_v I__8003 (
            .O(N__38644),
            .I(N__38619));
    Span4Mux_h I__8002 (
            .O(N__38641),
            .I(N__38619));
    InMux I__8001 (
            .O(N__38640),
            .I(N__38616));
    Odrv4 I__8000 (
            .O(N__38635),
            .I(n21079));
    Odrv4 I__7999 (
            .O(N__38628),
            .I(n21079));
    Odrv4 I__7998 (
            .O(N__38619),
            .I(n21079));
    LocalMux I__7997 (
            .O(N__38616),
            .I(n21079));
    CascadeMux I__7996 (
            .O(N__38607),
            .I(N__38603));
    InMux I__7995 (
            .O(N__38606),
            .I(N__38579));
    InMux I__7994 (
            .O(N__38603),
            .I(N__38574));
    InMux I__7993 (
            .O(N__38602),
            .I(N__38574));
    InMux I__7992 (
            .O(N__38601),
            .I(N__38571));
    InMux I__7991 (
            .O(N__38600),
            .I(N__38565));
    InMux I__7990 (
            .O(N__38599),
            .I(N__38565));
    InMux I__7989 (
            .O(N__38598),
            .I(N__38554));
    InMux I__7988 (
            .O(N__38597),
            .I(N__38544));
    InMux I__7987 (
            .O(N__38596),
            .I(N__38544));
    InMux I__7986 (
            .O(N__38595),
            .I(N__38544));
    InMux I__7985 (
            .O(N__38594),
            .I(N__38533));
    InMux I__7984 (
            .O(N__38593),
            .I(N__38533));
    InMux I__7983 (
            .O(N__38592),
            .I(N__38533));
    InMux I__7982 (
            .O(N__38591),
            .I(N__38533));
    InMux I__7981 (
            .O(N__38590),
            .I(N__38533));
    InMux I__7980 (
            .O(N__38589),
            .I(N__38528));
    InMux I__7979 (
            .O(N__38588),
            .I(N__38528));
    InMux I__7978 (
            .O(N__38587),
            .I(N__38515));
    InMux I__7977 (
            .O(N__38586),
            .I(N__38515));
    InMux I__7976 (
            .O(N__38585),
            .I(N__38515));
    InMux I__7975 (
            .O(N__38584),
            .I(N__38515));
    InMux I__7974 (
            .O(N__38583),
            .I(N__38515));
    InMux I__7973 (
            .O(N__38582),
            .I(N__38515));
    LocalMux I__7972 (
            .O(N__38579),
            .I(N__38510));
    LocalMux I__7971 (
            .O(N__38574),
            .I(N__38510));
    LocalMux I__7970 (
            .O(N__38571),
            .I(N__38507));
    InMux I__7969 (
            .O(N__38570),
            .I(N__38497));
    LocalMux I__7968 (
            .O(N__38565),
            .I(N__38494));
    CascadeMux I__7967 (
            .O(N__38564),
            .I(N__38491));
    InMux I__7966 (
            .O(N__38563),
            .I(N__38488));
    InMux I__7965 (
            .O(N__38562),
            .I(N__38481));
    InMux I__7964 (
            .O(N__38561),
            .I(N__38481));
    InMux I__7963 (
            .O(N__38560),
            .I(N__38481));
    InMux I__7962 (
            .O(N__38559),
            .I(N__38474));
    InMux I__7961 (
            .O(N__38558),
            .I(N__38474));
    InMux I__7960 (
            .O(N__38557),
            .I(N__38474));
    LocalMux I__7959 (
            .O(N__38554),
            .I(N__38471));
    InMux I__7958 (
            .O(N__38553),
            .I(N__38468));
    InMux I__7957 (
            .O(N__38552),
            .I(N__38463));
    InMux I__7956 (
            .O(N__38551),
            .I(N__38463));
    LocalMux I__7955 (
            .O(N__38544),
            .I(N__38460));
    LocalMux I__7954 (
            .O(N__38533),
            .I(N__38443));
    LocalMux I__7953 (
            .O(N__38528),
            .I(N__38438));
    LocalMux I__7952 (
            .O(N__38515),
            .I(N__38438));
    Span4Mux_v I__7951 (
            .O(N__38510),
            .I(N__38435));
    Span4Mux_v I__7950 (
            .O(N__38507),
            .I(N__38432));
    InMux I__7949 (
            .O(N__38506),
            .I(N__38427));
    InMux I__7948 (
            .O(N__38505),
            .I(N__38427));
    InMux I__7947 (
            .O(N__38504),
            .I(N__38422));
    InMux I__7946 (
            .O(N__38503),
            .I(N__38422));
    InMux I__7945 (
            .O(N__38502),
            .I(N__38415));
    InMux I__7944 (
            .O(N__38501),
            .I(N__38415));
    InMux I__7943 (
            .O(N__38500),
            .I(N__38415));
    LocalMux I__7942 (
            .O(N__38497),
            .I(N__38412));
    Span4Mux_v I__7941 (
            .O(N__38494),
            .I(N__38409));
    InMux I__7940 (
            .O(N__38491),
            .I(N__38394));
    LocalMux I__7939 (
            .O(N__38488),
            .I(N__38385));
    LocalMux I__7938 (
            .O(N__38481),
            .I(N__38385));
    LocalMux I__7937 (
            .O(N__38474),
            .I(N__38385));
    Span4Mux_h I__7936 (
            .O(N__38471),
            .I(N__38385));
    LocalMux I__7935 (
            .O(N__38468),
            .I(N__38378));
    LocalMux I__7934 (
            .O(N__38463),
            .I(N__38378));
    Span4Mux_v I__7933 (
            .O(N__38460),
            .I(N__38378));
    InMux I__7932 (
            .O(N__38459),
            .I(N__38371));
    InMux I__7931 (
            .O(N__38458),
            .I(N__38371));
    InMux I__7930 (
            .O(N__38457),
            .I(N__38371));
    InMux I__7929 (
            .O(N__38456),
            .I(N__38364));
    InMux I__7928 (
            .O(N__38455),
            .I(N__38364));
    InMux I__7927 (
            .O(N__38454),
            .I(N__38364));
    InMux I__7926 (
            .O(N__38453),
            .I(N__38353));
    InMux I__7925 (
            .O(N__38452),
            .I(N__38353));
    InMux I__7924 (
            .O(N__38451),
            .I(N__38353));
    InMux I__7923 (
            .O(N__38450),
            .I(N__38353));
    InMux I__7922 (
            .O(N__38449),
            .I(N__38353));
    InMux I__7921 (
            .O(N__38448),
            .I(N__38348));
    InMux I__7920 (
            .O(N__38447),
            .I(N__38348));
    InMux I__7919 (
            .O(N__38446),
            .I(N__38345));
    Sp12to4 I__7918 (
            .O(N__38443),
            .I(N__38342));
    Span4Mux_v I__7917 (
            .O(N__38438),
            .I(N__38335));
    Span4Mux_v I__7916 (
            .O(N__38435),
            .I(N__38335));
    Span4Mux_h I__7915 (
            .O(N__38432),
            .I(N__38335));
    LocalMux I__7914 (
            .O(N__38427),
            .I(N__38324));
    LocalMux I__7913 (
            .O(N__38422),
            .I(N__38324));
    LocalMux I__7912 (
            .O(N__38415),
            .I(N__38324));
    Sp12to4 I__7911 (
            .O(N__38412),
            .I(N__38324));
    Sp12to4 I__7910 (
            .O(N__38409),
            .I(N__38324));
    InMux I__7909 (
            .O(N__38408),
            .I(N__38317));
    InMux I__7908 (
            .O(N__38407),
            .I(N__38317));
    InMux I__7907 (
            .O(N__38406),
            .I(N__38317));
    InMux I__7906 (
            .O(N__38405),
            .I(N__38308));
    InMux I__7905 (
            .O(N__38404),
            .I(N__38308));
    InMux I__7904 (
            .O(N__38403),
            .I(N__38308));
    InMux I__7903 (
            .O(N__38402),
            .I(N__38308));
    InMux I__7902 (
            .O(N__38401),
            .I(N__38297));
    InMux I__7901 (
            .O(N__38400),
            .I(N__38297));
    InMux I__7900 (
            .O(N__38399),
            .I(N__38297));
    InMux I__7899 (
            .O(N__38398),
            .I(N__38297));
    InMux I__7898 (
            .O(N__38397),
            .I(N__38297));
    LocalMux I__7897 (
            .O(N__38394),
            .I(N__38288));
    Span4Mux_v I__7896 (
            .O(N__38385),
            .I(N__38288));
    Span4Mux_h I__7895 (
            .O(N__38378),
            .I(N__38288));
    LocalMux I__7894 (
            .O(N__38371),
            .I(N__38288));
    LocalMux I__7893 (
            .O(N__38364),
            .I(adc_state_0));
    LocalMux I__7892 (
            .O(N__38353),
            .I(adc_state_0));
    LocalMux I__7891 (
            .O(N__38348),
            .I(adc_state_0));
    LocalMux I__7890 (
            .O(N__38345),
            .I(adc_state_0));
    Odrv12 I__7889 (
            .O(N__38342),
            .I(adc_state_0));
    Odrv4 I__7888 (
            .O(N__38335),
            .I(adc_state_0));
    Odrv12 I__7887 (
            .O(N__38324),
            .I(adc_state_0));
    LocalMux I__7886 (
            .O(N__38317),
            .I(adc_state_0));
    LocalMux I__7885 (
            .O(N__38308),
            .I(adc_state_0));
    LocalMux I__7884 (
            .O(N__38297),
            .I(adc_state_0));
    Odrv4 I__7883 (
            .O(N__38288),
            .I(adc_state_0));
    CascadeMux I__7882 (
            .O(N__38265),
            .I(N__38260));
    CascadeMux I__7881 (
            .O(N__38264),
            .I(N__38257));
    InMux I__7880 (
            .O(N__38263),
            .I(N__38254));
    InMux I__7879 (
            .O(N__38260),
            .I(N__38251));
    InMux I__7878 (
            .O(N__38257),
            .I(N__38248));
    LocalMux I__7877 (
            .O(N__38254),
            .I(N__38245));
    LocalMux I__7876 (
            .O(N__38251),
            .I(cmd_rdadctmp_18));
    LocalMux I__7875 (
            .O(N__38248),
            .I(cmd_rdadctmp_18));
    Odrv12 I__7874 (
            .O(N__38245),
            .I(cmd_rdadctmp_18));
    InMux I__7873 (
            .O(N__38238),
            .I(N__38233));
    InMux I__7872 (
            .O(N__38237),
            .I(N__38230));
    CascadeMux I__7871 (
            .O(N__38236),
            .I(N__38227));
    LocalMux I__7870 (
            .O(N__38233),
            .I(N__38224));
    LocalMux I__7869 (
            .O(N__38230),
            .I(N__38221));
    InMux I__7868 (
            .O(N__38227),
            .I(N__38218));
    Span4Mux_v I__7867 (
            .O(N__38224),
            .I(N__38215));
    Span12Mux_s9_v I__7866 (
            .O(N__38221),
            .I(N__38212));
    LocalMux I__7865 (
            .O(N__38218),
            .I(buf_adcdata_iac_10));
    Odrv4 I__7864 (
            .O(N__38215),
            .I(buf_adcdata_iac_10));
    Odrv12 I__7863 (
            .O(N__38212),
            .I(buf_adcdata_iac_10));
    InMux I__7862 (
            .O(N__38205),
            .I(N__38202));
    LocalMux I__7861 (
            .O(N__38202),
            .I(n8_adj_1564));
    InMux I__7860 (
            .O(N__38199),
            .I(N__38196));
    LocalMux I__7859 (
            .O(N__38196),
            .I(N__38192));
    InMux I__7858 (
            .O(N__38195),
            .I(N__38189));
    Odrv4 I__7857 (
            .O(N__38192),
            .I(n7_adj_1563));
    LocalMux I__7856 (
            .O(N__38189),
            .I(n7_adj_1563));
    InMux I__7855 (
            .O(N__38184),
            .I(N__38179));
    InMux I__7854 (
            .O(N__38183),
            .I(N__38176));
    InMux I__7853 (
            .O(N__38182),
            .I(N__38173));
    LocalMux I__7852 (
            .O(N__38179),
            .I(N__38168));
    LocalMux I__7851 (
            .O(N__38176),
            .I(N__38168));
    LocalMux I__7850 (
            .O(N__38173),
            .I(data_index_4));
    Odrv4 I__7849 (
            .O(N__38168),
            .I(data_index_4));
    InMux I__7848 (
            .O(N__38163),
            .I(N__38160));
    LocalMux I__7847 (
            .O(N__38160),
            .I(N__38157));
    Span4Mux_v I__7846 (
            .O(N__38157),
            .I(N__38154));
    Odrv4 I__7845 (
            .O(N__38154),
            .I(n11611));
    SRMux I__7844 (
            .O(N__38151),
            .I(N__38146));
    SRMux I__7843 (
            .O(N__38150),
            .I(N__38143));
    SRMux I__7842 (
            .O(N__38149),
            .I(N__38140));
    LocalMux I__7841 (
            .O(N__38146),
            .I(N__38136));
    LocalMux I__7840 (
            .O(N__38143),
            .I(N__38133));
    LocalMux I__7839 (
            .O(N__38140),
            .I(N__38130));
    SRMux I__7838 (
            .O(N__38139),
            .I(N__38127));
    Span4Mux_h I__7837 (
            .O(N__38136),
            .I(N__38124));
    Span4Mux_v I__7836 (
            .O(N__38133),
            .I(N__38121));
    Span4Mux_h I__7835 (
            .O(N__38130),
            .I(N__38118));
    LocalMux I__7834 (
            .O(N__38127),
            .I(N__38115));
    Odrv4 I__7833 (
            .O(N__38124),
            .I(n14907));
    Odrv4 I__7832 (
            .O(N__38121),
            .I(n14907));
    Odrv4 I__7831 (
            .O(N__38118),
            .I(n14907));
    Odrv4 I__7830 (
            .O(N__38115),
            .I(n14907));
    InMux I__7829 (
            .O(N__38106),
            .I(bfn_14_15_0_));
    InMux I__7828 (
            .O(N__38103),
            .I(n19804));
    InMux I__7827 (
            .O(N__38100),
            .I(n19805));
    InMux I__7826 (
            .O(N__38097),
            .I(N__38092));
    InMux I__7825 (
            .O(N__38096),
            .I(N__38089));
    InMux I__7824 (
            .O(N__38095),
            .I(N__38086));
    LocalMux I__7823 (
            .O(N__38092),
            .I(data_index_3));
    LocalMux I__7822 (
            .O(N__38089),
            .I(data_index_3));
    LocalMux I__7821 (
            .O(N__38086),
            .I(data_index_3));
    InMux I__7820 (
            .O(N__38079),
            .I(N__38075));
    InMux I__7819 (
            .O(N__38078),
            .I(N__38072));
    LocalMux I__7818 (
            .O(N__38075),
            .I(n7_adj_1565));
    LocalMux I__7817 (
            .O(N__38072),
            .I(n7_adj_1565));
    InMux I__7816 (
            .O(N__38067),
            .I(n19806));
    InMux I__7815 (
            .O(N__38064),
            .I(n19807));
    InMux I__7814 (
            .O(N__38061),
            .I(n19808));
    InMux I__7813 (
            .O(N__38058),
            .I(N__38054));
    InMux I__7812 (
            .O(N__38057),
            .I(N__38051));
    LocalMux I__7811 (
            .O(N__38054),
            .I(N__38045));
    LocalMux I__7810 (
            .O(N__38051),
            .I(N__38045));
    InMux I__7809 (
            .O(N__38050),
            .I(N__38042));
    Span4Mux_h I__7808 (
            .O(N__38045),
            .I(N__38039));
    LocalMux I__7807 (
            .O(N__38042),
            .I(data_index_6));
    Odrv4 I__7806 (
            .O(N__38039),
            .I(data_index_6));
    CascadeMux I__7805 (
            .O(N__38034),
            .I(N__38030));
    InMux I__7804 (
            .O(N__38033),
            .I(N__38027));
    InMux I__7803 (
            .O(N__38030),
            .I(N__38024));
    LocalMux I__7802 (
            .O(N__38027),
            .I(N__38021));
    LocalMux I__7801 (
            .O(N__38024),
            .I(N__38018));
    Odrv12 I__7800 (
            .O(N__38021),
            .I(n7_adj_1561));
    Odrv4 I__7799 (
            .O(N__38018),
            .I(n7_adj_1561));
    InMux I__7798 (
            .O(N__38013),
            .I(n19809));
    InMux I__7797 (
            .O(N__38010),
            .I(N__38005));
    InMux I__7796 (
            .O(N__38009),
            .I(N__38002));
    InMux I__7795 (
            .O(N__38008),
            .I(N__37999));
    LocalMux I__7794 (
            .O(N__38005),
            .I(N__37994));
    LocalMux I__7793 (
            .O(N__38002),
            .I(N__37994));
    LocalMux I__7792 (
            .O(N__37999),
            .I(data_index_7));
    Odrv12 I__7791 (
            .O(N__37994),
            .I(data_index_7));
    InMux I__7790 (
            .O(N__37989),
            .I(N__37983));
    InMux I__7789 (
            .O(N__37988),
            .I(N__37983));
    LocalMux I__7788 (
            .O(N__37983),
            .I(N__37980));
    Odrv4 I__7787 (
            .O(N__37980),
            .I(n7_adj_1559));
    InMux I__7786 (
            .O(N__37977),
            .I(n19810));
    InMux I__7785 (
            .O(N__37974),
            .I(bfn_14_16_0_));
    InMux I__7784 (
            .O(N__37971),
            .I(bfn_14_14_0_));
    InMux I__7783 (
            .O(N__37968),
            .I(n19782));
    InMux I__7782 (
            .O(N__37965),
            .I(n19783));
    InMux I__7781 (
            .O(N__37962),
            .I(N__37959));
    LocalMux I__7780 (
            .O(N__37959),
            .I(N__37956));
    Span4Mux_h I__7779 (
            .O(N__37956),
            .I(N__37951));
    InMux I__7778 (
            .O(N__37955),
            .I(N__37948));
    InMux I__7777 (
            .O(N__37954),
            .I(N__37945));
    Span4Mux_v I__7776 (
            .O(N__37951),
            .I(N__37942));
    LocalMux I__7775 (
            .O(N__37948),
            .I(N__37939));
    LocalMux I__7774 (
            .O(N__37945),
            .I(data_cntvec_11));
    Odrv4 I__7773 (
            .O(N__37942),
            .I(data_cntvec_11));
    Odrv12 I__7772 (
            .O(N__37939),
            .I(data_cntvec_11));
    InMux I__7771 (
            .O(N__37932),
            .I(n19784));
    InMux I__7770 (
            .O(N__37929),
            .I(N__37926));
    LocalMux I__7769 (
            .O(N__37926),
            .I(N__37922));
    InMux I__7768 (
            .O(N__37925),
            .I(N__37919));
    Span4Mux_v I__7767 (
            .O(N__37922),
            .I(N__37916));
    LocalMux I__7766 (
            .O(N__37919),
            .I(data_cntvec_12));
    Odrv4 I__7765 (
            .O(N__37916),
            .I(data_cntvec_12));
    InMux I__7764 (
            .O(N__37911),
            .I(n19785));
    InMux I__7763 (
            .O(N__37908),
            .I(N__37905));
    LocalMux I__7762 (
            .O(N__37905),
            .I(N__37901));
    InMux I__7761 (
            .O(N__37904),
            .I(N__37898));
    Span4Mux_h I__7760 (
            .O(N__37901),
            .I(N__37895));
    LocalMux I__7759 (
            .O(N__37898),
            .I(data_cntvec_13));
    Odrv4 I__7758 (
            .O(N__37895),
            .I(data_cntvec_13));
    InMux I__7757 (
            .O(N__37890),
            .I(n19786));
    InMux I__7756 (
            .O(N__37887),
            .I(N__37884));
    LocalMux I__7755 (
            .O(N__37884),
            .I(N__37880));
    InMux I__7754 (
            .O(N__37883),
            .I(N__37877));
    Span12Mux_v I__7753 (
            .O(N__37880),
            .I(N__37874));
    LocalMux I__7752 (
            .O(N__37877),
            .I(data_cntvec_14));
    Odrv12 I__7751 (
            .O(N__37874),
            .I(data_cntvec_14));
    InMux I__7750 (
            .O(N__37869),
            .I(n19787));
    InMux I__7749 (
            .O(N__37866),
            .I(n19788));
    InMux I__7748 (
            .O(N__37863),
            .I(N__37860));
    LocalMux I__7747 (
            .O(N__37860),
            .I(N__37856));
    InMux I__7746 (
            .O(N__37859),
            .I(N__37853));
    Span4Mux_v I__7745 (
            .O(N__37856),
            .I(N__37850));
    LocalMux I__7744 (
            .O(N__37853),
            .I(data_cntvec_15));
    Odrv4 I__7743 (
            .O(N__37850),
            .I(data_cntvec_15));
    CEMux I__7742 (
            .O(N__37845),
            .I(N__37839));
    CEMux I__7741 (
            .O(N__37844),
            .I(N__37836));
    CEMux I__7740 (
            .O(N__37843),
            .I(N__37833));
    CEMux I__7739 (
            .O(N__37842),
            .I(N__37830));
    LocalMux I__7738 (
            .O(N__37839),
            .I(N__37827));
    LocalMux I__7737 (
            .O(N__37836),
            .I(N__37824));
    LocalMux I__7736 (
            .O(N__37833),
            .I(N__37821));
    LocalMux I__7735 (
            .O(N__37830),
            .I(N__37818));
    Span4Mux_h I__7734 (
            .O(N__37827),
            .I(N__37815));
    Span4Mux_h I__7733 (
            .O(N__37824),
            .I(N__37812));
    Span4Mux_h I__7732 (
            .O(N__37821),
            .I(N__37809));
    Span4Mux_h I__7731 (
            .O(N__37818),
            .I(N__37805));
    Span4Mux_v I__7730 (
            .O(N__37815),
            .I(N__37802));
    Span4Mux_h I__7729 (
            .O(N__37812),
            .I(N__37797));
    Span4Mux_h I__7728 (
            .O(N__37809),
            .I(N__37797));
    InMux I__7727 (
            .O(N__37808),
            .I(N__37794));
    Odrv4 I__7726 (
            .O(N__37805),
            .I(n11933));
    Odrv4 I__7725 (
            .O(N__37802),
            .I(n11933));
    Odrv4 I__7724 (
            .O(N__37797),
            .I(n11933));
    LocalMux I__7723 (
            .O(N__37794),
            .I(n11933));
    CascadeMux I__7722 (
            .O(N__37785),
            .I(N__37781));
    CascadeMux I__7721 (
            .O(N__37784),
            .I(N__37776));
    InMux I__7720 (
            .O(N__37781),
            .I(N__37773));
    InMux I__7719 (
            .O(N__37780),
            .I(N__37766));
    InMux I__7718 (
            .O(N__37779),
            .I(N__37766));
    InMux I__7717 (
            .O(N__37776),
            .I(N__37763));
    LocalMux I__7716 (
            .O(N__37773),
            .I(N__37760));
    InMux I__7715 (
            .O(N__37772),
            .I(N__37757));
    InMux I__7714 (
            .O(N__37771),
            .I(N__37754));
    LocalMux I__7713 (
            .O(N__37766),
            .I(N__37751));
    LocalMux I__7712 (
            .O(N__37763),
            .I(N__37748));
    Sp12to4 I__7711 (
            .O(N__37760),
            .I(N__37743));
    LocalMux I__7710 (
            .O(N__37757),
            .I(N__37743));
    LocalMux I__7709 (
            .O(N__37754),
            .I(N__37736));
    Span4Mux_v I__7708 (
            .O(N__37751),
            .I(N__37736));
    Span4Mux_h I__7707 (
            .O(N__37748),
            .I(N__37736));
    Span12Mux_v I__7706 (
            .O(N__37743),
            .I(N__37733));
    Odrv4 I__7705 (
            .O(N__37736),
            .I(iac_raw_buf_N_776));
    Odrv12 I__7704 (
            .O(N__37733),
            .I(iac_raw_buf_N_776));
    InMux I__7703 (
            .O(N__37728),
            .I(n19774));
    InMux I__7702 (
            .O(N__37725),
            .I(N__37722));
    LocalMux I__7701 (
            .O(N__37722),
            .I(N__37718));
    InMux I__7700 (
            .O(N__37721),
            .I(N__37714));
    Span4Mux_v I__7699 (
            .O(N__37718),
            .I(N__37711));
    InMux I__7698 (
            .O(N__37717),
            .I(N__37708));
    LocalMux I__7697 (
            .O(N__37714),
            .I(data_cntvec_2));
    Odrv4 I__7696 (
            .O(N__37711),
            .I(data_cntvec_2));
    LocalMux I__7695 (
            .O(N__37708),
            .I(data_cntvec_2));
    InMux I__7694 (
            .O(N__37701),
            .I(n19775));
    InMux I__7693 (
            .O(N__37698),
            .I(n19776));
    InMux I__7692 (
            .O(N__37695),
            .I(N__37692));
    LocalMux I__7691 (
            .O(N__37692),
            .I(N__37687));
    InMux I__7690 (
            .O(N__37691),
            .I(N__37684));
    InMux I__7689 (
            .O(N__37690),
            .I(N__37681));
    Span4Mux_h I__7688 (
            .O(N__37687),
            .I(N__37678));
    LocalMux I__7687 (
            .O(N__37684),
            .I(data_cntvec_4));
    LocalMux I__7686 (
            .O(N__37681),
            .I(data_cntvec_4));
    Odrv4 I__7685 (
            .O(N__37678),
            .I(data_cntvec_4));
    InMux I__7684 (
            .O(N__37671),
            .I(n19777));
    InMux I__7683 (
            .O(N__37668),
            .I(N__37664));
    InMux I__7682 (
            .O(N__37667),
            .I(N__37661));
    LocalMux I__7681 (
            .O(N__37664),
            .I(N__37657));
    LocalMux I__7680 (
            .O(N__37661),
            .I(N__37654));
    InMux I__7679 (
            .O(N__37660),
            .I(N__37651));
    Span4Mux_h I__7678 (
            .O(N__37657),
            .I(N__37648));
    Span4Mux_h I__7677 (
            .O(N__37654),
            .I(N__37645));
    LocalMux I__7676 (
            .O(N__37651),
            .I(data_cntvec_5));
    Odrv4 I__7675 (
            .O(N__37648),
            .I(data_cntvec_5));
    Odrv4 I__7674 (
            .O(N__37645),
            .I(data_cntvec_5));
    InMux I__7673 (
            .O(N__37638),
            .I(n19778));
    InMux I__7672 (
            .O(N__37635),
            .I(n19779));
    InMux I__7671 (
            .O(N__37632),
            .I(n19780));
    InMux I__7670 (
            .O(N__37629),
            .I(N__37626));
    LocalMux I__7669 (
            .O(N__37626),
            .I(N__37623));
    Span4Mux_h I__7668 (
            .O(N__37623),
            .I(N__37620));
    Span4Mux_h I__7667 (
            .O(N__37620),
            .I(N__37617));
    Odrv4 I__7666 (
            .O(N__37617),
            .I(n22380));
    InMux I__7665 (
            .O(N__37614),
            .I(N__37611));
    LocalMux I__7664 (
            .O(N__37611),
            .I(N__37608));
    Span4Mux_v I__7663 (
            .O(N__37608),
            .I(N__37605));
    Odrv4 I__7662 (
            .O(N__37605),
            .I(n30_adj_1679));
    CascadeMux I__7661 (
            .O(N__37602),
            .I(n8_adj_1689_cascade_));
    CascadeMux I__7660 (
            .O(N__37599),
            .I(n26_adj_1595_cascade_));
    CEMux I__7659 (
            .O(N__37596),
            .I(N__37593));
    LocalMux I__7658 (
            .O(N__37593),
            .I(n18_adj_1615));
    InMux I__7657 (
            .O(N__37590),
            .I(N__37586));
    InMux I__7656 (
            .O(N__37589),
            .I(N__37583));
    LocalMux I__7655 (
            .O(N__37586),
            .I(N__37579));
    LocalMux I__7654 (
            .O(N__37583),
            .I(N__37576));
    CascadeMux I__7653 (
            .O(N__37582),
            .I(N__37573));
    Span4Mux_h I__7652 (
            .O(N__37579),
            .I(N__37567));
    Span4Mux_h I__7651 (
            .O(N__37576),
            .I(N__37564));
    InMux I__7650 (
            .O(N__37573),
            .I(N__37557));
    InMux I__7649 (
            .O(N__37572),
            .I(N__37557));
    InMux I__7648 (
            .O(N__37571),
            .I(N__37557));
    InMux I__7647 (
            .O(N__37570),
            .I(N__37554));
    Odrv4 I__7646 (
            .O(N__37567),
            .I(n16818));
    Odrv4 I__7645 (
            .O(N__37564),
            .I(n16818));
    LocalMux I__7644 (
            .O(N__37557),
            .I(n16818));
    LocalMux I__7643 (
            .O(N__37554),
            .I(n16818));
    InMux I__7642 (
            .O(N__37545),
            .I(N__37542));
    LocalMux I__7641 (
            .O(N__37542),
            .I(n21714));
    CascadeMux I__7640 (
            .O(N__37539),
            .I(n7_cascade_));
    InMux I__7639 (
            .O(N__37536),
            .I(N__37533));
    LocalMux I__7638 (
            .O(N__37533),
            .I(N__37528));
    InMux I__7637 (
            .O(N__37532),
            .I(N__37525));
    InMux I__7636 (
            .O(N__37531),
            .I(N__37519));
    Span4Mux_v I__7635 (
            .O(N__37528),
            .I(N__37514));
    LocalMux I__7634 (
            .O(N__37525),
            .I(N__37514));
    InMux I__7633 (
            .O(N__37524),
            .I(N__37509));
    InMux I__7632 (
            .O(N__37523),
            .I(N__37509));
    InMux I__7631 (
            .O(N__37522),
            .I(N__37506));
    LocalMux I__7630 (
            .O(N__37519),
            .I(N__37503));
    Span4Mux_h I__7629 (
            .O(N__37514),
            .I(N__37498));
    LocalMux I__7628 (
            .O(N__37509),
            .I(N__37498));
    LocalMux I__7627 (
            .O(N__37506),
            .I(N__37493));
    Span4Mux_h I__7626 (
            .O(N__37503),
            .I(N__37488));
    Span4Mux_h I__7625 (
            .O(N__37498),
            .I(N__37488));
    InMux I__7624 (
            .O(N__37497),
            .I(N__37483));
    InMux I__7623 (
            .O(N__37496),
            .I(N__37483));
    Odrv12 I__7622 (
            .O(N__37493),
            .I(n12107));
    Odrv4 I__7621 (
            .O(N__37488),
            .I(n12107));
    LocalMux I__7620 (
            .O(N__37483),
            .I(n12107));
    InMux I__7619 (
            .O(N__37476),
            .I(N__37473));
    LocalMux I__7618 (
            .O(N__37473),
            .I(N__37469));
    InMux I__7617 (
            .O(N__37472),
            .I(N__37466));
    Span4Mux_h I__7616 (
            .O(N__37469),
            .I(N__37461));
    LocalMux I__7615 (
            .O(N__37466),
            .I(N__37461));
    Span4Mux_v I__7614 (
            .O(N__37461),
            .I(N__37458));
    Sp12to4 I__7613 (
            .O(N__37458),
            .I(N__37455));
    Odrv12 I__7612 (
            .O(N__37455),
            .I(n14_adj_1544));
    InMux I__7611 (
            .O(N__37452),
            .I(N__37449));
    LocalMux I__7610 (
            .O(N__37449),
            .I(N__37446));
    Span4Mux_v I__7609 (
            .O(N__37446),
            .I(N__37442));
    InMux I__7608 (
            .O(N__37445),
            .I(N__37439));
    Sp12to4 I__7607 (
            .O(N__37442),
            .I(N__37436));
    LocalMux I__7606 (
            .O(N__37439),
            .I(n14_adj_1575));
    Odrv12 I__7605 (
            .O(N__37436),
            .I(n14_adj_1575));
    InMux I__7604 (
            .O(N__37431),
            .I(N__37428));
    LocalMux I__7603 (
            .O(N__37428),
            .I(N__37425));
    Odrv12 I__7602 (
            .O(N__37425),
            .I(n19_adj_1666));
    CascadeMux I__7601 (
            .O(N__37422),
            .I(N__37419));
    InMux I__7600 (
            .O(N__37419),
            .I(N__37416));
    LocalMux I__7599 (
            .O(N__37416),
            .I(n20_adj_1667));
    InMux I__7598 (
            .O(N__37413),
            .I(N__37410));
    LocalMux I__7597 (
            .O(N__37410),
            .I(n16_adj_1664));
    InMux I__7596 (
            .O(N__37407),
            .I(N__37404));
    LocalMux I__7595 (
            .O(N__37404),
            .I(N__37401));
    Odrv12 I__7594 (
            .O(N__37401),
            .I(n17_adj_1665));
    CascadeMux I__7593 (
            .O(N__37398),
            .I(n22413_cascade_));
    CascadeMux I__7592 (
            .O(N__37395),
            .I(N__37392));
    InMux I__7591 (
            .O(N__37392),
            .I(N__37389));
    LocalMux I__7590 (
            .O(N__37389),
            .I(N__37386));
    Span4Mux_v I__7589 (
            .O(N__37386),
            .I(N__37383));
    Odrv4 I__7588 (
            .O(N__37383),
            .I(n21671));
    InMux I__7587 (
            .O(N__37380),
            .I(N__37377));
    LocalMux I__7586 (
            .O(N__37377),
            .I(N__37374));
    Span4Mux_v I__7585 (
            .O(N__37374),
            .I(N__37371));
    Span4Mux_h I__7584 (
            .O(N__37371),
            .I(N__37368));
    Odrv4 I__7583 (
            .O(N__37368),
            .I(n23_adj_1668));
    CascadeMux I__7582 (
            .O(N__37365),
            .I(n22569_cascade_));
    InMux I__7581 (
            .O(N__37362),
            .I(N__37359));
    LocalMux I__7580 (
            .O(N__37359),
            .I(n21702));
    InMux I__7579 (
            .O(N__37356),
            .I(N__37353));
    LocalMux I__7578 (
            .O(N__37353),
            .I(n22416));
    CascadeMux I__7577 (
            .O(N__37350),
            .I(n22572_cascade_));
    CascadeMux I__7576 (
            .O(N__37347),
            .I(n30_adj_1669_cascade_));
    InMux I__7575 (
            .O(N__37344),
            .I(N__37341));
    LocalMux I__7574 (
            .O(N__37341),
            .I(N__37338));
    Odrv4 I__7573 (
            .O(N__37338),
            .I(n22404));
    InMux I__7572 (
            .O(N__37335),
            .I(N__37332));
    LocalMux I__7571 (
            .O(N__37332),
            .I(N__37329));
    Span4Mux_h I__7570 (
            .O(N__37329),
            .I(N__37326));
    Odrv4 I__7569 (
            .O(N__37326),
            .I(n19_adj_1673));
    CascadeMux I__7568 (
            .O(N__37323),
            .I(N__37320));
    InMux I__7567 (
            .O(N__37320),
            .I(N__37317));
    LocalMux I__7566 (
            .O(N__37317),
            .I(n20_adj_1674));
    InMux I__7565 (
            .O(N__37314),
            .I(N__37304));
    InMux I__7564 (
            .O(N__37313),
            .I(N__37304));
    InMux I__7563 (
            .O(N__37312),
            .I(N__37304));
    InMux I__7562 (
            .O(N__37311),
            .I(N__37301));
    LocalMux I__7561 (
            .O(N__37304),
            .I(\comm_spi.bit_cnt_1 ));
    LocalMux I__7560 (
            .O(N__37301),
            .I(\comm_spi.bit_cnt_1 ));
    InMux I__7559 (
            .O(N__37296),
            .I(N__37289));
    InMux I__7558 (
            .O(N__37295),
            .I(N__37289));
    InMux I__7557 (
            .O(N__37294),
            .I(N__37286));
    LocalMux I__7556 (
            .O(N__37289),
            .I(\comm_spi.bit_cnt_2 ));
    LocalMux I__7555 (
            .O(N__37286),
            .I(\comm_spi.bit_cnt_2 ));
    CascadeMux I__7554 (
            .O(N__37281),
            .I(N__37278));
    InMux I__7553 (
            .O(N__37278),
            .I(N__37265));
    InMux I__7552 (
            .O(N__37277),
            .I(N__37265));
    InMux I__7551 (
            .O(N__37276),
            .I(N__37265));
    InMux I__7550 (
            .O(N__37275),
            .I(N__37265));
    InMux I__7549 (
            .O(N__37274),
            .I(N__37262));
    LocalMux I__7548 (
            .O(N__37265),
            .I(\comm_spi.bit_cnt_0 ));
    LocalMux I__7547 (
            .O(N__37262),
            .I(\comm_spi.bit_cnt_0 ));
    CascadeMux I__7546 (
            .O(N__37257),
            .I(N__37254));
    InMux I__7545 (
            .O(N__37254),
            .I(N__37251));
    LocalMux I__7544 (
            .O(N__37251),
            .I(N__37246));
    InMux I__7543 (
            .O(N__37250),
            .I(N__37243));
    InMux I__7542 (
            .O(N__37249),
            .I(N__37240));
    Span4Mux_h I__7541 (
            .O(N__37246),
            .I(N__37237));
    LocalMux I__7540 (
            .O(N__37243),
            .I(N__37234));
    LocalMux I__7539 (
            .O(N__37240),
            .I(N__37231));
    Span4Mux_h I__7538 (
            .O(N__37237),
            .I(N__37228));
    Span4Mux_h I__7537 (
            .O(N__37234),
            .I(N__37225));
    Span4Mux_v I__7536 (
            .O(N__37231),
            .I(N__37222));
    Span4Mux_v I__7535 (
            .O(N__37228),
            .I(N__37219));
    Span4Mux_h I__7534 (
            .O(N__37225),
            .I(N__37216));
    Span4Mux_h I__7533 (
            .O(N__37222),
            .I(N__37213));
    Odrv4 I__7532 (
            .O(N__37219),
            .I(n14_adj_1579));
    Odrv4 I__7531 (
            .O(N__37216),
            .I(n14_adj_1579));
    Odrv4 I__7530 (
            .O(N__37213),
            .I(n14_adj_1579));
    InMux I__7529 (
            .O(N__37206),
            .I(N__37203));
    LocalMux I__7528 (
            .O(N__37203),
            .I(N__37200));
    Span4Mux_v I__7527 (
            .O(N__37200),
            .I(N__37197));
    Span4Mux_h I__7526 (
            .O(N__37197),
            .I(N__37193));
    InMux I__7525 (
            .O(N__37196),
            .I(N__37190));
    Span4Mux_h I__7524 (
            .O(N__37193),
            .I(N__37187));
    LocalMux I__7523 (
            .O(N__37190),
            .I(n14_adj_1572));
    Odrv4 I__7522 (
            .O(N__37187),
            .I(n14_adj_1572));
    InMux I__7521 (
            .O(N__37182),
            .I(N__37179));
    LocalMux I__7520 (
            .O(N__37179),
            .I(N__37176));
    Odrv4 I__7519 (
            .O(N__37176),
            .I(n4_adj_1637));
    CascadeMux I__7518 (
            .O(N__37173),
            .I(\comm_spi.imosi_cascade_ ));
    SRMux I__7517 (
            .O(N__37170),
            .I(N__37167));
    LocalMux I__7516 (
            .O(N__37167),
            .I(N__37164));
    Span4Mux_h I__7515 (
            .O(N__37164),
            .I(N__37161));
    Odrv4 I__7514 (
            .O(N__37161),
            .I(\comm_spi.DOUT_7__N_786 ));
    SRMux I__7513 (
            .O(N__37158),
            .I(N__37155));
    LocalMux I__7512 (
            .O(N__37155),
            .I(N__37152));
    Odrv12 I__7511 (
            .O(N__37152),
            .I(\comm_spi.imosi_N_792 ));
    CascadeMux I__7510 (
            .O(N__37149),
            .I(n12_adj_1542_cascade_));
    CascadeMux I__7509 (
            .O(N__37146),
            .I(n19986_cascade_));
    InMux I__7508 (
            .O(N__37143),
            .I(N__37140));
    LocalMux I__7507 (
            .O(N__37140),
            .I(n30_adj_1530));
    InMux I__7506 (
            .O(N__37137),
            .I(N__37134));
    LocalMux I__7505 (
            .O(N__37134),
            .I(n33));
    CascadeMux I__7504 (
            .O(N__37131),
            .I(n34_cascade_));
    InMux I__7503 (
            .O(N__37128),
            .I(N__37125));
    LocalMux I__7502 (
            .O(N__37125),
            .I(n31));
    CascadeMux I__7501 (
            .O(N__37122),
            .I(n49_cascade_));
    InMux I__7500 (
            .O(N__37119),
            .I(N__37116));
    LocalMux I__7499 (
            .O(N__37116),
            .I(n32));
    InMux I__7498 (
            .O(N__37113),
            .I(N__37110));
    LocalMux I__7497 (
            .O(N__37110),
            .I(N__37106));
    InMux I__7496 (
            .O(N__37109),
            .I(N__37103));
    Span4Mux_h I__7495 (
            .O(N__37106),
            .I(N__37100));
    LocalMux I__7494 (
            .O(N__37103),
            .I(acadc_skipcnt_13));
    Odrv4 I__7493 (
            .O(N__37100),
            .I(acadc_skipcnt_13));
    InMux I__7492 (
            .O(N__37095),
            .I(n19801));
    InMux I__7491 (
            .O(N__37092),
            .I(N__37089));
    LocalMux I__7490 (
            .O(N__37089),
            .I(N__37086));
    Span4Mux_v I__7489 (
            .O(N__37086),
            .I(N__37082));
    InMux I__7488 (
            .O(N__37085),
            .I(N__37079));
    Sp12to4 I__7487 (
            .O(N__37082),
            .I(N__37076));
    LocalMux I__7486 (
            .O(N__37079),
            .I(acadc_skipcnt_14));
    Odrv12 I__7485 (
            .O(N__37076),
            .I(acadc_skipcnt_14));
    InMux I__7484 (
            .O(N__37071),
            .I(n19802));
    InMux I__7483 (
            .O(N__37068),
            .I(n19803));
    CascadeMux I__7482 (
            .O(N__37065),
            .I(N__37062));
    InMux I__7481 (
            .O(N__37062),
            .I(N__37059));
    LocalMux I__7480 (
            .O(N__37059),
            .I(N__37055));
    InMux I__7479 (
            .O(N__37058),
            .I(N__37052));
    Span12Mux_v I__7478 (
            .O(N__37055),
            .I(N__37049));
    LocalMux I__7477 (
            .O(N__37052),
            .I(acadc_skipcnt_15));
    Odrv12 I__7476 (
            .O(N__37049),
            .I(acadc_skipcnt_15));
    CEMux I__7475 (
            .O(N__37044),
            .I(N__37039));
    CEMux I__7474 (
            .O(N__37043),
            .I(N__37036));
    CEMux I__7473 (
            .O(N__37042),
            .I(N__37032));
    LocalMux I__7472 (
            .O(N__37039),
            .I(N__37027));
    LocalMux I__7471 (
            .O(N__37036),
            .I(N__37027));
    InMux I__7470 (
            .O(N__37035),
            .I(N__37024));
    LocalMux I__7469 (
            .O(N__37032),
            .I(N__37021));
    Span4Mux_v I__7468 (
            .O(N__37027),
            .I(N__37018));
    LocalMux I__7467 (
            .O(N__37024),
            .I(N__37015));
    Span4Mux_v I__7466 (
            .O(N__37021),
            .I(N__37010));
    Span4Mux_h I__7465 (
            .O(N__37018),
            .I(N__37010));
    Span4Mux_h I__7464 (
            .O(N__37015),
            .I(N__37007));
    Span4Mux_h I__7463 (
            .O(N__37010),
            .I(N__37002));
    Span4Mux_v I__7462 (
            .O(N__37007),
            .I(N__37002));
    Odrv4 I__7461 (
            .O(N__37002),
            .I(n11989));
    SRMux I__7460 (
            .O(N__36999),
            .I(N__36995));
    SRMux I__7459 (
            .O(N__36998),
            .I(N__36992));
    LocalMux I__7458 (
            .O(N__36995),
            .I(N__36989));
    LocalMux I__7457 (
            .O(N__36992),
            .I(N__36986));
    Span4Mux_v I__7456 (
            .O(N__36989),
            .I(N__36983));
    Sp12to4 I__7455 (
            .O(N__36986),
            .I(N__36980));
    Span4Mux_v I__7454 (
            .O(N__36983),
            .I(N__36977));
    Odrv12 I__7453 (
            .O(N__36980),
            .I(n14915));
    Odrv4 I__7452 (
            .O(N__36977),
            .I(n14915));
    InMux I__7451 (
            .O(N__36972),
            .I(N__36967));
    InMux I__7450 (
            .O(N__36971),
            .I(N__36964));
    InMux I__7449 (
            .O(N__36970),
            .I(N__36961));
    LocalMux I__7448 (
            .O(N__36967),
            .I(\comm_spi.n23083 ));
    LocalMux I__7447 (
            .O(N__36964),
            .I(\comm_spi.n23083 ));
    LocalMux I__7446 (
            .O(N__36961),
            .I(\comm_spi.n23083 ));
    InMux I__7445 (
            .O(N__36954),
            .I(N__36951));
    LocalMux I__7444 (
            .O(N__36951),
            .I(N__36947));
    InMux I__7443 (
            .O(N__36950),
            .I(N__36944));
    Span4Mux_h I__7442 (
            .O(N__36947),
            .I(N__36939));
    LocalMux I__7441 (
            .O(N__36944),
            .I(N__36939));
    Span4Mux_v I__7440 (
            .O(N__36939),
            .I(N__36936));
    Odrv4 I__7439 (
            .O(N__36936),
            .I(\comm_spi.n14846 ));
    InMux I__7438 (
            .O(N__36933),
            .I(N__36930));
    LocalMux I__7437 (
            .O(N__36930),
            .I(N__36926));
    InMux I__7436 (
            .O(N__36929),
            .I(N__36923));
    Span4Mux_h I__7435 (
            .O(N__36926),
            .I(N__36918));
    LocalMux I__7434 (
            .O(N__36923),
            .I(N__36918));
    Span4Mux_v I__7433 (
            .O(N__36918),
            .I(N__36915));
    Odrv4 I__7432 (
            .O(N__36915),
            .I(\comm_spi.n14847 ));
    InMux I__7431 (
            .O(N__36912),
            .I(N__36908));
    InMux I__7430 (
            .O(N__36911),
            .I(N__36905));
    LocalMux I__7429 (
            .O(N__36908),
            .I(N__36899));
    LocalMux I__7428 (
            .O(N__36905),
            .I(N__36899));
    InMux I__7427 (
            .O(N__36904),
            .I(N__36896));
    Odrv4 I__7426 (
            .O(N__36899),
            .I(\comm_spi.n14808 ));
    LocalMux I__7425 (
            .O(N__36896),
            .I(\comm_spi.n14808 ));
    InMux I__7424 (
            .O(N__36891),
            .I(N__36888));
    LocalMux I__7423 (
            .O(N__36888),
            .I(N__36883));
    InMux I__7422 (
            .O(N__36887),
            .I(N__36880));
    InMux I__7421 (
            .O(N__36886),
            .I(N__36877));
    Span4Mux_v I__7420 (
            .O(N__36883),
            .I(N__36874));
    LocalMux I__7419 (
            .O(N__36880),
            .I(\comm_spi.n14809 ));
    LocalMux I__7418 (
            .O(N__36877),
            .I(\comm_spi.n14809 ));
    Odrv4 I__7417 (
            .O(N__36874),
            .I(\comm_spi.n14809 ));
    CascadeMux I__7416 (
            .O(N__36867),
            .I(N__36864));
    InMux I__7415 (
            .O(N__36864),
            .I(N__36860));
    InMux I__7414 (
            .O(N__36863),
            .I(N__36857));
    LocalMux I__7413 (
            .O(N__36860),
            .I(N__36854));
    LocalMux I__7412 (
            .O(N__36857),
            .I(acadc_skipcnt_5));
    Odrv4 I__7411 (
            .O(N__36854),
            .I(acadc_skipcnt_5));
    InMux I__7410 (
            .O(N__36849),
            .I(n19793));
    CascadeMux I__7409 (
            .O(N__36846),
            .I(N__36843));
    InMux I__7408 (
            .O(N__36843),
            .I(N__36839));
    InMux I__7407 (
            .O(N__36842),
            .I(N__36836));
    LocalMux I__7406 (
            .O(N__36839),
            .I(N__36833));
    LocalMux I__7405 (
            .O(N__36836),
            .I(acadc_skipcnt_6));
    Odrv12 I__7404 (
            .O(N__36833),
            .I(acadc_skipcnt_6));
    InMux I__7403 (
            .O(N__36828),
            .I(n19794));
    CascadeMux I__7402 (
            .O(N__36825),
            .I(N__36822));
    InMux I__7401 (
            .O(N__36822),
            .I(N__36819));
    LocalMux I__7400 (
            .O(N__36819),
            .I(N__36815));
    InMux I__7399 (
            .O(N__36818),
            .I(N__36812));
    Span4Mux_v I__7398 (
            .O(N__36815),
            .I(N__36809));
    LocalMux I__7397 (
            .O(N__36812),
            .I(acadc_skipcnt_7));
    Odrv4 I__7396 (
            .O(N__36809),
            .I(acadc_skipcnt_7));
    InMux I__7395 (
            .O(N__36804),
            .I(n19795));
    InMux I__7394 (
            .O(N__36801),
            .I(N__36798));
    LocalMux I__7393 (
            .O(N__36798),
            .I(N__36794));
    InMux I__7392 (
            .O(N__36797),
            .I(N__36791));
    Span4Mux_h I__7391 (
            .O(N__36794),
            .I(N__36788));
    LocalMux I__7390 (
            .O(N__36791),
            .I(acadc_skipcnt_8));
    Odrv4 I__7389 (
            .O(N__36788),
            .I(acadc_skipcnt_8));
    InMux I__7388 (
            .O(N__36783),
            .I(n19796));
    InMux I__7387 (
            .O(N__36780),
            .I(N__36777));
    LocalMux I__7386 (
            .O(N__36777),
            .I(N__36773));
    InMux I__7385 (
            .O(N__36776),
            .I(N__36770));
    Span4Mux_h I__7384 (
            .O(N__36773),
            .I(N__36767));
    LocalMux I__7383 (
            .O(N__36770),
            .I(acadc_skipcnt_9));
    Odrv4 I__7382 (
            .O(N__36767),
            .I(acadc_skipcnt_9));
    InMux I__7381 (
            .O(N__36762),
            .I(bfn_13_20_0_));
    InMux I__7380 (
            .O(N__36759),
            .I(n19798));
    CascadeMux I__7379 (
            .O(N__36756),
            .I(N__36753));
    InMux I__7378 (
            .O(N__36753),
            .I(N__36750));
    LocalMux I__7377 (
            .O(N__36750),
            .I(N__36747));
    Sp12to4 I__7376 (
            .O(N__36747),
            .I(N__36743));
    InMux I__7375 (
            .O(N__36746),
            .I(N__36740));
    Span12Mux_v I__7374 (
            .O(N__36743),
            .I(N__36737));
    LocalMux I__7373 (
            .O(N__36740),
            .I(acadc_skipcnt_11));
    Odrv12 I__7372 (
            .O(N__36737),
            .I(acadc_skipcnt_11));
    InMux I__7371 (
            .O(N__36732),
            .I(n19799));
    InMux I__7370 (
            .O(N__36729),
            .I(n19800));
    InMux I__7369 (
            .O(N__36726),
            .I(N__36723));
    LocalMux I__7368 (
            .O(N__36723),
            .I(N__36720));
    Span4Mux_v I__7367 (
            .O(N__36720),
            .I(N__36716));
    InMux I__7366 (
            .O(N__36719),
            .I(N__36713));
    Span4Mux_h I__7365 (
            .O(N__36716),
            .I(N__36710));
    LocalMux I__7364 (
            .O(N__36713),
            .I(acadc_skipcnt_1));
    Odrv4 I__7363 (
            .O(N__36710),
            .I(acadc_skipcnt_1));
    InMux I__7362 (
            .O(N__36705),
            .I(bfn_13_19_0_));
    InMux I__7361 (
            .O(N__36702),
            .I(N__36699));
    LocalMux I__7360 (
            .O(N__36699),
            .I(N__36695));
    InMux I__7359 (
            .O(N__36698),
            .I(N__36692));
    Span4Mux_h I__7358 (
            .O(N__36695),
            .I(N__36689));
    LocalMux I__7357 (
            .O(N__36692),
            .I(acadc_skipcnt_2));
    Odrv4 I__7356 (
            .O(N__36689),
            .I(acadc_skipcnt_2));
    InMux I__7355 (
            .O(N__36684),
            .I(n19790));
    InMux I__7354 (
            .O(N__36681),
            .I(N__36677));
    InMux I__7353 (
            .O(N__36680),
            .I(N__36674));
    LocalMux I__7352 (
            .O(N__36677),
            .I(N__36671));
    LocalMux I__7351 (
            .O(N__36674),
            .I(N__36666));
    Span4Mux_v I__7350 (
            .O(N__36671),
            .I(N__36666));
    Odrv4 I__7349 (
            .O(N__36666),
            .I(acadc_skipcnt_3));
    InMux I__7348 (
            .O(N__36663),
            .I(n19791));
    CascadeMux I__7347 (
            .O(N__36660),
            .I(N__36657));
    InMux I__7346 (
            .O(N__36657),
            .I(N__36654));
    LocalMux I__7345 (
            .O(N__36654),
            .I(N__36650));
    InMux I__7344 (
            .O(N__36653),
            .I(N__36647));
    Span4Mux_v I__7343 (
            .O(N__36650),
            .I(N__36644));
    LocalMux I__7342 (
            .O(N__36647),
            .I(acadc_skipcnt_4));
    Odrv4 I__7341 (
            .O(N__36644),
            .I(acadc_skipcnt_4));
    InMux I__7340 (
            .O(N__36639),
            .I(n19792));
    CascadeMux I__7339 (
            .O(N__36636),
            .I(n8_adj_1566_cascade_));
    InMux I__7338 (
            .O(N__36633),
            .I(N__36630));
    LocalMux I__7337 (
            .O(N__36630),
            .I(N__36627));
    Span4Mux_h I__7336 (
            .O(N__36627),
            .I(N__36624));
    Odrv4 I__7335 (
            .O(N__36624),
            .I(\SIG_DDS.tmp_buf_6 ));
    InMux I__7334 (
            .O(N__36621),
            .I(N__36618));
    LocalMux I__7333 (
            .O(N__36618),
            .I(N__36615));
    Odrv4 I__7332 (
            .O(N__36615),
            .I(\SIG_DDS.tmp_buf_7 ));
    InMux I__7331 (
            .O(N__36612),
            .I(N__36609));
    LocalMux I__7330 (
            .O(N__36609),
            .I(N__36606));
    Span4Mux_h I__7329 (
            .O(N__36606),
            .I(N__36602));
    InMux I__7328 (
            .O(N__36605),
            .I(N__36599));
    Span4Mux_h I__7327 (
            .O(N__36602),
            .I(N__36596));
    LocalMux I__7326 (
            .O(N__36599),
            .I(\SIG_DDS.bit_cnt_3 ));
    Odrv4 I__7325 (
            .O(N__36596),
            .I(\SIG_DDS.bit_cnt_3 ));
    InMux I__7324 (
            .O(N__36591),
            .I(N__36588));
    LocalMux I__7323 (
            .O(N__36588),
            .I(N__36585));
    Span4Mux_v I__7322 (
            .O(N__36585),
            .I(N__36582));
    Span4Mux_h I__7321 (
            .O(N__36582),
            .I(N__36579));
    Odrv4 I__7320 (
            .O(N__36579),
            .I(\SIG_DDS.n21744 ));
    InMux I__7319 (
            .O(N__36576),
            .I(N__36573));
    LocalMux I__7318 (
            .O(N__36573),
            .I(N__36570));
    Span4Mux_v I__7317 (
            .O(N__36570),
            .I(N__36565));
    InMux I__7316 (
            .O(N__36569),
            .I(N__36562));
    InMux I__7315 (
            .O(N__36568),
            .I(N__36559));
    Span4Mux_h I__7314 (
            .O(N__36565),
            .I(N__36556));
    LocalMux I__7313 (
            .O(N__36562),
            .I(N__36553));
    LocalMux I__7312 (
            .O(N__36559),
            .I(buf_dds1_7));
    Odrv4 I__7311 (
            .O(N__36556),
            .I(buf_dds1_7));
    Odrv12 I__7310 (
            .O(N__36553),
            .I(buf_dds1_7));
    InMux I__7309 (
            .O(N__36546),
            .I(N__36542));
    CascadeMux I__7308 (
            .O(N__36545),
            .I(N__36539));
    LocalMux I__7307 (
            .O(N__36542),
            .I(N__36536));
    InMux I__7306 (
            .O(N__36539),
            .I(N__36533));
    Span4Mux_v I__7305 (
            .O(N__36536),
            .I(N__36530));
    LocalMux I__7304 (
            .O(N__36533),
            .I(acadc_skipcnt_0));
    Odrv4 I__7303 (
            .O(N__36530),
            .I(acadc_skipcnt_0));
    SRMux I__7302 (
            .O(N__36525),
            .I(N__36522));
    LocalMux I__7301 (
            .O(N__36522),
            .I(N__36519));
    Span4Mux_v I__7300 (
            .O(N__36519),
            .I(N__36516));
    Odrv4 I__7299 (
            .O(N__36516),
            .I(n21226));
    InMux I__7298 (
            .O(N__36513),
            .I(N__36507));
    InMux I__7297 (
            .O(N__36512),
            .I(N__36507));
    LocalMux I__7296 (
            .O(N__36507),
            .I(N__36504));
    Odrv4 I__7295 (
            .O(N__36504),
            .I(n20011));
    InMux I__7294 (
            .O(N__36501),
            .I(N__36498));
    LocalMux I__7293 (
            .O(N__36498),
            .I(N__36495));
    Span4Mux_h I__7292 (
            .O(N__36495),
            .I(N__36492));
    Span4Mux_v I__7291 (
            .O(N__36492),
            .I(N__36489));
    Odrv4 I__7290 (
            .O(N__36489),
            .I(n19_adj_1616));
    InMux I__7289 (
            .O(N__36486),
            .I(N__36482));
    InMux I__7288 (
            .O(N__36485),
            .I(N__36478));
    LocalMux I__7287 (
            .O(N__36482),
            .I(N__36475));
    InMux I__7286 (
            .O(N__36481),
            .I(N__36472));
    LocalMux I__7285 (
            .O(N__36478),
            .I(N__36467));
    Span4Mux_v I__7284 (
            .O(N__36475),
            .I(N__36467));
    LocalMux I__7283 (
            .O(N__36472),
            .I(N__36462));
    Span4Mux_h I__7282 (
            .O(N__36467),
            .I(N__36459));
    InMux I__7281 (
            .O(N__36466),
            .I(N__36454));
    InMux I__7280 (
            .O(N__36465),
            .I(N__36454));
    Span4Mux_v I__7279 (
            .O(N__36462),
            .I(N__36451));
    Span4Mux_h I__7278 (
            .O(N__36459),
            .I(N__36448));
    LocalMux I__7277 (
            .O(N__36454),
            .I(n14_adj_1547));
    Odrv4 I__7276 (
            .O(N__36451),
            .I(n14_adj_1547));
    Odrv4 I__7275 (
            .O(N__36448),
            .I(n14_adj_1547));
    CascadeMux I__7274 (
            .O(N__36441),
            .I(n8_adj_1564_cascade_));
    CascadeMux I__7273 (
            .O(N__36438),
            .I(N__36435));
    CascadeBuf I__7272 (
            .O(N__36435),
            .I(N__36432));
    CascadeMux I__7271 (
            .O(N__36432),
            .I(N__36429));
    CascadeBuf I__7270 (
            .O(N__36429),
            .I(N__36426));
    CascadeMux I__7269 (
            .O(N__36426),
            .I(N__36423));
    CascadeBuf I__7268 (
            .O(N__36423),
            .I(N__36420));
    CascadeMux I__7267 (
            .O(N__36420),
            .I(N__36417));
    CascadeBuf I__7266 (
            .O(N__36417),
            .I(N__36414));
    CascadeMux I__7265 (
            .O(N__36414),
            .I(N__36411));
    CascadeBuf I__7264 (
            .O(N__36411),
            .I(N__36408));
    CascadeMux I__7263 (
            .O(N__36408),
            .I(N__36405));
    CascadeBuf I__7262 (
            .O(N__36405),
            .I(N__36402));
    CascadeMux I__7261 (
            .O(N__36402),
            .I(N__36399));
    CascadeBuf I__7260 (
            .O(N__36399),
            .I(N__36396));
    CascadeMux I__7259 (
            .O(N__36396),
            .I(N__36393));
    CascadeBuf I__7258 (
            .O(N__36393),
            .I(N__36389));
    CascadeMux I__7257 (
            .O(N__36392),
            .I(N__36386));
    CascadeMux I__7256 (
            .O(N__36389),
            .I(N__36383));
    CascadeBuf I__7255 (
            .O(N__36386),
            .I(N__36380));
    CascadeBuf I__7254 (
            .O(N__36383),
            .I(N__36377));
    CascadeMux I__7253 (
            .O(N__36380),
            .I(N__36374));
    CascadeMux I__7252 (
            .O(N__36377),
            .I(N__36371));
    InMux I__7251 (
            .O(N__36374),
            .I(N__36368));
    InMux I__7250 (
            .O(N__36371),
            .I(N__36365));
    LocalMux I__7249 (
            .O(N__36368),
            .I(N__36362));
    LocalMux I__7248 (
            .O(N__36365),
            .I(N__36359));
    Span12Mux_h I__7247 (
            .O(N__36362),
            .I(N__36354));
    Span12Mux_h I__7246 (
            .O(N__36359),
            .I(N__36354));
    Odrv12 I__7245 (
            .O(N__36354),
            .I(data_index_9_N_212_4));
    CascadeMux I__7244 (
            .O(N__36351),
            .I(N__36348));
    InMux I__7243 (
            .O(N__36348),
            .I(N__36345));
    LocalMux I__7242 (
            .O(N__36345),
            .I(N__36341));
    CascadeMux I__7241 (
            .O(N__36344),
            .I(N__36338));
    Span4Mux_v I__7240 (
            .O(N__36341),
            .I(N__36335));
    InMux I__7239 (
            .O(N__36338),
            .I(N__36332));
    Span4Mux_h I__7238 (
            .O(N__36335),
            .I(N__36328));
    LocalMux I__7237 (
            .O(N__36332),
            .I(N__36325));
    InMux I__7236 (
            .O(N__36331),
            .I(N__36322));
    Odrv4 I__7235 (
            .O(N__36328),
            .I(cmd_rdadctmp_9));
    Odrv4 I__7234 (
            .O(N__36325),
            .I(cmd_rdadctmp_9));
    LocalMux I__7233 (
            .O(N__36322),
            .I(cmd_rdadctmp_9));
    InMux I__7232 (
            .O(N__36315),
            .I(N__36312));
    LocalMux I__7231 (
            .O(N__36312),
            .I(N__36309));
    Span4Mux_v I__7230 (
            .O(N__36309),
            .I(N__36306));
    Sp12to4 I__7229 (
            .O(N__36306),
            .I(N__36303));
    Span12Mux_h I__7228 (
            .O(N__36303),
            .I(N__36298));
    InMux I__7227 (
            .O(N__36302),
            .I(N__36293));
    InMux I__7226 (
            .O(N__36301),
            .I(N__36293));
    Odrv12 I__7225 (
            .O(N__36298),
            .I(buf_adcdata_iac_1));
    LocalMux I__7224 (
            .O(N__36293),
            .I(buf_adcdata_iac_1));
    InMux I__7223 (
            .O(N__36288),
            .I(N__36284));
    InMux I__7222 (
            .O(N__36287),
            .I(N__36281));
    LocalMux I__7221 (
            .O(N__36284),
            .I(N__36278));
    LocalMux I__7220 (
            .O(N__36281),
            .I(N__36274));
    Span4Mux_h I__7219 (
            .O(N__36278),
            .I(N__36271));
    InMux I__7218 (
            .O(N__36277),
            .I(N__36268));
    Span4Mux_v I__7217 (
            .O(N__36274),
            .I(N__36263));
    Span4Mux_v I__7216 (
            .O(N__36271),
            .I(N__36263));
    LocalMux I__7215 (
            .O(N__36268),
            .I(buf_dds1_12));
    Odrv4 I__7214 (
            .O(N__36263),
            .I(buf_dds1_12));
    InMux I__7213 (
            .O(N__36258),
            .I(N__36253));
    InMux I__7212 (
            .O(N__36257),
            .I(N__36250));
    InMux I__7211 (
            .O(N__36256),
            .I(N__36247));
    LocalMux I__7210 (
            .O(N__36253),
            .I(N__36244));
    LocalMux I__7209 (
            .O(N__36250),
            .I(buf_dds0_12));
    LocalMux I__7208 (
            .O(N__36247),
            .I(buf_dds0_12));
    Odrv4 I__7207 (
            .O(N__36244),
            .I(buf_dds0_12));
    CascadeMux I__7206 (
            .O(N__36237),
            .I(N__36234));
    InMux I__7205 (
            .O(N__36234),
            .I(N__36231));
    LocalMux I__7204 (
            .O(N__36231),
            .I(N__36228));
    Odrv4 I__7203 (
            .O(N__36228),
            .I(n8_adj_1566));
    IoInMux I__7202 (
            .O(N__36225),
            .I(N__36222));
    LocalMux I__7201 (
            .O(N__36222),
            .I(N__36219));
    Sp12to4 I__7200 (
            .O(N__36219),
            .I(N__36216));
    Span12Mux_v I__7199 (
            .O(N__36216),
            .I(N__36211));
    InMux I__7198 (
            .O(N__36215),
            .I(N__36208));
    InMux I__7197 (
            .O(N__36214),
            .I(N__36205));
    Odrv12 I__7196 (
            .O(N__36211),
            .I(SELIRNG1));
    LocalMux I__7195 (
            .O(N__36208),
            .I(SELIRNG1));
    LocalMux I__7194 (
            .O(N__36205),
            .I(SELIRNG1));
    InMux I__7193 (
            .O(N__36198),
            .I(N__36193));
    InMux I__7192 (
            .O(N__36197),
            .I(N__36190));
    CascadeMux I__7191 (
            .O(N__36196),
            .I(N__36187));
    LocalMux I__7190 (
            .O(N__36193),
            .I(N__36182));
    LocalMux I__7189 (
            .O(N__36190),
            .I(N__36182));
    InMux I__7188 (
            .O(N__36187),
            .I(N__36179));
    Span4Mux_h I__7187 (
            .O(N__36182),
            .I(N__36176));
    LocalMux I__7186 (
            .O(N__36179),
            .I(n14_adj_1546));
    Odrv4 I__7185 (
            .O(N__36176),
            .I(n14_adj_1546));
    InMux I__7184 (
            .O(N__36171),
            .I(N__36167));
    InMux I__7183 (
            .O(N__36170),
            .I(N__36162));
    LocalMux I__7182 (
            .O(N__36167),
            .I(N__36159));
    CascadeMux I__7181 (
            .O(N__36166),
            .I(N__36156));
    InMux I__7180 (
            .O(N__36165),
            .I(N__36153));
    LocalMux I__7179 (
            .O(N__36162),
            .I(N__36150));
    Span4Mux_v I__7178 (
            .O(N__36159),
            .I(N__36147));
    InMux I__7177 (
            .O(N__36156),
            .I(N__36144));
    LocalMux I__7176 (
            .O(N__36153),
            .I(N__36139));
    Span4Mux_v I__7175 (
            .O(N__36150),
            .I(N__36139));
    Span4Mux_h I__7174 (
            .O(N__36147),
            .I(N__36136));
    LocalMux I__7173 (
            .O(N__36144),
            .I(n14_adj_1549));
    Odrv4 I__7172 (
            .O(N__36139),
            .I(n14_adj_1549));
    Odrv4 I__7171 (
            .O(N__36136),
            .I(n14_adj_1549));
    InMux I__7170 (
            .O(N__36129),
            .I(N__36125));
    InMux I__7169 (
            .O(N__36128),
            .I(N__36122));
    LocalMux I__7168 (
            .O(N__36125),
            .I(n8_adj_1562));
    LocalMux I__7167 (
            .O(N__36122),
            .I(n8_adj_1562));
    CascadeMux I__7166 (
            .O(N__36117),
            .I(N__36114));
    CascadeBuf I__7165 (
            .O(N__36114),
            .I(N__36111));
    CascadeMux I__7164 (
            .O(N__36111),
            .I(N__36108));
    CascadeBuf I__7163 (
            .O(N__36108),
            .I(N__36105));
    CascadeMux I__7162 (
            .O(N__36105),
            .I(N__36102));
    CascadeBuf I__7161 (
            .O(N__36102),
            .I(N__36099));
    CascadeMux I__7160 (
            .O(N__36099),
            .I(N__36096));
    CascadeBuf I__7159 (
            .O(N__36096),
            .I(N__36093));
    CascadeMux I__7158 (
            .O(N__36093),
            .I(N__36090));
    CascadeBuf I__7157 (
            .O(N__36090),
            .I(N__36087));
    CascadeMux I__7156 (
            .O(N__36087),
            .I(N__36084));
    CascadeBuf I__7155 (
            .O(N__36084),
            .I(N__36081));
    CascadeMux I__7154 (
            .O(N__36081),
            .I(N__36077));
    CascadeMux I__7153 (
            .O(N__36080),
            .I(N__36074));
    CascadeBuf I__7152 (
            .O(N__36077),
            .I(N__36071));
    CascadeBuf I__7151 (
            .O(N__36074),
            .I(N__36068));
    CascadeMux I__7150 (
            .O(N__36071),
            .I(N__36065));
    CascadeMux I__7149 (
            .O(N__36068),
            .I(N__36062));
    CascadeBuf I__7148 (
            .O(N__36065),
            .I(N__36059));
    InMux I__7147 (
            .O(N__36062),
            .I(N__36056));
    CascadeMux I__7146 (
            .O(N__36059),
            .I(N__36053));
    LocalMux I__7145 (
            .O(N__36056),
            .I(N__36050));
    CascadeBuf I__7144 (
            .O(N__36053),
            .I(N__36047));
    Span4Mux_h I__7143 (
            .O(N__36050),
            .I(N__36044));
    CascadeMux I__7142 (
            .O(N__36047),
            .I(N__36041));
    Span4Mux_v I__7141 (
            .O(N__36044),
            .I(N__36038));
    InMux I__7140 (
            .O(N__36041),
            .I(N__36035));
    Span4Mux_v I__7139 (
            .O(N__36038),
            .I(N__36032));
    LocalMux I__7138 (
            .O(N__36035),
            .I(N__36029));
    Sp12to4 I__7137 (
            .O(N__36032),
            .I(N__36024));
    Span12Mux_s11_v I__7136 (
            .O(N__36029),
            .I(N__36024));
    Odrv12 I__7135 (
            .O(N__36024),
            .I(data_index_9_N_212_6));
    InMux I__7134 (
            .O(N__36021),
            .I(N__36018));
    LocalMux I__7133 (
            .O(N__36018),
            .I(n17_adj_1553));
    IoInMux I__7132 (
            .O(N__36015),
            .I(N__36012));
    LocalMux I__7131 (
            .O(N__36012),
            .I(N__36009));
    Span4Mux_s0_h I__7130 (
            .O(N__36009),
            .I(N__36006));
    Span4Mux_v I__7129 (
            .O(N__36006),
            .I(N__36003));
    Span4Mux_v I__7128 (
            .O(N__36003),
            .I(N__36000));
    Span4Mux_h I__7127 (
            .O(N__36000),
            .I(N__35997));
    Span4Mux_h I__7126 (
            .O(N__35997),
            .I(N__35993));
    InMux I__7125 (
            .O(N__35996),
            .I(N__35990));
    Span4Mux_h I__7124 (
            .O(N__35993),
            .I(N__35984));
    LocalMux I__7123 (
            .O(N__35990),
            .I(N__35984));
    CascadeMux I__7122 (
            .O(N__35989),
            .I(N__35981));
    Span4Mux_h I__7121 (
            .O(N__35984),
            .I(N__35978));
    InMux I__7120 (
            .O(N__35981),
            .I(N__35975));
    Span4Mux_v I__7119 (
            .O(N__35978),
            .I(N__35972));
    LocalMux I__7118 (
            .O(N__35975),
            .I(AMPV_POW));
    Odrv4 I__7117 (
            .O(N__35972),
            .I(AMPV_POW));
    CascadeMux I__7116 (
            .O(N__35967),
            .I(N__35964));
    CascadeBuf I__7115 (
            .O(N__35964),
            .I(N__35961));
    CascadeMux I__7114 (
            .O(N__35961),
            .I(N__35958));
    CascadeBuf I__7113 (
            .O(N__35958),
            .I(N__35955));
    CascadeMux I__7112 (
            .O(N__35955),
            .I(N__35952));
    CascadeBuf I__7111 (
            .O(N__35952),
            .I(N__35949));
    CascadeMux I__7110 (
            .O(N__35949),
            .I(N__35946));
    CascadeBuf I__7109 (
            .O(N__35946),
            .I(N__35943));
    CascadeMux I__7108 (
            .O(N__35943),
            .I(N__35940));
    CascadeBuf I__7107 (
            .O(N__35940),
            .I(N__35937));
    CascadeMux I__7106 (
            .O(N__35937),
            .I(N__35934));
    CascadeBuf I__7105 (
            .O(N__35934),
            .I(N__35931));
    CascadeMux I__7104 (
            .O(N__35931),
            .I(N__35928));
    CascadeBuf I__7103 (
            .O(N__35928),
            .I(N__35925));
    CascadeMux I__7102 (
            .O(N__35925),
            .I(N__35922));
    CascadeBuf I__7101 (
            .O(N__35922),
            .I(N__35918));
    CascadeMux I__7100 (
            .O(N__35921),
            .I(N__35915));
    CascadeMux I__7099 (
            .O(N__35918),
            .I(N__35912));
    CascadeBuf I__7098 (
            .O(N__35915),
            .I(N__35909));
    CascadeBuf I__7097 (
            .O(N__35912),
            .I(N__35906));
    CascadeMux I__7096 (
            .O(N__35909),
            .I(N__35903));
    CascadeMux I__7095 (
            .O(N__35906),
            .I(N__35900));
    InMux I__7094 (
            .O(N__35903),
            .I(N__35897));
    InMux I__7093 (
            .O(N__35900),
            .I(N__35894));
    LocalMux I__7092 (
            .O(N__35897),
            .I(N__35891));
    LocalMux I__7091 (
            .O(N__35894),
            .I(N__35888));
    Span12Mux_h I__7090 (
            .O(N__35891),
            .I(N__35883));
    Span12Mux_h I__7089 (
            .O(N__35888),
            .I(N__35883));
    Odrv12 I__7088 (
            .O(N__35883),
            .I(data_index_9_N_212_3));
    InMux I__7087 (
            .O(N__35880),
            .I(N__35877));
    LocalMux I__7086 (
            .O(N__35877),
            .I(N__35867));
    CascadeMux I__7085 (
            .O(N__35876),
            .I(N__35862));
    InMux I__7084 (
            .O(N__35875),
            .I(N__35852));
    InMux I__7083 (
            .O(N__35874),
            .I(N__35852));
    InMux I__7082 (
            .O(N__35873),
            .I(N__35852));
    InMux I__7081 (
            .O(N__35872),
            .I(N__35847));
    InMux I__7080 (
            .O(N__35871),
            .I(N__35847));
    InMux I__7079 (
            .O(N__35870),
            .I(N__35844));
    Span12Mux_h I__7078 (
            .O(N__35867),
            .I(N__35841));
    InMux I__7077 (
            .O(N__35866),
            .I(N__35834));
    InMux I__7076 (
            .O(N__35865),
            .I(N__35834));
    InMux I__7075 (
            .O(N__35862),
            .I(N__35834));
    InMux I__7074 (
            .O(N__35861),
            .I(N__35829));
    InMux I__7073 (
            .O(N__35860),
            .I(N__35829));
    InMux I__7072 (
            .O(N__35859),
            .I(N__35826));
    LocalMux I__7071 (
            .O(N__35852),
            .I(eis_state_1));
    LocalMux I__7070 (
            .O(N__35847),
            .I(eis_state_1));
    LocalMux I__7069 (
            .O(N__35844),
            .I(eis_state_1));
    Odrv12 I__7068 (
            .O(N__35841),
            .I(eis_state_1));
    LocalMux I__7067 (
            .O(N__35834),
            .I(eis_state_1));
    LocalMux I__7066 (
            .O(N__35829),
            .I(eis_state_1));
    LocalMux I__7065 (
            .O(N__35826),
            .I(eis_state_1));
    InMux I__7064 (
            .O(N__35811),
            .I(N__35808));
    LocalMux I__7063 (
            .O(N__35808),
            .I(N__35804));
    InMux I__7062 (
            .O(N__35807),
            .I(N__35801));
    Span4Mux_v I__7061 (
            .O(N__35804),
            .I(N__35795));
    LocalMux I__7060 (
            .O(N__35801),
            .I(N__35795));
    InMux I__7059 (
            .O(N__35800),
            .I(N__35788));
    Sp12to4 I__7058 (
            .O(N__35795),
            .I(N__35785));
    CascadeMux I__7057 (
            .O(N__35794),
            .I(N__35778));
    InMux I__7056 (
            .O(N__35793),
            .I(N__35768));
    InMux I__7055 (
            .O(N__35792),
            .I(N__35768));
    InMux I__7054 (
            .O(N__35791),
            .I(N__35768));
    LocalMux I__7053 (
            .O(N__35788),
            .I(N__35763));
    Span12Mux_v I__7052 (
            .O(N__35785),
            .I(N__35763));
    InMux I__7051 (
            .O(N__35784),
            .I(N__35752));
    InMux I__7050 (
            .O(N__35783),
            .I(N__35752));
    InMux I__7049 (
            .O(N__35782),
            .I(N__35752));
    InMux I__7048 (
            .O(N__35781),
            .I(N__35752));
    InMux I__7047 (
            .O(N__35778),
            .I(N__35752));
    InMux I__7046 (
            .O(N__35777),
            .I(N__35745));
    InMux I__7045 (
            .O(N__35776),
            .I(N__35745));
    InMux I__7044 (
            .O(N__35775),
            .I(N__35745));
    LocalMux I__7043 (
            .O(N__35768),
            .I(eis_state_2));
    Odrv12 I__7042 (
            .O(N__35763),
            .I(eis_state_2));
    LocalMux I__7041 (
            .O(N__35752),
            .I(eis_state_2));
    LocalMux I__7040 (
            .O(N__35745),
            .I(eis_state_2));
    InMux I__7039 (
            .O(N__35736),
            .I(N__35728));
    SRMux I__7038 (
            .O(N__35735),
            .I(N__35725));
    InMux I__7037 (
            .O(N__35734),
            .I(N__35720));
    InMux I__7036 (
            .O(N__35733),
            .I(N__35720));
    SRMux I__7035 (
            .O(N__35732),
            .I(N__35717));
    InMux I__7034 (
            .O(N__35731),
            .I(N__35714));
    LocalMux I__7033 (
            .O(N__35728),
            .I(N__35711));
    LocalMux I__7032 (
            .O(N__35725),
            .I(N__35703));
    LocalMux I__7031 (
            .O(N__35720),
            .I(N__35698));
    LocalMux I__7030 (
            .O(N__35717),
            .I(N__35698));
    LocalMux I__7029 (
            .O(N__35714),
            .I(N__35695));
    Span4Mux_h I__7028 (
            .O(N__35711),
            .I(N__35692));
    InMux I__7027 (
            .O(N__35710),
            .I(N__35689));
    InMux I__7026 (
            .O(N__35709),
            .I(N__35686));
    InMux I__7025 (
            .O(N__35708),
            .I(N__35681));
    InMux I__7024 (
            .O(N__35707),
            .I(N__35681));
    InMux I__7023 (
            .O(N__35706),
            .I(N__35678));
    Span4Mux_h I__7022 (
            .O(N__35703),
            .I(N__35675));
    Span12Mux_h I__7021 (
            .O(N__35698),
            .I(N__35672));
    Span4Mux_v I__7020 (
            .O(N__35695),
            .I(N__35667));
    Span4Mux_v I__7019 (
            .O(N__35692),
            .I(N__35667));
    LocalMux I__7018 (
            .O(N__35689),
            .I(N__35664));
    LocalMux I__7017 (
            .O(N__35686),
            .I(N__35661));
    LocalMux I__7016 (
            .O(N__35681),
            .I(N__35658));
    LocalMux I__7015 (
            .O(N__35678),
            .I(acadc_rst));
    Odrv4 I__7014 (
            .O(N__35675),
            .I(acadc_rst));
    Odrv12 I__7013 (
            .O(N__35672),
            .I(acadc_rst));
    Odrv4 I__7012 (
            .O(N__35667),
            .I(acadc_rst));
    Odrv12 I__7011 (
            .O(N__35664),
            .I(acadc_rst));
    Odrv4 I__7010 (
            .O(N__35661),
            .I(acadc_rst));
    Odrv4 I__7009 (
            .O(N__35658),
            .I(acadc_rst));
    InMux I__7008 (
            .O(N__35643),
            .I(N__35640));
    LocalMux I__7007 (
            .O(N__35640),
            .I(n66));
    InMux I__7006 (
            .O(N__35637),
            .I(N__35634));
    LocalMux I__7005 (
            .O(N__35634),
            .I(N__35631));
    Span4Mux_h I__7004 (
            .O(N__35631),
            .I(N__35626));
    InMux I__7003 (
            .O(N__35630),
            .I(N__35623));
    InMux I__7002 (
            .O(N__35629),
            .I(N__35620));
    Span4Mux_h I__7001 (
            .O(N__35626),
            .I(N__35617));
    LocalMux I__7000 (
            .O(N__35623),
            .I(N__35614));
    LocalMux I__6999 (
            .O(N__35620),
            .I(buf_dds1_14));
    Odrv4 I__6998 (
            .O(N__35617),
            .I(buf_dds1_14));
    Odrv4 I__6997 (
            .O(N__35614),
            .I(buf_dds1_14));
    InMux I__6996 (
            .O(N__35607),
            .I(N__35604));
    LocalMux I__6995 (
            .O(N__35604),
            .I(N__35599));
    InMux I__6994 (
            .O(N__35603),
            .I(N__35596));
    CascadeMux I__6993 (
            .O(N__35602),
            .I(N__35593));
    Span4Mux_v I__6992 (
            .O(N__35599),
            .I(N__35590));
    LocalMux I__6991 (
            .O(N__35596),
            .I(N__35587));
    InMux I__6990 (
            .O(N__35593),
            .I(N__35584));
    Span4Mux_h I__6989 (
            .O(N__35590),
            .I(N__35581));
    Span4Mux_h I__6988 (
            .O(N__35587),
            .I(N__35578));
    LocalMux I__6987 (
            .O(N__35584),
            .I(buf_dds1_1));
    Odrv4 I__6986 (
            .O(N__35581),
            .I(buf_dds1_1));
    Odrv4 I__6985 (
            .O(N__35578),
            .I(buf_dds1_1));
    InMux I__6984 (
            .O(N__35571),
            .I(N__35562));
    InMux I__6983 (
            .O(N__35570),
            .I(N__35562));
    InMux I__6982 (
            .O(N__35569),
            .I(N__35562));
    LocalMux I__6981 (
            .O(N__35562),
            .I(N__35552));
    InMux I__6980 (
            .O(N__35561),
            .I(N__35547));
    InMux I__6979 (
            .O(N__35560),
            .I(N__35547));
    InMux I__6978 (
            .O(N__35559),
            .I(N__35544));
    InMux I__6977 (
            .O(N__35558),
            .I(N__35539));
    InMux I__6976 (
            .O(N__35557),
            .I(N__35539));
    CascadeMux I__6975 (
            .O(N__35556),
            .I(N__35534));
    InMux I__6974 (
            .O(N__35555),
            .I(N__35530));
    Span4Mux_v I__6973 (
            .O(N__35552),
            .I(N__35525));
    LocalMux I__6972 (
            .O(N__35547),
            .I(N__35525));
    LocalMux I__6971 (
            .O(N__35544),
            .I(N__35520));
    LocalMux I__6970 (
            .O(N__35539),
            .I(N__35520));
    InMux I__6969 (
            .O(N__35538),
            .I(N__35511));
    InMux I__6968 (
            .O(N__35537),
            .I(N__35511));
    InMux I__6967 (
            .O(N__35534),
            .I(N__35511));
    InMux I__6966 (
            .O(N__35533),
            .I(N__35511));
    LocalMux I__6965 (
            .O(N__35530),
            .I(N__35505));
    Span4Mux_v I__6964 (
            .O(N__35525),
            .I(N__35502));
    Span4Mux_v I__6963 (
            .O(N__35520),
            .I(N__35499));
    LocalMux I__6962 (
            .O(N__35511),
            .I(N__35496));
    InMux I__6961 (
            .O(N__35510),
            .I(N__35489));
    InMux I__6960 (
            .O(N__35509),
            .I(N__35489));
    InMux I__6959 (
            .O(N__35508),
            .I(N__35489));
    Odrv12 I__6958 (
            .O(N__35505),
            .I(n12662));
    Odrv4 I__6957 (
            .O(N__35502),
            .I(n12662));
    Odrv4 I__6956 (
            .O(N__35499),
            .I(n12662));
    Odrv4 I__6955 (
            .O(N__35496),
            .I(n12662));
    LocalMux I__6954 (
            .O(N__35489),
            .I(n12662));
    CascadeMux I__6953 (
            .O(N__35478),
            .I(N__35475));
    InMux I__6952 (
            .O(N__35475),
            .I(N__35472));
    LocalMux I__6951 (
            .O(N__35472),
            .I(N__35469));
    Span4Mux_h I__6950 (
            .O(N__35469),
            .I(N__35466));
    Odrv4 I__6949 (
            .O(N__35466),
            .I(n5_adj_1536));
    CascadeMux I__6948 (
            .O(N__35463),
            .I(n7_adj_1650_cascade_));
    InMux I__6947 (
            .O(N__35460),
            .I(N__35457));
    LocalMux I__6946 (
            .O(N__35457),
            .I(N__35453));
    InMux I__6945 (
            .O(N__35456),
            .I(N__35450));
    Span4Mux_v I__6944 (
            .O(N__35453),
            .I(N__35445));
    LocalMux I__6943 (
            .O(N__35450),
            .I(N__35445));
    Odrv4 I__6942 (
            .O(N__35445),
            .I(n12));
    InMux I__6941 (
            .O(N__35442),
            .I(N__35439));
    LocalMux I__6940 (
            .O(N__35439),
            .I(N__35436));
    Span4Mux_h I__6939 (
            .O(N__35436),
            .I(N__35433));
    Odrv4 I__6938 (
            .O(N__35433),
            .I(n16_adj_1645));
    CascadeMux I__6937 (
            .O(N__35430),
            .I(n22641_cascade_));
    InMux I__6936 (
            .O(N__35427),
            .I(N__35424));
    LocalMux I__6935 (
            .O(N__35424),
            .I(N__35420));
    CascadeMux I__6934 (
            .O(N__35423),
            .I(N__35417));
    Span4Mux_v I__6933 (
            .O(N__35420),
            .I(N__35414));
    InMux I__6932 (
            .O(N__35417),
            .I(N__35411));
    Span4Mux_h I__6931 (
            .O(N__35414),
            .I(N__35408));
    LocalMux I__6930 (
            .O(N__35411),
            .I(data_idxvec_2));
    Odrv4 I__6929 (
            .O(N__35408),
            .I(data_idxvec_2));
    CascadeMux I__6928 (
            .O(N__35403),
            .I(n26_adj_1647_cascade_));
    InMux I__6927 (
            .O(N__35400),
            .I(N__35397));
    LocalMux I__6926 (
            .O(N__35397),
            .I(N__35394));
    Span4Mux_h I__6925 (
            .O(N__35394),
            .I(N__35389));
    InMux I__6924 (
            .O(N__35393),
            .I(N__35384));
    InMux I__6923 (
            .O(N__35392),
            .I(N__35384));
    Odrv4 I__6922 (
            .O(N__35389),
            .I(acadc_skipCount_2));
    LocalMux I__6921 (
            .O(N__35384),
            .I(acadc_skipCount_2));
    CascadeMux I__6920 (
            .O(N__35379),
            .I(n22383_cascade_));
    InMux I__6919 (
            .O(N__35376),
            .I(N__35371));
    CascadeMux I__6918 (
            .O(N__35375),
            .I(N__35368));
    CascadeMux I__6917 (
            .O(N__35374),
            .I(N__35365));
    LocalMux I__6916 (
            .O(N__35371),
            .I(N__35362));
    InMux I__6915 (
            .O(N__35368),
            .I(N__35357));
    InMux I__6914 (
            .O(N__35365),
            .I(N__35357));
    Odrv12 I__6913 (
            .O(N__35362),
            .I(req_data_cnt_2));
    LocalMux I__6912 (
            .O(N__35357),
            .I(req_data_cnt_2));
    InMux I__6911 (
            .O(N__35352),
            .I(N__35349));
    LocalMux I__6910 (
            .O(N__35349),
            .I(n22644));
    CascadeMux I__6909 (
            .O(N__35346),
            .I(n22386_cascade_));
    CascadeMux I__6908 (
            .O(N__35343),
            .I(n30_adj_1648_cascade_));
    CascadeMux I__6907 (
            .O(N__35340),
            .I(N__35337));
    InMux I__6906 (
            .O(N__35337),
            .I(N__35332));
    InMux I__6905 (
            .O(N__35336),
            .I(N__35329));
    InMux I__6904 (
            .O(N__35335),
            .I(N__35326));
    LocalMux I__6903 (
            .O(N__35332),
            .I(N__35323));
    LocalMux I__6902 (
            .O(N__35329),
            .I(req_data_cnt_4));
    LocalMux I__6901 (
            .O(N__35326),
            .I(req_data_cnt_4));
    Odrv4 I__6900 (
            .O(N__35323),
            .I(req_data_cnt_4));
    InMux I__6899 (
            .O(N__35316),
            .I(N__35313));
    LocalMux I__6898 (
            .O(N__35313),
            .I(n18_adj_1644));
    InMux I__6897 (
            .O(N__35310),
            .I(N__35306));
    CascadeMux I__6896 (
            .O(N__35309),
            .I(N__35303));
    LocalMux I__6895 (
            .O(N__35306),
            .I(N__35300));
    InMux I__6894 (
            .O(N__35303),
            .I(N__35296));
    Span4Mux_v I__6893 (
            .O(N__35300),
            .I(N__35293));
    InMux I__6892 (
            .O(N__35299),
            .I(N__35290));
    LocalMux I__6891 (
            .O(N__35296),
            .I(N__35287));
    Odrv4 I__6890 (
            .O(N__35293),
            .I(buf_dds0_13));
    LocalMux I__6889 (
            .O(N__35290),
            .I(buf_dds0_13));
    Odrv4 I__6888 (
            .O(N__35287),
            .I(buf_dds0_13));
    CascadeMux I__6887 (
            .O(N__35280),
            .I(N__35276));
    InMux I__6886 (
            .O(N__35279),
            .I(N__35273));
    InMux I__6885 (
            .O(N__35276),
            .I(N__35270));
    LocalMux I__6884 (
            .O(N__35273),
            .I(N__35267));
    LocalMux I__6883 (
            .O(N__35270),
            .I(N__35264));
    Span4Mux_h I__6882 (
            .O(N__35267),
            .I(N__35261));
    Odrv4 I__6881 (
            .O(N__35264),
            .I(n9269));
    Odrv4 I__6880 (
            .O(N__35261),
            .I(n9269));
    CascadeMux I__6879 (
            .O(N__35256),
            .I(n12082_cascade_));
    InMux I__6878 (
            .O(N__35253),
            .I(N__35250));
    LocalMux I__6877 (
            .O(N__35250),
            .I(N__35247));
    Span4Mux_h I__6876 (
            .O(N__35247),
            .I(N__35243));
    InMux I__6875 (
            .O(N__35246),
            .I(N__35240));
    Span4Mux_h I__6874 (
            .O(N__35243),
            .I(N__35237));
    LocalMux I__6873 (
            .O(N__35240),
            .I(N__35234));
    Span4Mux_v I__6872 (
            .O(N__35237),
            .I(N__35231));
    Odrv4 I__6871 (
            .O(N__35234),
            .I(n14_adj_1573));
    Odrv4 I__6870 (
            .O(N__35231),
            .I(n14_adj_1573));
    SRMux I__6869 (
            .O(N__35226),
            .I(N__35223));
    LocalMux I__6868 (
            .O(N__35223),
            .I(N__35220));
    Span4Mux_v I__6867 (
            .O(N__35220),
            .I(N__35217));
    Odrv4 I__6866 (
            .O(N__35217),
            .I(\comm_spi.data_tx_7__N_817 ));
    CascadeMux I__6865 (
            .O(N__35214),
            .I(N__35211));
    InMux I__6864 (
            .O(N__35211),
            .I(N__35207));
    InMux I__6863 (
            .O(N__35210),
            .I(N__35203));
    LocalMux I__6862 (
            .O(N__35207),
            .I(N__35200));
    InMux I__6861 (
            .O(N__35206),
            .I(N__35197));
    LocalMux I__6860 (
            .O(N__35203),
            .I(N__35192));
    Span4Mux_v I__6859 (
            .O(N__35200),
            .I(N__35192));
    LocalMux I__6858 (
            .O(N__35197),
            .I(req_data_cnt_10));
    Odrv4 I__6857 (
            .O(N__35192),
            .I(req_data_cnt_10));
    InMux I__6856 (
            .O(N__35187),
            .I(N__35184));
    LocalMux I__6855 (
            .O(N__35184),
            .I(N__35181));
    Span4Mux_v I__6854 (
            .O(N__35181),
            .I(N__35178));
    Odrv4 I__6853 (
            .O(N__35178),
            .I(n19_adj_1646));
    CascadeMux I__6852 (
            .O(N__35175),
            .I(N__35172));
    InMux I__6851 (
            .O(N__35172),
            .I(N__35169));
    LocalMux I__6850 (
            .O(N__35169),
            .I(N__35166));
    Span4Mux_v I__6849 (
            .O(N__35166),
            .I(N__35163));
    Span4Mux_h I__6848 (
            .O(N__35163),
            .I(N__35160));
    Sp12to4 I__6847 (
            .O(N__35160),
            .I(N__35156));
    InMux I__6846 (
            .O(N__35159),
            .I(N__35153));
    Odrv12 I__6845 (
            .O(N__35156),
            .I(buf_readRTD_2));
    LocalMux I__6844 (
            .O(N__35153),
            .I(buf_readRTD_2));
    InMux I__6843 (
            .O(N__35148),
            .I(N__35145));
    LocalMux I__6842 (
            .O(N__35145),
            .I(N__35141));
    InMux I__6841 (
            .O(N__35144),
            .I(N__35138));
    Span4Mux_h I__6840 (
            .O(N__35141),
            .I(N__35135));
    LocalMux I__6839 (
            .O(N__35138),
            .I(secclk_cnt_9));
    Odrv4 I__6838 (
            .O(N__35135),
            .I(secclk_cnt_9));
    InMux I__6837 (
            .O(N__35130),
            .I(N__35126));
    InMux I__6836 (
            .O(N__35129),
            .I(N__35123));
    LocalMux I__6835 (
            .O(N__35126),
            .I(N__35120));
    LocalMux I__6834 (
            .O(N__35123),
            .I(secclk_cnt_17));
    Odrv4 I__6833 (
            .O(N__35120),
            .I(secclk_cnt_17));
    InMux I__6832 (
            .O(N__35115),
            .I(N__35112));
    LocalMux I__6831 (
            .O(N__35112),
            .I(n10));
    InMux I__6830 (
            .O(N__35109),
            .I(N__35106));
    LocalMux I__6829 (
            .O(N__35106),
            .I(N__35103));
    Span4Mux_v I__6828 (
            .O(N__35103),
            .I(N__35100));
    Span4Mux_h I__6827 (
            .O(N__35100),
            .I(N__35097));
    Odrv4 I__6826 (
            .O(N__35097),
            .I(n19_adj_1683));
    CascadeMux I__6825 (
            .O(N__35094),
            .I(N__35091));
    InMux I__6824 (
            .O(N__35091),
            .I(N__35088));
    LocalMux I__6823 (
            .O(N__35088),
            .I(N__35085));
    Span4Mux_h I__6822 (
            .O(N__35085),
            .I(N__35082));
    Span4Mux_h I__6821 (
            .O(N__35082),
            .I(N__35079));
    Odrv4 I__6820 (
            .O(N__35079),
            .I(n20_adj_1684));
    InMux I__6819 (
            .O(N__35076),
            .I(N__35073));
    LocalMux I__6818 (
            .O(N__35073),
            .I(N__35070));
    Span4Mux_v I__6817 (
            .O(N__35070),
            .I(N__35066));
    CascadeMux I__6816 (
            .O(N__35069),
            .I(N__35063));
    Span4Mux_h I__6815 (
            .O(N__35066),
            .I(N__35060));
    InMux I__6814 (
            .O(N__35063),
            .I(N__35057));
    Odrv4 I__6813 (
            .O(N__35060),
            .I(buf_adcdata_vdc_11));
    LocalMux I__6812 (
            .O(N__35057),
            .I(buf_adcdata_vdc_11));
    InMux I__6811 (
            .O(N__35052),
            .I(N__35049));
    LocalMux I__6810 (
            .O(N__35049),
            .I(N__35046));
    Sp12to4 I__6809 (
            .O(N__35046),
            .I(N__35041));
    InMux I__6808 (
            .O(N__35045),
            .I(N__35038));
    InMux I__6807 (
            .O(N__35044),
            .I(N__35035));
    Span12Mux_v I__6806 (
            .O(N__35041),
            .I(N__35030));
    LocalMux I__6805 (
            .O(N__35038),
            .I(N__35030));
    LocalMux I__6804 (
            .O(N__35035),
            .I(buf_adcdata_vac_11));
    Odrv12 I__6803 (
            .O(N__35030),
            .I(buf_adcdata_vac_11));
    InMux I__6802 (
            .O(N__35025),
            .I(N__35022));
    LocalMux I__6801 (
            .O(N__35022),
            .I(N__35018));
    InMux I__6800 (
            .O(N__35021),
            .I(N__35015));
    Odrv12 I__6799 (
            .O(N__35018),
            .I(buf_readRTD_12));
    LocalMux I__6798 (
            .O(N__35015),
            .I(buf_readRTD_12));
    InMux I__6797 (
            .O(N__35010),
            .I(N__35005));
    InMux I__6796 (
            .O(N__35009),
            .I(N__35000));
    InMux I__6795 (
            .O(N__35008),
            .I(N__35000));
    LocalMux I__6794 (
            .O(N__35005),
            .I(N__34993));
    LocalMux I__6793 (
            .O(N__35000),
            .I(N__34993));
    CascadeMux I__6792 (
            .O(N__34999),
            .I(N__34990));
    InMux I__6791 (
            .O(N__34998),
            .I(N__34987));
    Span4Mux_v I__6790 (
            .O(N__34993),
            .I(N__34984));
    InMux I__6789 (
            .O(N__34990),
            .I(N__34981));
    LocalMux I__6788 (
            .O(N__34987),
            .I(N__34978));
    Odrv4 I__6787 (
            .O(N__34984),
            .I(buf_cfgRTD_4));
    LocalMux I__6786 (
            .O(N__34981),
            .I(buf_cfgRTD_4));
    Odrv4 I__6785 (
            .O(N__34978),
            .I(buf_cfgRTD_4));
    InMux I__6784 (
            .O(N__34971),
            .I(N__34968));
    LocalMux I__6783 (
            .O(N__34968),
            .I(N__34964));
    CascadeMux I__6782 (
            .O(N__34967),
            .I(N__34961));
    Span4Mux_h I__6781 (
            .O(N__34964),
            .I(N__34957));
    InMux I__6780 (
            .O(N__34961),
            .I(N__34954));
    InMux I__6779 (
            .O(N__34960),
            .I(N__34951));
    Span4Mux_h I__6778 (
            .O(N__34957),
            .I(N__34948));
    LocalMux I__6777 (
            .O(N__34954),
            .I(buf_dds1_13));
    LocalMux I__6776 (
            .O(N__34951),
            .I(buf_dds1_13));
    Odrv4 I__6775 (
            .O(N__34948),
            .I(buf_dds1_13));
    InMux I__6774 (
            .O(N__34941),
            .I(N__34934));
    InMux I__6773 (
            .O(N__34940),
            .I(N__34934));
    InMux I__6772 (
            .O(N__34939),
            .I(N__34931));
    LocalMux I__6771 (
            .O(N__34934),
            .I(N__34928));
    LocalMux I__6770 (
            .O(N__34931),
            .I(N__34923));
    Span4Mux_v I__6769 (
            .O(N__34928),
            .I(N__34923));
    Span4Mux_h I__6768 (
            .O(N__34923),
            .I(N__34920));
    Span4Mux_h I__6767 (
            .O(N__34920),
            .I(N__34915));
    InMux I__6766 (
            .O(N__34919),
            .I(N__34912));
    InMux I__6765 (
            .O(N__34918),
            .I(N__34909));
    Odrv4 I__6764 (
            .O(N__34915),
            .I(buf_cfgRTD_5));
    LocalMux I__6763 (
            .O(N__34912),
            .I(buf_cfgRTD_5));
    LocalMux I__6762 (
            .O(N__34909),
            .I(buf_cfgRTD_5));
    InMux I__6761 (
            .O(N__34902),
            .I(N__34899));
    LocalMux I__6760 (
            .O(N__34899),
            .I(N__34896));
    Span4Mux_h I__6759 (
            .O(N__34896),
            .I(N__34893));
    Span4Mux_h I__6758 (
            .O(N__34893),
            .I(N__34889));
    InMux I__6757 (
            .O(N__34892),
            .I(N__34886));
    Odrv4 I__6756 (
            .O(N__34889),
            .I(buf_readRTD_13));
    LocalMux I__6755 (
            .O(N__34886),
            .I(buf_readRTD_13));
    InMux I__6754 (
            .O(N__34881),
            .I(N__34874));
    InMux I__6753 (
            .O(N__34880),
            .I(N__34874));
    InMux I__6752 (
            .O(N__34879),
            .I(N__34871));
    LocalMux I__6751 (
            .O(N__34874),
            .I(req_data_cnt_12));
    LocalMux I__6750 (
            .O(N__34871),
            .I(req_data_cnt_12));
    InMux I__6749 (
            .O(N__34866),
            .I(N__34863));
    LocalMux I__6748 (
            .O(N__34863),
            .I(n22));
    InMux I__6747 (
            .O(N__34860),
            .I(N__34856));
    InMux I__6746 (
            .O(N__34859),
            .I(N__34852));
    LocalMux I__6745 (
            .O(N__34856),
            .I(N__34848));
    InMux I__6744 (
            .O(N__34855),
            .I(N__34845));
    LocalMux I__6743 (
            .O(N__34852),
            .I(N__34842));
    InMux I__6742 (
            .O(N__34851),
            .I(N__34839));
    Span4Mux_v I__6741 (
            .O(N__34848),
            .I(N__34836));
    LocalMux I__6740 (
            .O(N__34845),
            .I(N__34833));
    Span4Mux_v I__6739 (
            .O(N__34842),
            .I(N__34830));
    LocalMux I__6738 (
            .O(N__34839),
            .I(N__34827));
    Sp12to4 I__6737 (
            .O(N__34836),
            .I(N__34822));
    Sp12to4 I__6736 (
            .O(N__34833),
            .I(N__34822));
    Span4Mux_h I__6735 (
            .O(N__34830),
            .I(N__34819));
    Sp12to4 I__6734 (
            .O(N__34827),
            .I(N__34816));
    Span12Mux_h I__6733 (
            .O(N__34822),
            .I(N__34813));
    Odrv4 I__6732 (
            .O(N__34819),
            .I(n14_adj_1548));
    Odrv12 I__6731 (
            .O(N__34816),
            .I(n14_adj_1548));
    Odrv12 I__6730 (
            .O(N__34813),
            .I(n14_adj_1548));
    InMux I__6729 (
            .O(N__34806),
            .I(N__34801));
    InMux I__6728 (
            .O(N__34805),
            .I(N__34798));
    InMux I__6727 (
            .O(N__34804),
            .I(N__34795));
    LocalMux I__6726 (
            .O(N__34801),
            .I(\comm_spi.n23095 ));
    LocalMux I__6725 (
            .O(N__34798),
            .I(\comm_spi.n23095 ));
    LocalMux I__6724 (
            .O(N__34795),
            .I(\comm_spi.n23095 ));
    SRMux I__6723 (
            .O(N__34788),
            .I(N__34785));
    LocalMux I__6722 (
            .O(N__34785),
            .I(N__34782));
    Span4Mux_h I__6721 (
            .O(N__34782),
            .I(N__34779));
    Odrv4 I__6720 (
            .O(N__34779),
            .I(\comm_spi.data_tx_7__N_807 ));
    InMux I__6719 (
            .O(N__34776),
            .I(N__34773));
    LocalMux I__6718 (
            .O(N__34773),
            .I(N__34770));
    Span4Mux_h I__6717 (
            .O(N__34770),
            .I(N__34765));
    InMux I__6716 (
            .O(N__34769),
            .I(N__34760));
    InMux I__6715 (
            .O(N__34768),
            .I(N__34760));
    Odrv4 I__6714 (
            .O(N__34765),
            .I(req_data_cnt_13));
    LocalMux I__6713 (
            .O(N__34760),
            .I(req_data_cnt_13));
    InMux I__6712 (
            .O(N__34755),
            .I(\ADC_VDC.n19924 ));
    InMux I__6711 (
            .O(N__34752),
            .I(N__34747));
    InMux I__6710 (
            .O(N__34751),
            .I(N__34742));
    InMux I__6709 (
            .O(N__34750),
            .I(N__34742));
    LocalMux I__6708 (
            .O(N__34747),
            .I(\ADC_VDC.bit_cnt_7 ));
    LocalMux I__6707 (
            .O(N__34742),
            .I(\ADC_VDC.bit_cnt_7 ));
    SRMux I__6706 (
            .O(N__34737),
            .I(N__34734));
    LocalMux I__6705 (
            .O(N__34734),
            .I(N__34731));
    Odrv4 I__6704 (
            .O(N__34731),
            .I(\ADC_VDC.n15273 ));
    CascadeMux I__6703 (
            .O(N__34728),
            .I(N__34725));
    InMux I__6702 (
            .O(N__34725),
            .I(N__34722));
    LocalMux I__6701 (
            .O(N__34722),
            .I(N__34719));
    Odrv4 I__6700 (
            .O(N__34719),
            .I(n21_adj_1594));
    SRMux I__6699 (
            .O(N__34716),
            .I(N__34711));
    SRMux I__6698 (
            .O(N__34715),
            .I(N__34708));
    SRMux I__6697 (
            .O(N__34714),
            .I(N__34705));
    LocalMux I__6696 (
            .O(N__34711),
            .I(N__34702));
    LocalMux I__6695 (
            .O(N__34708),
            .I(N__34697));
    LocalMux I__6694 (
            .O(N__34705),
            .I(N__34697));
    Span4Mux_h I__6693 (
            .O(N__34702),
            .I(N__34694));
    Sp12to4 I__6692 (
            .O(N__34697),
            .I(N__34690));
    Span4Mux_h I__6691 (
            .O(N__34694),
            .I(N__34687));
    InMux I__6690 (
            .O(N__34693),
            .I(N__34684));
    Odrv12 I__6689 (
            .O(N__34690),
            .I(n14899));
    Odrv4 I__6688 (
            .O(N__34687),
            .I(n14899));
    LocalMux I__6687 (
            .O(N__34684),
            .I(n14899));
    IoInMux I__6686 (
            .O(N__34677),
            .I(N__34674));
    LocalMux I__6685 (
            .O(N__34674),
            .I(N__34671));
    IoSpan4Mux I__6684 (
            .O(N__34671),
            .I(N__34668));
    Span4Mux_s3_v I__6683 (
            .O(N__34668),
            .I(N__34665));
    Sp12to4 I__6682 (
            .O(N__34665),
            .I(N__34661));
    InMux I__6681 (
            .O(N__34664),
            .I(N__34658));
    Span12Mux_h I__6680 (
            .O(N__34661),
            .I(N__34655));
    LocalMux I__6679 (
            .O(N__34658),
            .I(N__34652));
    Odrv12 I__6678 (
            .O(N__34655),
            .I(TEST_LED));
    Odrv4 I__6677 (
            .O(N__34652),
            .I(TEST_LED));
    InMux I__6676 (
            .O(N__34647),
            .I(N__34644));
    LocalMux I__6675 (
            .O(N__34644),
            .I(N__34640));
    InMux I__6674 (
            .O(N__34643),
            .I(N__34637));
    Span4Mux_h I__6673 (
            .O(N__34640),
            .I(N__34634));
    LocalMux I__6672 (
            .O(N__34637),
            .I(secclk_cnt_15));
    Odrv4 I__6671 (
            .O(N__34634),
            .I(secclk_cnt_15));
    InMux I__6670 (
            .O(N__34629),
            .I(N__34626));
    LocalMux I__6669 (
            .O(N__34626),
            .I(N__34622));
    InMux I__6668 (
            .O(N__34625),
            .I(N__34619));
    Span4Mux_v I__6667 (
            .O(N__34622),
            .I(N__34616));
    LocalMux I__6666 (
            .O(N__34619),
            .I(secclk_cnt_8));
    Odrv4 I__6665 (
            .O(N__34616),
            .I(secclk_cnt_8));
    CascadeMux I__6664 (
            .O(N__34611),
            .I(N__34607));
    InMux I__6663 (
            .O(N__34610),
            .I(N__34604));
    InMux I__6662 (
            .O(N__34607),
            .I(N__34601));
    LocalMux I__6661 (
            .O(N__34604),
            .I(N__34596));
    LocalMux I__6660 (
            .O(N__34601),
            .I(N__34596));
    Odrv4 I__6659 (
            .O(N__34596),
            .I(secclk_cnt_1));
    InMux I__6658 (
            .O(N__34593),
            .I(N__34589));
    InMux I__6657 (
            .O(N__34592),
            .I(N__34586));
    LocalMux I__6656 (
            .O(N__34589),
            .I(N__34583));
    LocalMux I__6655 (
            .O(N__34586),
            .I(secclk_cnt_5));
    Odrv4 I__6654 (
            .O(N__34583),
            .I(secclk_cnt_5));
    InMux I__6653 (
            .O(N__34578),
            .I(N__34575));
    LocalMux I__6652 (
            .O(N__34575),
            .I(n25));
    InMux I__6651 (
            .O(N__34572),
            .I(N__34568));
    InMux I__6650 (
            .O(N__34571),
            .I(N__34565));
    LocalMux I__6649 (
            .O(N__34568),
            .I(N__34562));
    LocalMux I__6648 (
            .O(N__34565),
            .I(N__34557));
    Span4Mux_v I__6647 (
            .O(N__34562),
            .I(N__34557));
    Odrv4 I__6646 (
            .O(N__34557),
            .I(secclk_cnt_18));
    InMux I__6645 (
            .O(N__34554),
            .I(N__34550));
    InMux I__6644 (
            .O(N__34553),
            .I(N__34547));
    LocalMux I__6643 (
            .O(N__34550),
            .I(N__34542));
    LocalMux I__6642 (
            .O(N__34547),
            .I(N__34542));
    Odrv4 I__6641 (
            .O(N__34542),
            .I(secclk_cnt_0));
    CascadeMux I__6640 (
            .O(N__34539),
            .I(N__34536));
    InMux I__6639 (
            .O(N__34536),
            .I(N__34533));
    LocalMux I__6638 (
            .O(N__34533),
            .I(N__34529));
    InMux I__6637 (
            .O(N__34532),
            .I(N__34526));
    Span4Mux_h I__6636 (
            .O(N__34529),
            .I(N__34523));
    LocalMux I__6635 (
            .O(N__34526),
            .I(secclk_cnt_11));
    Odrv4 I__6634 (
            .O(N__34523),
            .I(secclk_cnt_11));
    InMux I__6633 (
            .O(N__34518),
            .I(N__34514));
    InMux I__6632 (
            .O(N__34517),
            .I(N__34511));
    LocalMux I__6631 (
            .O(N__34514),
            .I(N__34508));
    LocalMux I__6630 (
            .O(N__34511),
            .I(secclk_cnt_4));
    Odrv12 I__6629 (
            .O(N__34508),
            .I(secclk_cnt_4));
    CascadeMux I__6628 (
            .O(N__34503),
            .I(N__34500));
    InMux I__6627 (
            .O(N__34500),
            .I(N__34497));
    LocalMux I__6626 (
            .O(N__34497),
            .I(n28_adj_1554));
    InMux I__6625 (
            .O(N__34494),
            .I(N__34491));
    LocalMux I__6624 (
            .O(N__34491),
            .I(N__34488));
    Span4Mux_h I__6623 (
            .O(N__34488),
            .I(N__34484));
    CascadeMux I__6622 (
            .O(N__34487),
            .I(N__34481));
    Span4Mux_v I__6621 (
            .O(N__34484),
            .I(N__34477));
    InMux I__6620 (
            .O(N__34481),
            .I(N__34474));
    InMux I__6619 (
            .O(N__34480),
            .I(N__34471));
    Span4Mux_h I__6618 (
            .O(N__34477),
            .I(N__34466));
    LocalMux I__6617 (
            .O(N__34474),
            .I(N__34466));
    LocalMux I__6616 (
            .O(N__34471),
            .I(req_data_cnt_15));
    Odrv4 I__6615 (
            .O(N__34466),
            .I(req_data_cnt_15));
    InMux I__6614 (
            .O(N__34461),
            .I(N__34458));
    LocalMux I__6613 (
            .O(N__34458),
            .I(n24));
    InMux I__6612 (
            .O(N__34455),
            .I(N__34452));
    LocalMux I__6611 (
            .O(N__34452),
            .I(\comm_spi.n14822 ));
    CascadeMux I__6610 (
            .O(N__34449),
            .I(\comm_spi.n23089_cascade_ ));
    InMux I__6609 (
            .O(N__34446),
            .I(N__34443));
    LocalMux I__6608 (
            .O(N__34443),
            .I(\comm_spi.n14823 ));
    CascadeMux I__6607 (
            .O(N__34440),
            .I(N__34437));
    InMux I__6606 (
            .O(N__34437),
            .I(N__34433));
    CascadeMux I__6605 (
            .O(N__34436),
            .I(N__34430));
    LocalMux I__6604 (
            .O(N__34433),
            .I(N__34426));
    InMux I__6603 (
            .O(N__34430),
            .I(N__34423));
    InMux I__6602 (
            .O(N__34429),
            .I(N__34419));
    Span4Mux_v I__6601 (
            .O(N__34426),
            .I(N__34414));
    LocalMux I__6600 (
            .O(N__34423),
            .I(N__34414));
    InMux I__6599 (
            .O(N__34422),
            .I(N__34411));
    LocalMux I__6598 (
            .O(N__34419),
            .I(\ADC_VDC.bit_cnt_0 ));
    Odrv4 I__6597 (
            .O(N__34414),
            .I(\ADC_VDC.bit_cnt_0 ));
    LocalMux I__6596 (
            .O(N__34411),
            .I(\ADC_VDC.bit_cnt_0 ));
    InMux I__6595 (
            .O(N__34404),
            .I(bfn_13_6_0_));
    InMux I__6594 (
            .O(N__34401),
            .I(N__34398));
    LocalMux I__6593 (
            .O(N__34398),
            .I(N__34394));
    InMux I__6592 (
            .O(N__34397),
            .I(N__34390));
    Span4Mux_h I__6591 (
            .O(N__34394),
            .I(N__34387));
    InMux I__6590 (
            .O(N__34393),
            .I(N__34384));
    LocalMux I__6589 (
            .O(N__34390),
            .I(\ADC_VDC.bit_cnt_1 ));
    Odrv4 I__6588 (
            .O(N__34387),
            .I(\ADC_VDC.bit_cnt_1 ));
    LocalMux I__6587 (
            .O(N__34384),
            .I(\ADC_VDC.bit_cnt_1 ));
    InMux I__6586 (
            .O(N__34377),
            .I(\ADC_VDC.n19918 ));
    InMux I__6585 (
            .O(N__34374),
            .I(N__34370));
    InMux I__6584 (
            .O(N__34373),
            .I(N__34366));
    LocalMux I__6583 (
            .O(N__34370),
            .I(N__34363));
    InMux I__6582 (
            .O(N__34369),
            .I(N__34360));
    LocalMux I__6581 (
            .O(N__34366),
            .I(N__34354));
    Span4Mux_v I__6580 (
            .O(N__34363),
            .I(N__34354));
    LocalMux I__6579 (
            .O(N__34360),
            .I(N__34351));
    InMux I__6578 (
            .O(N__34359),
            .I(N__34348));
    Odrv4 I__6577 (
            .O(N__34354),
            .I(\ADC_VDC.bit_cnt_2 ));
    Odrv4 I__6576 (
            .O(N__34351),
            .I(\ADC_VDC.bit_cnt_2 ));
    LocalMux I__6575 (
            .O(N__34348),
            .I(\ADC_VDC.bit_cnt_2 ));
    InMux I__6574 (
            .O(N__34341),
            .I(\ADC_VDC.n19919 ));
    InMux I__6573 (
            .O(N__34338),
            .I(N__34334));
    InMux I__6572 (
            .O(N__34337),
            .I(N__34330));
    LocalMux I__6571 (
            .O(N__34334),
            .I(N__34327));
    InMux I__6570 (
            .O(N__34333),
            .I(N__34323));
    LocalMux I__6569 (
            .O(N__34330),
            .I(N__34318));
    Span4Mux_v I__6568 (
            .O(N__34327),
            .I(N__34318));
    InMux I__6567 (
            .O(N__34326),
            .I(N__34315));
    LocalMux I__6566 (
            .O(N__34323),
            .I(\ADC_VDC.bit_cnt_3 ));
    Odrv4 I__6565 (
            .O(N__34318),
            .I(\ADC_VDC.bit_cnt_3 ));
    LocalMux I__6564 (
            .O(N__34315),
            .I(\ADC_VDC.bit_cnt_3 ));
    InMux I__6563 (
            .O(N__34308),
            .I(\ADC_VDC.n19920 ));
    InMux I__6562 (
            .O(N__34305),
            .I(N__34302));
    LocalMux I__6561 (
            .O(N__34302),
            .I(N__34298));
    InMux I__6560 (
            .O(N__34301),
            .I(N__34293));
    Span4Mux_h I__6559 (
            .O(N__34298),
            .I(N__34290));
    InMux I__6558 (
            .O(N__34297),
            .I(N__34285));
    InMux I__6557 (
            .O(N__34296),
            .I(N__34285));
    LocalMux I__6556 (
            .O(N__34293),
            .I(\ADC_VDC.bit_cnt_4 ));
    Odrv4 I__6555 (
            .O(N__34290),
            .I(\ADC_VDC.bit_cnt_4 ));
    LocalMux I__6554 (
            .O(N__34285),
            .I(\ADC_VDC.bit_cnt_4 ));
    InMux I__6553 (
            .O(N__34278),
            .I(\ADC_VDC.n19921 ));
    CascadeMux I__6552 (
            .O(N__34275),
            .I(N__34270));
    InMux I__6551 (
            .O(N__34274),
            .I(N__34267));
    InMux I__6550 (
            .O(N__34273),
            .I(N__34262));
    InMux I__6549 (
            .O(N__34270),
            .I(N__34262));
    LocalMux I__6548 (
            .O(N__34267),
            .I(\ADC_VDC.bit_cnt_5 ));
    LocalMux I__6547 (
            .O(N__34262),
            .I(\ADC_VDC.bit_cnt_5 ));
    InMux I__6546 (
            .O(N__34257),
            .I(\ADC_VDC.n19922 ));
    InMux I__6545 (
            .O(N__34254),
            .I(N__34249));
    InMux I__6544 (
            .O(N__34253),
            .I(N__34244));
    InMux I__6543 (
            .O(N__34252),
            .I(N__34244));
    LocalMux I__6542 (
            .O(N__34249),
            .I(\ADC_VDC.bit_cnt_6 ));
    LocalMux I__6541 (
            .O(N__34244),
            .I(\ADC_VDC.bit_cnt_6 ));
    InMux I__6540 (
            .O(N__34239),
            .I(\ADC_VDC.n19923 ));
    CascadeMux I__6539 (
            .O(N__34236),
            .I(N__34233));
    CascadeBuf I__6538 (
            .O(N__34233),
            .I(N__34230));
    CascadeMux I__6537 (
            .O(N__34230),
            .I(N__34227));
    CascadeBuf I__6536 (
            .O(N__34227),
            .I(N__34224));
    CascadeMux I__6535 (
            .O(N__34224),
            .I(N__34221));
    CascadeBuf I__6534 (
            .O(N__34221),
            .I(N__34218));
    CascadeMux I__6533 (
            .O(N__34218),
            .I(N__34215));
    CascadeBuf I__6532 (
            .O(N__34215),
            .I(N__34212));
    CascadeMux I__6531 (
            .O(N__34212),
            .I(N__34209));
    CascadeBuf I__6530 (
            .O(N__34209),
            .I(N__34206));
    CascadeMux I__6529 (
            .O(N__34206),
            .I(N__34203));
    CascadeBuf I__6528 (
            .O(N__34203),
            .I(N__34200));
    CascadeMux I__6527 (
            .O(N__34200),
            .I(N__34197));
    CascadeBuf I__6526 (
            .O(N__34197),
            .I(N__34194));
    CascadeMux I__6525 (
            .O(N__34194),
            .I(N__34190));
    CascadeMux I__6524 (
            .O(N__34193),
            .I(N__34187));
    CascadeBuf I__6523 (
            .O(N__34190),
            .I(N__34184));
    CascadeBuf I__6522 (
            .O(N__34187),
            .I(N__34181));
    CascadeMux I__6521 (
            .O(N__34184),
            .I(N__34178));
    CascadeMux I__6520 (
            .O(N__34181),
            .I(N__34175));
    CascadeBuf I__6519 (
            .O(N__34178),
            .I(N__34172));
    InMux I__6518 (
            .O(N__34175),
            .I(N__34169));
    CascadeMux I__6517 (
            .O(N__34172),
            .I(N__34166));
    LocalMux I__6516 (
            .O(N__34169),
            .I(N__34163));
    InMux I__6515 (
            .O(N__34166),
            .I(N__34160));
    Span4Mux_h I__6514 (
            .O(N__34163),
            .I(N__34157));
    LocalMux I__6513 (
            .O(N__34160),
            .I(N__34154));
    Sp12to4 I__6512 (
            .O(N__34157),
            .I(N__34150));
    Span4Mux_v I__6511 (
            .O(N__34154),
            .I(N__34147));
    InMux I__6510 (
            .O(N__34153),
            .I(N__34144));
    Span12Mux_v I__6509 (
            .O(N__34150),
            .I(N__34141));
    Sp12to4 I__6508 (
            .O(N__34147),
            .I(N__34138));
    LocalMux I__6507 (
            .O(N__34144),
            .I(data_count_6));
    Odrv12 I__6506 (
            .O(N__34141),
            .I(data_count_6));
    Odrv12 I__6505 (
            .O(N__34138),
            .I(data_count_6));
    InMux I__6504 (
            .O(N__34131),
            .I(n19770));
    CascadeMux I__6503 (
            .O(N__34128),
            .I(N__34125));
    CascadeBuf I__6502 (
            .O(N__34125),
            .I(N__34122));
    CascadeMux I__6501 (
            .O(N__34122),
            .I(N__34119));
    CascadeBuf I__6500 (
            .O(N__34119),
            .I(N__34116));
    CascadeMux I__6499 (
            .O(N__34116),
            .I(N__34113));
    CascadeBuf I__6498 (
            .O(N__34113),
            .I(N__34110));
    CascadeMux I__6497 (
            .O(N__34110),
            .I(N__34107));
    CascadeBuf I__6496 (
            .O(N__34107),
            .I(N__34104));
    CascadeMux I__6495 (
            .O(N__34104),
            .I(N__34101));
    CascadeBuf I__6494 (
            .O(N__34101),
            .I(N__34098));
    CascadeMux I__6493 (
            .O(N__34098),
            .I(N__34095));
    CascadeBuf I__6492 (
            .O(N__34095),
            .I(N__34092));
    CascadeMux I__6491 (
            .O(N__34092),
            .I(N__34088));
    CascadeMux I__6490 (
            .O(N__34091),
            .I(N__34085));
    CascadeBuf I__6489 (
            .O(N__34088),
            .I(N__34082));
    CascadeBuf I__6488 (
            .O(N__34085),
            .I(N__34079));
    CascadeMux I__6487 (
            .O(N__34082),
            .I(N__34076));
    CascadeMux I__6486 (
            .O(N__34079),
            .I(N__34073));
    CascadeBuf I__6485 (
            .O(N__34076),
            .I(N__34070));
    InMux I__6484 (
            .O(N__34073),
            .I(N__34067));
    CascadeMux I__6483 (
            .O(N__34070),
            .I(N__34064));
    LocalMux I__6482 (
            .O(N__34067),
            .I(N__34061));
    CascadeBuf I__6481 (
            .O(N__34064),
            .I(N__34058));
    Span4Mux_h I__6480 (
            .O(N__34061),
            .I(N__34055));
    CascadeMux I__6479 (
            .O(N__34058),
            .I(N__34052));
    Span4Mux_h I__6478 (
            .O(N__34055),
            .I(N__34049));
    InMux I__6477 (
            .O(N__34052),
            .I(N__34046));
    Sp12to4 I__6476 (
            .O(N__34049),
            .I(N__34042));
    LocalMux I__6475 (
            .O(N__34046),
            .I(N__34039));
    InMux I__6474 (
            .O(N__34045),
            .I(N__34036));
    Span12Mux_v I__6473 (
            .O(N__34042),
            .I(N__34033));
    Span12Mux_s8_v I__6472 (
            .O(N__34039),
            .I(N__34030));
    LocalMux I__6471 (
            .O(N__34036),
            .I(data_count_7));
    Odrv12 I__6470 (
            .O(N__34033),
            .I(data_count_7));
    Odrv12 I__6469 (
            .O(N__34030),
            .I(data_count_7));
    InMux I__6468 (
            .O(N__34023),
            .I(n19771));
    CascadeMux I__6467 (
            .O(N__34020),
            .I(N__34017));
    CascadeBuf I__6466 (
            .O(N__34017),
            .I(N__34014));
    CascadeMux I__6465 (
            .O(N__34014),
            .I(N__34011));
    CascadeBuf I__6464 (
            .O(N__34011),
            .I(N__34008));
    CascadeMux I__6463 (
            .O(N__34008),
            .I(N__34005));
    CascadeBuf I__6462 (
            .O(N__34005),
            .I(N__34002));
    CascadeMux I__6461 (
            .O(N__34002),
            .I(N__33999));
    CascadeBuf I__6460 (
            .O(N__33999),
            .I(N__33996));
    CascadeMux I__6459 (
            .O(N__33996),
            .I(N__33993));
    CascadeBuf I__6458 (
            .O(N__33993),
            .I(N__33990));
    CascadeMux I__6457 (
            .O(N__33990),
            .I(N__33987));
    CascadeBuf I__6456 (
            .O(N__33987),
            .I(N__33984));
    CascadeMux I__6455 (
            .O(N__33984),
            .I(N__33981));
    CascadeBuf I__6454 (
            .O(N__33981),
            .I(N__33978));
    CascadeMux I__6453 (
            .O(N__33978),
            .I(N__33974));
    CascadeMux I__6452 (
            .O(N__33977),
            .I(N__33971));
    CascadeBuf I__6451 (
            .O(N__33974),
            .I(N__33968));
    CascadeBuf I__6450 (
            .O(N__33971),
            .I(N__33965));
    CascadeMux I__6449 (
            .O(N__33968),
            .I(N__33962));
    CascadeMux I__6448 (
            .O(N__33965),
            .I(N__33959));
    CascadeBuf I__6447 (
            .O(N__33962),
            .I(N__33956));
    InMux I__6446 (
            .O(N__33959),
            .I(N__33953));
    CascadeMux I__6445 (
            .O(N__33956),
            .I(N__33950));
    LocalMux I__6444 (
            .O(N__33953),
            .I(N__33947));
    InMux I__6443 (
            .O(N__33950),
            .I(N__33944));
    Span4Mux_v I__6442 (
            .O(N__33947),
            .I(N__33941));
    LocalMux I__6441 (
            .O(N__33944),
            .I(N__33938));
    Sp12to4 I__6440 (
            .O(N__33941),
            .I(N__33934));
    Span4Mux_v I__6439 (
            .O(N__33938),
            .I(N__33931));
    InMux I__6438 (
            .O(N__33937),
            .I(N__33928));
    Span12Mux_h I__6437 (
            .O(N__33934),
            .I(N__33925));
    Sp12to4 I__6436 (
            .O(N__33931),
            .I(N__33922));
    LocalMux I__6435 (
            .O(N__33928),
            .I(data_count_8));
    Odrv12 I__6434 (
            .O(N__33925),
            .I(data_count_8));
    Odrv12 I__6433 (
            .O(N__33922),
            .I(data_count_8));
    InMux I__6432 (
            .O(N__33915),
            .I(bfn_12_19_0_));
    InMux I__6431 (
            .O(N__33912),
            .I(n19773));
    CascadeMux I__6430 (
            .O(N__33909),
            .I(N__33906));
    CascadeBuf I__6429 (
            .O(N__33906),
            .I(N__33903));
    CascadeMux I__6428 (
            .O(N__33903),
            .I(N__33900));
    CascadeBuf I__6427 (
            .O(N__33900),
            .I(N__33897));
    CascadeMux I__6426 (
            .O(N__33897),
            .I(N__33894));
    CascadeBuf I__6425 (
            .O(N__33894),
            .I(N__33891));
    CascadeMux I__6424 (
            .O(N__33891),
            .I(N__33888));
    CascadeBuf I__6423 (
            .O(N__33888),
            .I(N__33885));
    CascadeMux I__6422 (
            .O(N__33885),
            .I(N__33882));
    CascadeBuf I__6421 (
            .O(N__33882),
            .I(N__33879));
    CascadeMux I__6420 (
            .O(N__33879),
            .I(N__33876));
    CascadeBuf I__6419 (
            .O(N__33876),
            .I(N__33873));
    CascadeMux I__6418 (
            .O(N__33873),
            .I(N__33870));
    CascadeBuf I__6417 (
            .O(N__33870),
            .I(N__33867));
    CascadeMux I__6416 (
            .O(N__33867),
            .I(N__33864));
    CascadeBuf I__6415 (
            .O(N__33864),
            .I(N__33860));
    CascadeMux I__6414 (
            .O(N__33863),
            .I(N__33857));
    CascadeMux I__6413 (
            .O(N__33860),
            .I(N__33854));
    CascadeBuf I__6412 (
            .O(N__33857),
            .I(N__33851));
    CascadeBuf I__6411 (
            .O(N__33854),
            .I(N__33848));
    CascadeMux I__6410 (
            .O(N__33851),
            .I(N__33845));
    CascadeMux I__6409 (
            .O(N__33848),
            .I(N__33842));
    InMux I__6408 (
            .O(N__33845),
            .I(N__33839));
    InMux I__6407 (
            .O(N__33842),
            .I(N__33836));
    LocalMux I__6406 (
            .O(N__33839),
            .I(N__33832));
    LocalMux I__6405 (
            .O(N__33836),
            .I(N__33829));
    InMux I__6404 (
            .O(N__33835),
            .I(N__33826));
    Span12Mux_h I__6403 (
            .O(N__33832),
            .I(N__33821));
    Span12Mux_h I__6402 (
            .O(N__33829),
            .I(N__33821));
    LocalMux I__6401 (
            .O(N__33826),
            .I(data_count_9));
    Odrv12 I__6400 (
            .O(N__33821),
            .I(data_count_9));
    InMux I__6399 (
            .O(N__33816),
            .I(N__33813));
    LocalMux I__6398 (
            .O(N__33813),
            .I(\comm_spi.n23089 ));
    InMux I__6397 (
            .O(N__33810),
            .I(N__33807));
    LocalMux I__6396 (
            .O(N__33807),
            .I(N__33804));
    Span4Mux_v I__6395 (
            .O(N__33804),
            .I(N__33800));
    InMux I__6394 (
            .O(N__33803),
            .I(N__33797));
    Span4Mux_h I__6393 (
            .O(N__33800),
            .I(N__33791));
    LocalMux I__6392 (
            .O(N__33797),
            .I(N__33791));
    InMux I__6391 (
            .O(N__33796),
            .I(N__33788));
    Odrv4 I__6390 (
            .O(N__33791),
            .I(cmd_rdadctmp_16));
    LocalMux I__6389 (
            .O(N__33788),
            .I(cmd_rdadctmp_16));
    CascadeMux I__6388 (
            .O(N__33783),
            .I(N__33780));
    InMux I__6387 (
            .O(N__33780),
            .I(N__33777));
    LocalMux I__6386 (
            .O(N__33777),
            .I(N__33773));
    CascadeMux I__6385 (
            .O(N__33776),
            .I(N__33769));
    Span4Mux_h I__6384 (
            .O(N__33773),
            .I(N__33766));
    InMux I__6383 (
            .O(N__33772),
            .I(N__33761));
    InMux I__6382 (
            .O(N__33769),
            .I(N__33761));
    Odrv4 I__6381 (
            .O(N__33766),
            .I(cmd_rdadctmp_17));
    LocalMux I__6380 (
            .O(N__33761),
            .I(cmd_rdadctmp_17));
    CascadeMux I__6379 (
            .O(N__33756),
            .I(N__33753));
    CascadeBuf I__6378 (
            .O(N__33753),
            .I(N__33750));
    CascadeMux I__6377 (
            .O(N__33750),
            .I(N__33747));
    CascadeBuf I__6376 (
            .O(N__33747),
            .I(N__33744));
    CascadeMux I__6375 (
            .O(N__33744),
            .I(N__33741));
    CascadeBuf I__6374 (
            .O(N__33741),
            .I(N__33738));
    CascadeMux I__6373 (
            .O(N__33738),
            .I(N__33735));
    CascadeBuf I__6372 (
            .O(N__33735),
            .I(N__33732));
    CascadeMux I__6371 (
            .O(N__33732),
            .I(N__33729));
    CascadeBuf I__6370 (
            .O(N__33729),
            .I(N__33726));
    CascadeMux I__6369 (
            .O(N__33726),
            .I(N__33723));
    CascadeBuf I__6368 (
            .O(N__33723),
            .I(N__33720));
    CascadeMux I__6367 (
            .O(N__33720),
            .I(N__33717));
    CascadeBuf I__6366 (
            .O(N__33717),
            .I(N__33714));
    CascadeMux I__6365 (
            .O(N__33714),
            .I(N__33710));
    CascadeMux I__6364 (
            .O(N__33713),
            .I(N__33707));
    CascadeBuf I__6363 (
            .O(N__33710),
            .I(N__33704));
    CascadeBuf I__6362 (
            .O(N__33707),
            .I(N__33701));
    CascadeMux I__6361 (
            .O(N__33704),
            .I(N__33698));
    CascadeMux I__6360 (
            .O(N__33701),
            .I(N__33695));
    CascadeBuf I__6359 (
            .O(N__33698),
            .I(N__33692));
    InMux I__6358 (
            .O(N__33695),
            .I(N__33689));
    CascadeMux I__6357 (
            .O(N__33692),
            .I(N__33686));
    LocalMux I__6356 (
            .O(N__33689),
            .I(N__33683));
    InMux I__6355 (
            .O(N__33686),
            .I(N__33680));
    Span4Mux_h I__6354 (
            .O(N__33683),
            .I(N__33677));
    LocalMux I__6353 (
            .O(N__33680),
            .I(N__33674));
    Sp12to4 I__6352 (
            .O(N__33677),
            .I(N__33670));
    Span4Mux_v I__6351 (
            .O(N__33674),
            .I(N__33667));
    InMux I__6350 (
            .O(N__33673),
            .I(N__33664));
    Span12Mux_v I__6349 (
            .O(N__33670),
            .I(N__33659));
    Sp12to4 I__6348 (
            .O(N__33667),
            .I(N__33659));
    LocalMux I__6347 (
            .O(N__33664),
            .I(data_count_0));
    Odrv12 I__6346 (
            .O(N__33659),
            .I(data_count_0));
    CascadeMux I__6345 (
            .O(N__33654),
            .I(N__33651));
    CascadeBuf I__6344 (
            .O(N__33651),
            .I(N__33648));
    CascadeMux I__6343 (
            .O(N__33648),
            .I(N__33645));
    CascadeBuf I__6342 (
            .O(N__33645),
            .I(N__33642));
    CascadeMux I__6341 (
            .O(N__33642),
            .I(N__33639));
    CascadeBuf I__6340 (
            .O(N__33639),
            .I(N__33636));
    CascadeMux I__6339 (
            .O(N__33636),
            .I(N__33633));
    CascadeBuf I__6338 (
            .O(N__33633),
            .I(N__33630));
    CascadeMux I__6337 (
            .O(N__33630),
            .I(N__33627));
    CascadeBuf I__6336 (
            .O(N__33627),
            .I(N__33624));
    CascadeMux I__6335 (
            .O(N__33624),
            .I(N__33621));
    CascadeBuf I__6334 (
            .O(N__33621),
            .I(N__33618));
    CascadeMux I__6333 (
            .O(N__33618),
            .I(N__33615));
    CascadeBuf I__6332 (
            .O(N__33615),
            .I(N__33612));
    CascadeMux I__6331 (
            .O(N__33612),
            .I(N__33608));
    CascadeMux I__6330 (
            .O(N__33611),
            .I(N__33605));
    CascadeBuf I__6329 (
            .O(N__33608),
            .I(N__33602));
    CascadeBuf I__6328 (
            .O(N__33605),
            .I(N__33599));
    CascadeMux I__6327 (
            .O(N__33602),
            .I(N__33596));
    CascadeMux I__6326 (
            .O(N__33599),
            .I(N__33593));
    CascadeBuf I__6325 (
            .O(N__33596),
            .I(N__33590));
    InMux I__6324 (
            .O(N__33593),
            .I(N__33587));
    CascadeMux I__6323 (
            .O(N__33590),
            .I(N__33584));
    LocalMux I__6322 (
            .O(N__33587),
            .I(N__33581));
    InMux I__6321 (
            .O(N__33584),
            .I(N__33578));
    Span4Mux_v I__6320 (
            .O(N__33581),
            .I(N__33575));
    LocalMux I__6319 (
            .O(N__33578),
            .I(N__33572));
    Sp12to4 I__6318 (
            .O(N__33575),
            .I(N__33568));
    Span4Mux_v I__6317 (
            .O(N__33572),
            .I(N__33565));
    InMux I__6316 (
            .O(N__33571),
            .I(N__33562));
    Span12Mux_h I__6315 (
            .O(N__33568),
            .I(N__33559));
    Sp12to4 I__6314 (
            .O(N__33565),
            .I(N__33556));
    LocalMux I__6313 (
            .O(N__33562),
            .I(data_count_1));
    Odrv12 I__6312 (
            .O(N__33559),
            .I(data_count_1));
    Odrv12 I__6311 (
            .O(N__33556),
            .I(data_count_1));
    InMux I__6310 (
            .O(N__33549),
            .I(n19765));
    CascadeMux I__6309 (
            .O(N__33546),
            .I(N__33543));
    CascadeBuf I__6308 (
            .O(N__33543),
            .I(N__33540));
    CascadeMux I__6307 (
            .O(N__33540),
            .I(N__33537));
    CascadeBuf I__6306 (
            .O(N__33537),
            .I(N__33534));
    CascadeMux I__6305 (
            .O(N__33534),
            .I(N__33531));
    CascadeBuf I__6304 (
            .O(N__33531),
            .I(N__33528));
    CascadeMux I__6303 (
            .O(N__33528),
            .I(N__33525));
    CascadeBuf I__6302 (
            .O(N__33525),
            .I(N__33522));
    CascadeMux I__6301 (
            .O(N__33522),
            .I(N__33519));
    CascadeBuf I__6300 (
            .O(N__33519),
            .I(N__33516));
    CascadeMux I__6299 (
            .O(N__33516),
            .I(N__33513));
    CascadeBuf I__6298 (
            .O(N__33513),
            .I(N__33510));
    CascadeMux I__6297 (
            .O(N__33510),
            .I(N__33507));
    CascadeBuf I__6296 (
            .O(N__33507),
            .I(N__33504));
    CascadeMux I__6295 (
            .O(N__33504),
            .I(N__33501));
    CascadeBuf I__6294 (
            .O(N__33501),
            .I(N__33497));
    CascadeMux I__6293 (
            .O(N__33500),
            .I(N__33494));
    CascadeMux I__6292 (
            .O(N__33497),
            .I(N__33491));
    CascadeBuf I__6291 (
            .O(N__33494),
            .I(N__33488));
    CascadeBuf I__6290 (
            .O(N__33491),
            .I(N__33485));
    CascadeMux I__6289 (
            .O(N__33488),
            .I(N__33482));
    CascadeMux I__6288 (
            .O(N__33485),
            .I(N__33479));
    InMux I__6287 (
            .O(N__33482),
            .I(N__33476));
    InMux I__6286 (
            .O(N__33479),
            .I(N__33473));
    LocalMux I__6285 (
            .O(N__33476),
            .I(N__33470));
    LocalMux I__6284 (
            .O(N__33473),
            .I(N__33467));
    Span4Mux_h I__6283 (
            .O(N__33470),
            .I(N__33464));
    Span4Mux_v I__6282 (
            .O(N__33467),
            .I(N__33461));
    Sp12to4 I__6281 (
            .O(N__33464),
            .I(N__33457));
    Span4Mux_h I__6280 (
            .O(N__33461),
            .I(N__33454));
    InMux I__6279 (
            .O(N__33460),
            .I(N__33451));
    Span12Mux_v I__6278 (
            .O(N__33457),
            .I(N__33448));
    Span4Mux_h I__6277 (
            .O(N__33454),
            .I(N__33445));
    LocalMux I__6276 (
            .O(N__33451),
            .I(data_count_2));
    Odrv12 I__6275 (
            .O(N__33448),
            .I(data_count_2));
    Odrv4 I__6274 (
            .O(N__33445),
            .I(data_count_2));
    InMux I__6273 (
            .O(N__33438),
            .I(n19766));
    CascadeMux I__6272 (
            .O(N__33435),
            .I(N__33432));
    CascadeBuf I__6271 (
            .O(N__33432),
            .I(N__33429));
    CascadeMux I__6270 (
            .O(N__33429),
            .I(N__33426));
    CascadeBuf I__6269 (
            .O(N__33426),
            .I(N__33423));
    CascadeMux I__6268 (
            .O(N__33423),
            .I(N__33420));
    CascadeBuf I__6267 (
            .O(N__33420),
            .I(N__33417));
    CascadeMux I__6266 (
            .O(N__33417),
            .I(N__33414));
    CascadeBuf I__6265 (
            .O(N__33414),
            .I(N__33411));
    CascadeMux I__6264 (
            .O(N__33411),
            .I(N__33408));
    CascadeBuf I__6263 (
            .O(N__33408),
            .I(N__33405));
    CascadeMux I__6262 (
            .O(N__33405),
            .I(N__33402));
    CascadeBuf I__6261 (
            .O(N__33402),
            .I(N__33399));
    CascadeMux I__6260 (
            .O(N__33399),
            .I(N__33396));
    CascadeBuf I__6259 (
            .O(N__33396),
            .I(N__33393));
    CascadeMux I__6258 (
            .O(N__33393),
            .I(N__33390));
    CascadeBuf I__6257 (
            .O(N__33390),
            .I(N__33386));
    CascadeMux I__6256 (
            .O(N__33389),
            .I(N__33383));
    CascadeMux I__6255 (
            .O(N__33386),
            .I(N__33380));
    CascadeBuf I__6254 (
            .O(N__33383),
            .I(N__33377));
    CascadeBuf I__6253 (
            .O(N__33380),
            .I(N__33374));
    CascadeMux I__6252 (
            .O(N__33377),
            .I(N__33371));
    CascadeMux I__6251 (
            .O(N__33374),
            .I(N__33368));
    InMux I__6250 (
            .O(N__33371),
            .I(N__33365));
    InMux I__6249 (
            .O(N__33368),
            .I(N__33362));
    LocalMux I__6248 (
            .O(N__33365),
            .I(N__33359));
    LocalMux I__6247 (
            .O(N__33362),
            .I(N__33356));
    Span4Mux_h I__6246 (
            .O(N__33359),
            .I(N__33353));
    Span4Mux_v I__6245 (
            .O(N__33356),
            .I(N__33350));
    Span4Mux_h I__6244 (
            .O(N__33353),
            .I(N__33346));
    Span4Mux_h I__6243 (
            .O(N__33350),
            .I(N__33343));
    InMux I__6242 (
            .O(N__33349),
            .I(N__33340));
    Sp12to4 I__6241 (
            .O(N__33346),
            .I(N__33337));
    Span4Mux_h I__6240 (
            .O(N__33343),
            .I(N__33334));
    LocalMux I__6239 (
            .O(N__33340),
            .I(data_count_3));
    Odrv12 I__6238 (
            .O(N__33337),
            .I(data_count_3));
    Odrv4 I__6237 (
            .O(N__33334),
            .I(data_count_3));
    InMux I__6236 (
            .O(N__33327),
            .I(n19767));
    CascadeMux I__6235 (
            .O(N__33324),
            .I(N__33321));
    CascadeBuf I__6234 (
            .O(N__33321),
            .I(N__33318));
    CascadeMux I__6233 (
            .O(N__33318),
            .I(N__33315));
    CascadeBuf I__6232 (
            .O(N__33315),
            .I(N__33312));
    CascadeMux I__6231 (
            .O(N__33312),
            .I(N__33309));
    CascadeBuf I__6230 (
            .O(N__33309),
            .I(N__33306));
    CascadeMux I__6229 (
            .O(N__33306),
            .I(N__33303));
    CascadeBuf I__6228 (
            .O(N__33303),
            .I(N__33300));
    CascadeMux I__6227 (
            .O(N__33300),
            .I(N__33297));
    CascadeBuf I__6226 (
            .O(N__33297),
            .I(N__33294));
    CascadeMux I__6225 (
            .O(N__33294),
            .I(N__33291));
    CascadeBuf I__6224 (
            .O(N__33291),
            .I(N__33288));
    CascadeMux I__6223 (
            .O(N__33288),
            .I(N__33285));
    CascadeBuf I__6222 (
            .O(N__33285),
            .I(N__33282));
    CascadeMux I__6221 (
            .O(N__33282),
            .I(N__33279));
    CascadeBuf I__6220 (
            .O(N__33279),
            .I(N__33276));
    CascadeMux I__6219 (
            .O(N__33276),
            .I(N__33272));
    CascadeMux I__6218 (
            .O(N__33275),
            .I(N__33269));
    CascadeBuf I__6217 (
            .O(N__33272),
            .I(N__33266));
    CascadeBuf I__6216 (
            .O(N__33269),
            .I(N__33263));
    CascadeMux I__6215 (
            .O(N__33266),
            .I(N__33260));
    CascadeMux I__6214 (
            .O(N__33263),
            .I(N__33257));
    InMux I__6213 (
            .O(N__33260),
            .I(N__33254));
    InMux I__6212 (
            .O(N__33257),
            .I(N__33251));
    LocalMux I__6211 (
            .O(N__33254),
            .I(N__33248));
    LocalMux I__6210 (
            .O(N__33251),
            .I(N__33244));
    Span4Mux_v I__6209 (
            .O(N__33248),
            .I(N__33241));
    InMux I__6208 (
            .O(N__33247),
            .I(N__33238));
    Span12Mux_v I__6207 (
            .O(N__33244),
            .I(N__33235));
    Sp12to4 I__6206 (
            .O(N__33241),
            .I(N__33232));
    LocalMux I__6205 (
            .O(N__33238),
            .I(data_count_4));
    Odrv12 I__6204 (
            .O(N__33235),
            .I(data_count_4));
    Odrv12 I__6203 (
            .O(N__33232),
            .I(data_count_4));
    InMux I__6202 (
            .O(N__33225),
            .I(n19768));
    CascadeMux I__6201 (
            .O(N__33222),
            .I(N__33219));
    CascadeBuf I__6200 (
            .O(N__33219),
            .I(N__33216));
    CascadeMux I__6199 (
            .O(N__33216),
            .I(N__33213));
    CascadeBuf I__6198 (
            .O(N__33213),
            .I(N__33210));
    CascadeMux I__6197 (
            .O(N__33210),
            .I(N__33207));
    CascadeBuf I__6196 (
            .O(N__33207),
            .I(N__33204));
    CascadeMux I__6195 (
            .O(N__33204),
            .I(N__33201));
    CascadeBuf I__6194 (
            .O(N__33201),
            .I(N__33198));
    CascadeMux I__6193 (
            .O(N__33198),
            .I(N__33195));
    CascadeBuf I__6192 (
            .O(N__33195),
            .I(N__33192));
    CascadeMux I__6191 (
            .O(N__33192),
            .I(N__33189));
    CascadeBuf I__6190 (
            .O(N__33189),
            .I(N__33186));
    CascadeMux I__6189 (
            .O(N__33186),
            .I(N__33183));
    CascadeBuf I__6188 (
            .O(N__33183),
            .I(N__33179));
    CascadeMux I__6187 (
            .O(N__33182),
            .I(N__33176));
    CascadeMux I__6186 (
            .O(N__33179),
            .I(N__33173));
    CascadeBuf I__6185 (
            .O(N__33176),
            .I(N__33170));
    CascadeBuf I__6184 (
            .O(N__33173),
            .I(N__33167));
    CascadeMux I__6183 (
            .O(N__33170),
            .I(N__33164));
    CascadeMux I__6182 (
            .O(N__33167),
            .I(N__33161));
    InMux I__6181 (
            .O(N__33164),
            .I(N__33158));
    CascadeBuf I__6180 (
            .O(N__33161),
            .I(N__33155));
    LocalMux I__6179 (
            .O(N__33158),
            .I(N__33152));
    CascadeMux I__6178 (
            .O(N__33155),
            .I(N__33149));
    Span4Mux_v I__6177 (
            .O(N__33152),
            .I(N__33146));
    InMux I__6176 (
            .O(N__33149),
            .I(N__33143));
    Sp12to4 I__6175 (
            .O(N__33146),
            .I(N__33139));
    LocalMux I__6174 (
            .O(N__33143),
            .I(N__33136));
    InMux I__6173 (
            .O(N__33142),
            .I(N__33133));
    Span12Mux_h I__6172 (
            .O(N__33139),
            .I(N__33130));
    Span4Mux_v I__6171 (
            .O(N__33136),
            .I(N__33127));
    LocalMux I__6170 (
            .O(N__33133),
            .I(N__33120));
    Span12Mux_v I__6169 (
            .O(N__33130),
            .I(N__33120));
    Sp12to4 I__6168 (
            .O(N__33127),
            .I(N__33120));
    Odrv12 I__6167 (
            .O(N__33120),
            .I(data_count_5));
    InMux I__6166 (
            .O(N__33117),
            .I(n19769));
    CascadeMux I__6165 (
            .O(N__33114),
            .I(N__33110));
    InMux I__6164 (
            .O(N__33113),
            .I(N__33107));
    InMux I__6163 (
            .O(N__33110),
            .I(N__33104));
    LocalMux I__6162 (
            .O(N__33107),
            .I(N__33101));
    LocalMux I__6161 (
            .O(N__33104),
            .I(N__33098));
    Span4Mux_v I__6160 (
            .O(N__33101),
            .I(N__33092));
    Span4Mux_v I__6159 (
            .O(N__33098),
            .I(N__33092));
    InMux I__6158 (
            .O(N__33097),
            .I(N__33089));
    Odrv4 I__6157 (
            .O(N__33092),
            .I(cmd_rdadctmp_21));
    LocalMux I__6156 (
            .O(N__33089),
            .I(cmd_rdadctmp_21));
    CascadeMux I__6155 (
            .O(N__33084),
            .I(N__33080));
    CascadeMux I__6154 (
            .O(N__33083),
            .I(N__33076));
    InMux I__6153 (
            .O(N__33080),
            .I(N__33073));
    InMux I__6152 (
            .O(N__33079),
            .I(N__33070));
    InMux I__6151 (
            .O(N__33076),
            .I(N__33067));
    LocalMux I__6150 (
            .O(N__33073),
            .I(N__33064));
    LocalMux I__6149 (
            .O(N__33070),
            .I(N__33061));
    LocalMux I__6148 (
            .O(N__33067),
            .I(N__33056));
    Span4Mux_v I__6147 (
            .O(N__33064),
            .I(N__33056));
    Span12Mux_h I__6146 (
            .O(N__33061),
            .I(N__33053));
    Odrv4 I__6145 (
            .O(N__33056),
            .I(buf_adcdata_iac_13));
    Odrv12 I__6144 (
            .O(N__33053),
            .I(buf_adcdata_iac_13));
    InMux I__6143 (
            .O(N__33048),
            .I(N__33045));
    LocalMux I__6142 (
            .O(N__33045),
            .I(N__33042));
    Span12Mux_h I__6141 (
            .O(N__33042),
            .I(N__33037));
    InMux I__6140 (
            .O(N__33041),
            .I(N__33032));
    InMux I__6139 (
            .O(N__33040),
            .I(N__33032));
    Odrv12 I__6138 (
            .O(N__33037),
            .I(acadc_skipCount_13));
    LocalMux I__6137 (
            .O(N__33032),
            .I(acadc_skipCount_13));
    InMux I__6136 (
            .O(N__33027),
            .I(N__33024));
    LocalMux I__6135 (
            .O(N__33024),
            .I(N__33020));
    InMux I__6134 (
            .O(N__33023),
            .I(N__33017));
    Sp12to4 I__6133 (
            .O(N__33020),
            .I(N__33013));
    LocalMux I__6132 (
            .O(N__33017),
            .I(N__33010));
    InMux I__6131 (
            .O(N__33016),
            .I(N__33007));
    Span12Mux_v I__6130 (
            .O(N__33013),
            .I(N__33004));
    Odrv4 I__6129 (
            .O(N__33010),
            .I(buf_dds0_5));
    LocalMux I__6128 (
            .O(N__33007),
            .I(buf_dds0_5));
    Odrv12 I__6127 (
            .O(N__33004),
            .I(buf_dds0_5));
    InMux I__6126 (
            .O(N__32997),
            .I(N__32992));
    InMux I__6125 (
            .O(N__32996),
            .I(N__32989));
    InMux I__6124 (
            .O(N__32995),
            .I(N__32986));
    LocalMux I__6123 (
            .O(N__32992),
            .I(N__32983));
    LocalMux I__6122 (
            .O(N__32989),
            .I(buf_dds0_3));
    LocalMux I__6121 (
            .O(N__32986),
            .I(buf_dds0_3));
    Odrv4 I__6120 (
            .O(N__32983),
            .I(buf_dds0_3));
    InMux I__6119 (
            .O(N__32976),
            .I(N__32972));
    InMux I__6118 (
            .O(N__32975),
            .I(N__32968));
    LocalMux I__6117 (
            .O(N__32972),
            .I(N__32965));
    InMux I__6116 (
            .O(N__32971),
            .I(N__32962));
    LocalMux I__6115 (
            .O(N__32968),
            .I(acadc_skipCount_5));
    Odrv12 I__6114 (
            .O(N__32965),
            .I(acadc_skipCount_5));
    LocalMux I__6113 (
            .O(N__32962),
            .I(acadc_skipCount_5));
    InMux I__6112 (
            .O(N__32955),
            .I(N__32952));
    LocalMux I__6111 (
            .O(N__32952),
            .I(n20_adj_1670));
    CascadeMux I__6110 (
            .O(N__32949),
            .I(n8_adj_1560_cascade_));
    CascadeMux I__6109 (
            .O(N__32946),
            .I(N__32943));
    CascadeBuf I__6108 (
            .O(N__32943),
            .I(N__32940));
    CascadeMux I__6107 (
            .O(N__32940),
            .I(N__32937));
    CascadeBuf I__6106 (
            .O(N__32937),
            .I(N__32934));
    CascadeMux I__6105 (
            .O(N__32934),
            .I(N__32931));
    CascadeBuf I__6104 (
            .O(N__32931),
            .I(N__32928));
    CascadeMux I__6103 (
            .O(N__32928),
            .I(N__32925));
    CascadeBuf I__6102 (
            .O(N__32925),
            .I(N__32922));
    CascadeMux I__6101 (
            .O(N__32922),
            .I(N__32919));
    CascadeBuf I__6100 (
            .O(N__32919),
            .I(N__32916));
    CascadeMux I__6099 (
            .O(N__32916),
            .I(N__32913));
    CascadeBuf I__6098 (
            .O(N__32913),
            .I(N__32910));
    CascadeMux I__6097 (
            .O(N__32910),
            .I(N__32907));
    CascadeBuf I__6096 (
            .O(N__32907),
            .I(N__32904));
    CascadeMux I__6095 (
            .O(N__32904),
            .I(N__32901));
    CascadeBuf I__6094 (
            .O(N__32901),
            .I(N__32897));
    CascadeMux I__6093 (
            .O(N__32900),
            .I(N__32894));
    CascadeMux I__6092 (
            .O(N__32897),
            .I(N__32891));
    CascadeBuf I__6091 (
            .O(N__32894),
            .I(N__32888));
    CascadeBuf I__6090 (
            .O(N__32891),
            .I(N__32885));
    CascadeMux I__6089 (
            .O(N__32888),
            .I(N__32882));
    CascadeMux I__6088 (
            .O(N__32885),
            .I(N__32879));
    InMux I__6087 (
            .O(N__32882),
            .I(N__32876));
    InMux I__6086 (
            .O(N__32879),
            .I(N__32873));
    LocalMux I__6085 (
            .O(N__32876),
            .I(N__32870));
    LocalMux I__6084 (
            .O(N__32873),
            .I(N__32867));
    Span4Mux_h I__6083 (
            .O(N__32870),
            .I(N__32864));
    Span4Mux_h I__6082 (
            .O(N__32867),
            .I(N__32861));
    Span4Mux_v I__6081 (
            .O(N__32864),
            .I(N__32858));
    Span4Mux_h I__6080 (
            .O(N__32861),
            .I(N__32855));
    Span4Mux_h I__6079 (
            .O(N__32858),
            .I(N__32852));
    Span4Mux_v I__6078 (
            .O(N__32855),
            .I(N__32849));
    Odrv4 I__6077 (
            .O(N__32852),
            .I(data_index_9_N_212_7));
    Odrv4 I__6076 (
            .O(N__32849),
            .I(data_index_9_N_212_7));
    InMux I__6075 (
            .O(N__32844),
            .I(N__32841));
    LocalMux I__6074 (
            .O(N__32841),
            .I(n24_adj_1593));
    InMux I__6073 (
            .O(N__32838),
            .I(N__32835));
    LocalMux I__6072 (
            .O(N__32835),
            .I(N__32832));
    Odrv12 I__6071 (
            .O(N__32832),
            .I(n23_adj_1591));
    CascadeMux I__6070 (
            .O(N__32829),
            .I(n22_adj_1590_cascade_));
    InMux I__6069 (
            .O(N__32826),
            .I(N__32823));
    LocalMux I__6068 (
            .O(N__32823),
            .I(n18));
    CascadeMux I__6067 (
            .O(N__32820),
            .I(n30_adj_1543_cascade_));
    InMux I__6066 (
            .O(N__32817),
            .I(N__32810));
    InMux I__6065 (
            .O(N__32816),
            .I(N__32810));
    InMux I__6064 (
            .O(N__32815),
            .I(N__32807));
    LocalMux I__6063 (
            .O(N__32810),
            .I(N__32804));
    LocalMux I__6062 (
            .O(N__32807),
            .I(N__32801));
    Odrv4 I__6061 (
            .O(N__32804),
            .I(n31_adj_1537));
    Odrv4 I__6060 (
            .O(N__32801),
            .I(n31_adj_1537));
    CascadeMux I__6059 (
            .O(N__32796),
            .I(N__32793));
    InMux I__6058 (
            .O(N__32793),
            .I(N__32790));
    LocalMux I__6057 (
            .O(N__32790),
            .I(N__32787));
    Span4Mux_v I__6056 (
            .O(N__32787),
            .I(N__32783));
    CascadeMux I__6055 (
            .O(N__32786),
            .I(N__32780));
    Span4Mux_h I__6054 (
            .O(N__32783),
            .I(N__32776));
    InMux I__6053 (
            .O(N__32780),
            .I(N__32773));
    InMux I__6052 (
            .O(N__32779),
            .I(N__32770));
    Odrv4 I__6051 (
            .O(N__32776),
            .I(cmd_rdadctmp_26));
    LocalMux I__6050 (
            .O(N__32773),
            .I(cmd_rdadctmp_26));
    LocalMux I__6049 (
            .O(N__32770),
            .I(cmd_rdadctmp_26));
    InMux I__6048 (
            .O(N__32763),
            .I(N__32760));
    LocalMux I__6047 (
            .O(N__32760),
            .I(N__32757));
    Span4Mux_v I__6046 (
            .O(N__32757),
            .I(N__32753));
    InMux I__6045 (
            .O(N__32756),
            .I(N__32750));
    Span4Mux_h I__6044 (
            .O(N__32753),
            .I(N__32746));
    LocalMux I__6043 (
            .O(N__32750),
            .I(N__32743));
    InMux I__6042 (
            .O(N__32749),
            .I(N__32740));
    Span4Mux_h I__6041 (
            .O(N__32746),
            .I(N__32737));
    Span4Mux_v I__6040 (
            .O(N__32743),
            .I(N__32734));
    LocalMux I__6039 (
            .O(N__32740),
            .I(buf_adcdata_iac_18));
    Odrv4 I__6038 (
            .O(N__32737),
            .I(buf_adcdata_iac_18));
    Odrv4 I__6037 (
            .O(N__32734),
            .I(buf_adcdata_iac_18));
    InMux I__6036 (
            .O(N__32727),
            .I(N__32723));
    InMux I__6035 (
            .O(N__32726),
            .I(N__32720));
    LocalMux I__6034 (
            .O(N__32723),
            .I(N__32716));
    LocalMux I__6033 (
            .O(N__32720),
            .I(N__32713));
    InMux I__6032 (
            .O(N__32719),
            .I(N__32710));
    Span4Mux_v I__6031 (
            .O(N__32716),
            .I(N__32707));
    Span4Mux_h I__6030 (
            .O(N__32713),
            .I(N__32704));
    LocalMux I__6029 (
            .O(N__32710),
            .I(acadc_skipCount_8));
    Odrv4 I__6028 (
            .O(N__32707),
            .I(acadc_skipCount_8));
    Odrv4 I__6027 (
            .O(N__32704),
            .I(acadc_skipCount_8));
    CascadeMux I__6026 (
            .O(N__32697),
            .I(n14_adj_1538_cascade_));
    InMux I__6025 (
            .O(N__32694),
            .I(N__32691));
    LocalMux I__6024 (
            .O(N__32691),
            .I(n26_adj_1525));
    InMux I__6023 (
            .O(N__32688),
            .I(N__32684));
    InMux I__6022 (
            .O(N__32687),
            .I(N__32680));
    LocalMux I__6021 (
            .O(N__32684),
            .I(N__32677));
    InMux I__6020 (
            .O(N__32683),
            .I(N__32674));
    LocalMux I__6019 (
            .O(N__32680),
            .I(buf_dds1_3));
    Odrv12 I__6018 (
            .O(N__32677),
            .I(buf_dds1_3));
    LocalMux I__6017 (
            .O(N__32674),
            .I(buf_dds1_3));
    InMux I__6016 (
            .O(N__32667),
            .I(N__32664));
    LocalMux I__6015 (
            .O(N__32664),
            .I(N__32661));
    Span4Mux_h I__6014 (
            .O(N__32661),
            .I(N__32656));
    InMux I__6013 (
            .O(N__32660),
            .I(N__32651));
    InMux I__6012 (
            .O(N__32659),
            .I(N__32651));
    Odrv4 I__6011 (
            .O(N__32656),
            .I(acadc_skipCount_4));
    LocalMux I__6010 (
            .O(N__32651),
            .I(acadc_skipCount_4));
    InMux I__6009 (
            .O(N__32646),
            .I(N__32643));
    LocalMux I__6008 (
            .O(N__32643),
            .I(n8_adj_1560));
    CascadeMux I__6007 (
            .O(N__32640),
            .I(n30_adj_1631_cascade_));
    InMux I__6006 (
            .O(N__32637),
            .I(N__32634));
    LocalMux I__6005 (
            .O(N__32634),
            .I(N__32631));
    Sp12to4 I__6004 (
            .O(N__32631),
            .I(N__32628));
    Odrv12 I__6003 (
            .O(N__32628),
            .I(n9));
    InMux I__6002 (
            .O(N__32625),
            .I(N__32622));
    LocalMux I__6001 (
            .O(N__32622),
            .I(N__32619));
    Span4Mux_v I__6000 (
            .O(N__32619),
            .I(N__32616));
    Span4Mux_h I__5999 (
            .O(N__32616),
            .I(N__32613));
    Span4Mux_h I__5998 (
            .O(N__32613),
            .I(N__32610));
    Span4Mux_v I__5997 (
            .O(N__32610),
            .I(N__32607));
    Odrv4 I__5996 (
            .O(N__32607),
            .I(buf_data_iac_22));
    CascadeMux I__5995 (
            .O(N__32604),
            .I(N__32601));
    InMux I__5994 (
            .O(N__32601),
            .I(N__32597));
    CascadeMux I__5993 (
            .O(N__32600),
            .I(N__32594));
    LocalMux I__5992 (
            .O(N__32597),
            .I(N__32591));
    InMux I__5991 (
            .O(N__32594),
            .I(N__32588));
    Span4Mux_h I__5990 (
            .O(N__32591),
            .I(N__32585));
    LocalMux I__5989 (
            .O(N__32588),
            .I(data_idxvec_14));
    Odrv4 I__5988 (
            .O(N__32585),
            .I(data_idxvec_14));
    CascadeMux I__5987 (
            .O(N__32580),
            .I(N__32577));
    InMux I__5986 (
            .O(N__32577),
            .I(N__32574));
    LocalMux I__5985 (
            .O(N__32574),
            .I(N__32571));
    Span4Mux_v I__5984 (
            .O(N__32571),
            .I(N__32568));
    Span4Mux_h I__5983 (
            .O(N__32568),
            .I(N__32565));
    Odrv4 I__5982 (
            .O(N__32565),
            .I(n21330));
    CascadeMux I__5981 (
            .O(N__32562),
            .I(N__32558));
    InMux I__5980 (
            .O(N__32561),
            .I(N__32555));
    InMux I__5979 (
            .O(N__32558),
            .I(N__32551));
    LocalMux I__5978 (
            .O(N__32555),
            .I(N__32548));
    InMux I__5977 (
            .O(N__32554),
            .I(N__32545));
    LocalMux I__5976 (
            .O(N__32551),
            .I(acadc_skipCount_11));
    Odrv4 I__5975 (
            .O(N__32548),
            .I(acadc_skipCount_11));
    LocalMux I__5974 (
            .O(N__32545),
            .I(acadc_skipCount_11));
    CascadeMux I__5973 (
            .O(N__32538),
            .I(N__32535));
    InMux I__5972 (
            .O(N__32535),
            .I(N__32532));
    LocalMux I__5971 (
            .O(N__32532),
            .I(N__32529));
    Odrv4 I__5970 (
            .O(N__32529),
            .I(n23_adj_1677));
    InMux I__5969 (
            .O(N__32526),
            .I(N__32522));
    InMux I__5968 (
            .O(N__32525),
            .I(N__32519));
    LocalMux I__5967 (
            .O(N__32522),
            .I(N__32513));
    LocalMux I__5966 (
            .O(N__32519),
            .I(N__32513));
    InMux I__5965 (
            .O(N__32518),
            .I(N__32510));
    Span4Mux_v I__5964 (
            .O(N__32513),
            .I(N__32507));
    LocalMux I__5963 (
            .O(N__32510),
            .I(N__32502));
    Span4Mux_h I__5962 (
            .O(N__32507),
            .I(N__32502));
    Odrv4 I__5961 (
            .O(N__32502),
            .I(buf_dds1_9));
    InMux I__5960 (
            .O(N__32499),
            .I(N__32496));
    LocalMux I__5959 (
            .O(N__32496),
            .I(N__32493));
    Span4Mux_v I__5958 (
            .O(N__32493),
            .I(N__32490));
    Span4Mux_v I__5957 (
            .O(N__32490),
            .I(N__32486));
    CascadeMux I__5956 (
            .O(N__32489),
            .I(N__32483));
    Span4Mux_h I__5955 (
            .O(N__32486),
            .I(N__32480));
    InMux I__5954 (
            .O(N__32483),
            .I(N__32477));
    Odrv4 I__5953 (
            .O(N__32480),
            .I(buf_adcdata_vdc_14));
    LocalMux I__5952 (
            .O(N__32477),
            .I(buf_adcdata_vdc_14));
    InMux I__5951 (
            .O(N__32472),
            .I(N__32469));
    LocalMux I__5950 (
            .O(N__32469),
            .I(N__32465));
    InMux I__5949 (
            .O(N__32468),
            .I(N__32462));
    Span12Mux_v I__5948 (
            .O(N__32465),
            .I(N__32458));
    LocalMux I__5947 (
            .O(N__32462),
            .I(N__32455));
    InMux I__5946 (
            .O(N__32461),
            .I(N__32452));
    Span12Mux_h I__5945 (
            .O(N__32458),
            .I(N__32449));
    Span4Mux_h I__5944 (
            .O(N__32455),
            .I(N__32446));
    LocalMux I__5943 (
            .O(N__32452),
            .I(buf_adcdata_vac_14));
    Odrv12 I__5942 (
            .O(N__32449),
            .I(buf_adcdata_vac_14));
    Odrv4 I__5941 (
            .O(N__32446),
            .I(buf_adcdata_vac_14));
    InMux I__5940 (
            .O(N__32439),
            .I(N__32436));
    LocalMux I__5939 (
            .O(N__32436),
            .I(N__32433));
    Odrv4 I__5938 (
            .O(N__32433),
            .I(n20));
    CascadeMux I__5937 (
            .O(N__32430),
            .I(n17_cascade_));
    InMux I__5936 (
            .O(N__32427),
            .I(N__32424));
    LocalMux I__5935 (
            .O(N__32424),
            .I(n19_adj_1526));
    InMux I__5934 (
            .O(N__32421),
            .I(N__32415));
    InMux I__5933 (
            .O(N__32420),
            .I(N__32415));
    LocalMux I__5932 (
            .O(N__32415),
            .I(n29));
    InMux I__5931 (
            .O(N__32412),
            .I(N__32408));
    CascadeMux I__5930 (
            .O(N__32411),
            .I(N__32405));
    LocalMux I__5929 (
            .O(N__32408),
            .I(N__32402));
    InMux I__5928 (
            .O(N__32405),
            .I(N__32399));
    Span4Mux_v I__5927 (
            .O(N__32402),
            .I(N__32396));
    LocalMux I__5926 (
            .O(N__32399),
            .I(data_idxvec_13));
    Odrv4 I__5925 (
            .O(N__32396),
            .I(data_idxvec_13));
    CascadeMux I__5924 (
            .O(N__32391),
            .I(N__32387));
    InMux I__5923 (
            .O(N__32390),
            .I(N__32384));
    InMux I__5922 (
            .O(N__32387),
            .I(N__32381));
    LocalMux I__5921 (
            .O(N__32384),
            .I(N__32378));
    LocalMux I__5920 (
            .O(N__32381),
            .I(N__32372));
    Span4Mux_h I__5919 (
            .O(N__32378),
            .I(N__32372));
    InMux I__5918 (
            .O(N__32377),
            .I(N__32369));
    Odrv4 I__5917 (
            .O(N__32372),
            .I(comm_cmd_4));
    LocalMux I__5916 (
            .O(N__32369),
            .I(comm_cmd_4));
    CascadeMux I__5915 (
            .O(N__32364),
            .I(n16818_cascade_));
    InMux I__5914 (
            .O(N__32361),
            .I(N__32358));
    LocalMux I__5913 (
            .O(N__32358),
            .I(N__32355));
    Span4Mux_v I__5912 (
            .O(N__32355),
            .I(N__32352));
    Span4Mux_h I__5911 (
            .O(N__32352),
            .I(N__32349));
    Odrv4 I__5910 (
            .O(N__32349),
            .I(n16_adj_1628));
    InMux I__5909 (
            .O(N__32346),
            .I(N__32343));
    LocalMux I__5908 (
            .O(N__32343),
            .I(N__32340));
    Span4Mux_h I__5907 (
            .O(N__32340),
            .I(N__32337));
    Odrv4 I__5906 (
            .O(N__32337),
            .I(n22365));
    InMux I__5905 (
            .O(N__32334),
            .I(N__32331));
    LocalMux I__5904 (
            .O(N__32331),
            .I(N__32328));
    Span4Mux_v I__5903 (
            .O(N__32328),
            .I(N__32324));
    InMux I__5902 (
            .O(N__32327),
            .I(N__32321));
    Span4Mux_h I__5901 (
            .O(N__32324),
            .I(N__32318));
    LocalMux I__5900 (
            .O(N__32321),
            .I(data_idxvec_5));
    Odrv4 I__5899 (
            .O(N__32318),
            .I(data_idxvec_5));
    CascadeMux I__5898 (
            .O(N__32313),
            .I(n26_adj_1630_cascade_));
    CascadeMux I__5897 (
            .O(N__32310),
            .I(n22449_cascade_));
    InMux I__5896 (
            .O(N__32307),
            .I(N__32302));
    CascadeMux I__5895 (
            .O(N__32306),
            .I(N__32299));
    InMux I__5894 (
            .O(N__32305),
            .I(N__32296));
    LocalMux I__5893 (
            .O(N__32302),
            .I(N__32293));
    InMux I__5892 (
            .O(N__32299),
            .I(N__32290));
    LocalMux I__5891 (
            .O(N__32296),
            .I(req_data_cnt_5));
    Odrv4 I__5890 (
            .O(N__32293),
            .I(req_data_cnt_5));
    LocalMux I__5889 (
            .O(N__32290),
            .I(req_data_cnt_5));
    InMux I__5888 (
            .O(N__32283),
            .I(N__32280));
    LocalMux I__5887 (
            .O(N__32280),
            .I(n22368));
    CascadeMux I__5886 (
            .O(N__32277),
            .I(n22452_cascade_));
    InMux I__5885 (
            .O(N__32274),
            .I(N__32271));
    LocalMux I__5884 (
            .O(N__32271),
            .I(N__32267));
    InMux I__5883 (
            .O(N__32270),
            .I(N__32264));
    Span4Mux_h I__5882 (
            .O(N__32267),
            .I(N__32261));
    LocalMux I__5881 (
            .O(N__32264),
            .I(n14_adj_1551));
    Odrv4 I__5880 (
            .O(N__32261),
            .I(n14_adj_1551));
    InMux I__5879 (
            .O(N__32256),
            .I(N__32252));
    InMux I__5878 (
            .O(N__32255),
            .I(N__32249));
    LocalMux I__5877 (
            .O(N__32252),
            .I(N__32246));
    LocalMux I__5876 (
            .O(N__32249),
            .I(N__32242));
    Span12Mux_v I__5875 (
            .O(N__32246),
            .I(N__32239));
    InMux I__5874 (
            .O(N__32245),
            .I(N__32236));
    Span4Mux_v I__5873 (
            .O(N__32242),
            .I(N__32233));
    Odrv12 I__5872 (
            .O(N__32239),
            .I(buf_dds0_4));
    LocalMux I__5871 (
            .O(N__32236),
            .I(buf_dds0_4));
    Odrv4 I__5870 (
            .O(N__32233),
            .I(buf_dds0_4));
    CascadeMux I__5869 (
            .O(N__32226),
            .I(N__32223));
    InMux I__5868 (
            .O(N__32223),
            .I(N__32220));
    LocalMux I__5867 (
            .O(N__32220),
            .I(n23_adj_1661));
    InMux I__5866 (
            .O(N__32217),
            .I(N__32212));
    InMux I__5865 (
            .O(N__32216),
            .I(N__32207));
    InMux I__5864 (
            .O(N__32215),
            .I(N__32207));
    LocalMux I__5863 (
            .O(N__32212),
            .I(acadc_skipCount_14));
    LocalMux I__5862 (
            .O(N__32207),
            .I(acadc_skipCount_14));
    InMux I__5861 (
            .O(N__32202),
            .I(N__32199));
    LocalMux I__5860 (
            .O(N__32199),
            .I(N__32196));
    Span4Mux_v I__5859 (
            .O(N__32196),
            .I(N__32192));
    InMux I__5858 (
            .O(N__32195),
            .I(N__32189));
    Odrv4 I__5857 (
            .O(N__32192),
            .I(buf_adcdata_vdc_1));
    LocalMux I__5856 (
            .O(N__32189),
            .I(buf_adcdata_vdc_1));
    InMux I__5855 (
            .O(N__32184),
            .I(N__32181));
    LocalMux I__5854 (
            .O(N__32181),
            .I(N__32178));
    Span4Mux_h I__5853 (
            .O(N__32178),
            .I(N__32175));
    Span4Mux_v I__5852 (
            .O(N__32175),
            .I(N__32171));
    InMux I__5851 (
            .O(N__32174),
            .I(N__32168));
    Span4Mux_h I__5850 (
            .O(N__32171),
            .I(N__32163));
    LocalMux I__5849 (
            .O(N__32168),
            .I(N__32163));
    Span4Mux_h I__5848 (
            .O(N__32163),
            .I(N__32159));
    InMux I__5847 (
            .O(N__32162),
            .I(N__32156));
    Span4Mux_h I__5846 (
            .O(N__32159),
            .I(N__32153));
    LocalMux I__5845 (
            .O(N__32156),
            .I(buf_adcdata_vac_1));
    Odrv4 I__5844 (
            .O(N__32153),
            .I(buf_adcdata_vac_1));
    InMux I__5843 (
            .O(N__32148),
            .I(N__32145));
    LocalMux I__5842 (
            .O(N__32145),
            .I(N__32142));
    Span4Mux_v I__5841 (
            .O(N__32142),
            .I(N__32138));
    InMux I__5840 (
            .O(N__32141),
            .I(N__32135));
    Sp12to4 I__5839 (
            .O(N__32138),
            .I(N__32132));
    LocalMux I__5838 (
            .O(N__32135),
            .I(N__32129));
    Span12Mux_h I__5837 (
            .O(N__32132),
            .I(N__32125));
    Span4Mux_v I__5836 (
            .O(N__32129),
            .I(N__32122));
    InMux I__5835 (
            .O(N__32128),
            .I(N__32119));
    Span12Mux_v I__5834 (
            .O(N__32125),
            .I(N__32116));
    Span4Mux_v I__5833 (
            .O(N__32122),
            .I(N__32113));
    LocalMux I__5832 (
            .O(N__32119),
            .I(buf_adcdata_iac_20));
    Odrv12 I__5831 (
            .O(N__32116),
            .I(buf_adcdata_iac_20));
    Odrv4 I__5830 (
            .O(N__32113),
            .I(buf_adcdata_iac_20));
    IoInMux I__5829 (
            .O(N__32106),
            .I(N__32103));
    LocalMux I__5828 (
            .O(N__32103),
            .I(N__32100));
    Span4Mux_s1_h I__5827 (
            .O(N__32100),
            .I(N__32097));
    Sp12to4 I__5826 (
            .O(N__32097),
            .I(N__32094));
    Span12Mux_v I__5825 (
            .O(N__32094),
            .I(N__32091));
    Span12Mux_h I__5824 (
            .O(N__32091),
            .I(N__32086));
    InMux I__5823 (
            .O(N__32090),
            .I(N__32083));
    InMux I__5822 (
            .O(N__32089),
            .I(N__32080));
    Odrv12 I__5821 (
            .O(N__32086),
            .I(VAC_OSR0));
    LocalMux I__5820 (
            .O(N__32083),
            .I(VAC_OSR0));
    LocalMux I__5819 (
            .O(N__32080),
            .I(VAC_OSR0));
    CascadeMux I__5818 (
            .O(N__32073),
            .I(N__32070));
    InMux I__5817 (
            .O(N__32070),
            .I(N__32066));
    InMux I__5816 (
            .O(N__32069),
            .I(N__32063));
    LocalMux I__5815 (
            .O(N__32066),
            .I(N__32060));
    LocalMux I__5814 (
            .O(N__32063),
            .I(N__32057));
    Span4Mux_v I__5813 (
            .O(N__32060),
            .I(N__32054));
    Span4Mux_v I__5812 (
            .O(N__32057),
            .I(N__32049));
    Span4Mux_h I__5811 (
            .O(N__32054),
            .I(N__32049));
    Odrv4 I__5810 (
            .O(N__32049),
            .I(n30));
    InMux I__5809 (
            .O(N__32046),
            .I(N__32043));
    LocalMux I__5808 (
            .O(N__32043),
            .I(N__32039));
    InMux I__5807 (
            .O(N__32042),
            .I(N__32036));
    Span4Mux_v I__5806 (
            .O(N__32039),
            .I(N__32033));
    LocalMux I__5805 (
            .O(N__32036),
            .I(N__32030));
    Span4Mux_h I__5804 (
            .O(N__32033),
            .I(N__32025));
    Span4Mux_v I__5803 (
            .O(N__32030),
            .I(N__32025));
    Span4Mux_v I__5802 (
            .O(N__32025),
            .I(N__32022));
    Odrv4 I__5801 (
            .O(N__32022),
            .I(n14_adj_1574));
    InMux I__5800 (
            .O(N__32019),
            .I(N__32016));
    LocalMux I__5799 (
            .O(N__32016),
            .I(N__32013));
    Span4Mux_h I__5798 (
            .O(N__32013),
            .I(N__32010));
    Span4Mux_h I__5797 (
            .O(N__32010),
            .I(N__32007));
    Span4Mux_v I__5796 (
            .O(N__32007),
            .I(N__32004));
    Odrv4 I__5795 (
            .O(N__32004),
            .I(buf_data_iac_3));
    InMux I__5794 (
            .O(N__32001),
            .I(N__31998));
    LocalMux I__5793 (
            .O(N__31998),
            .I(N__31995));
    Odrv12 I__5792 (
            .O(N__31995),
            .I(n22_adj_1610));
    CascadeMux I__5791 (
            .O(N__31992),
            .I(N__31987));
    InMux I__5790 (
            .O(N__31991),
            .I(N__31982));
    InMux I__5789 (
            .O(N__31990),
            .I(N__31982));
    InMux I__5788 (
            .O(N__31987),
            .I(N__31979));
    LocalMux I__5787 (
            .O(N__31982),
            .I(req_data_cnt_14));
    LocalMux I__5786 (
            .O(N__31979),
            .I(req_data_cnt_14));
    InMux I__5785 (
            .O(N__31974),
            .I(N__31971));
    LocalMux I__5784 (
            .O(N__31971),
            .I(N__31968));
    Span12Mux_v I__5783 (
            .O(N__31968),
            .I(N__31963));
    InMux I__5782 (
            .O(N__31967),
            .I(N__31958));
    InMux I__5781 (
            .O(N__31966),
            .I(N__31958));
    Odrv12 I__5780 (
            .O(N__31963),
            .I(req_data_cnt_11));
    LocalMux I__5779 (
            .O(N__31958),
            .I(req_data_cnt_11));
    InMux I__5778 (
            .O(N__31953),
            .I(N__31950));
    LocalMux I__5777 (
            .O(N__31950),
            .I(n23));
    InMux I__5776 (
            .O(N__31947),
            .I(N__31944));
    LocalMux I__5775 (
            .O(N__31944),
            .I(\ADC_VDC.n21211 ));
    CEMux I__5774 (
            .O(N__31941),
            .I(N__31938));
    LocalMux I__5773 (
            .O(N__31938),
            .I(N__31935));
    Odrv4 I__5772 (
            .O(N__31935),
            .I(\ADC_VDC.n13368 ));
    InMux I__5771 (
            .O(N__31932),
            .I(N__31929));
    LocalMux I__5770 (
            .O(N__31929),
            .I(N__31925));
    InMux I__5769 (
            .O(N__31928),
            .I(N__31922));
    Span4Mux_h I__5768 (
            .O(N__31925),
            .I(N__31919));
    LocalMux I__5767 (
            .O(N__31922),
            .I(secclk_cnt_20));
    Odrv4 I__5766 (
            .O(N__31919),
            .I(secclk_cnt_20));
    CascadeMux I__5765 (
            .O(N__31914),
            .I(n20048_cascade_));
    InMux I__5764 (
            .O(N__31911),
            .I(N__31908));
    LocalMux I__5763 (
            .O(N__31908),
            .I(N__31905));
    Odrv4 I__5762 (
            .O(N__31905),
            .I(n14));
    InMux I__5761 (
            .O(N__31902),
            .I(N__31899));
    LocalMux I__5760 (
            .O(N__31899),
            .I(N__31896));
    Span4Mux_h I__5759 (
            .O(N__31896),
            .I(N__31892));
    InMux I__5758 (
            .O(N__31895),
            .I(N__31889));
    Odrv4 I__5757 (
            .O(N__31892),
            .I(buf_adcdata_vdc_20));
    LocalMux I__5756 (
            .O(N__31889),
            .I(buf_adcdata_vdc_20));
    InMux I__5755 (
            .O(N__31884),
            .I(N__31881));
    LocalMux I__5754 (
            .O(N__31881),
            .I(N__31878));
    Span4Mux_h I__5753 (
            .O(N__31878),
            .I(N__31875));
    Span4Mux_v I__5752 (
            .O(N__31875),
            .I(N__31872));
    Span4Mux_h I__5751 (
            .O(N__31872),
            .I(N__31868));
    InMux I__5750 (
            .O(N__31871),
            .I(N__31865));
    Span4Mux_h I__5749 (
            .O(N__31868),
            .I(N__31860));
    LocalMux I__5748 (
            .O(N__31865),
            .I(N__31860));
    Span4Mux_h I__5747 (
            .O(N__31860),
            .I(N__31856));
    InMux I__5746 (
            .O(N__31859),
            .I(N__31853));
    Span4Mux_v I__5745 (
            .O(N__31856),
            .I(N__31850));
    LocalMux I__5744 (
            .O(N__31853),
            .I(buf_adcdata_vac_20));
    Odrv4 I__5743 (
            .O(N__31850),
            .I(buf_adcdata_vac_20));
    InMux I__5742 (
            .O(N__31845),
            .I(N__31841));
    InMux I__5741 (
            .O(N__31844),
            .I(N__31838));
    LocalMux I__5740 (
            .O(N__31841),
            .I(secclk_cnt_6));
    LocalMux I__5739 (
            .O(N__31838),
            .I(secclk_cnt_6));
    InMux I__5738 (
            .O(N__31833),
            .I(N__31829));
    InMux I__5737 (
            .O(N__31832),
            .I(N__31826));
    LocalMux I__5736 (
            .O(N__31829),
            .I(secclk_cnt_14));
    LocalMux I__5735 (
            .O(N__31826),
            .I(secclk_cnt_14));
    CascadeMux I__5734 (
            .O(N__31821),
            .I(N__31818));
    InMux I__5733 (
            .O(N__31818),
            .I(N__31814));
    InMux I__5732 (
            .O(N__31817),
            .I(N__31811));
    LocalMux I__5731 (
            .O(N__31814),
            .I(N__31808));
    LocalMux I__5730 (
            .O(N__31811),
            .I(secclk_cnt_10));
    Odrv4 I__5729 (
            .O(N__31808),
            .I(secclk_cnt_10));
    InMux I__5728 (
            .O(N__31803),
            .I(N__31799));
    InMux I__5727 (
            .O(N__31802),
            .I(N__31796));
    LocalMux I__5726 (
            .O(N__31799),
            .I(secclk_cnt_3));
    LocalMux I__5725 (
            .O(N__31796),
            .I(secclk_cnt_3));
    InMux I__5724 (
            .O(N__31791),
            .I(N__31788));
    LocalMux I__5723 (
            .O(N__31788),
            .I(n27));
    InMux I__5722 (
            .O(N__31785),
            .I(N__31781));
    InMux I__5721 (
            .O(N__31784),
            .I(N__31778));
    LocalMux I__5720 (
            .O(N__31781),
            .I(secclk_cnt_2));
    LocalMux I__5719 (
            .O(N__31778),
            .I(secclk_cnt_2));
    InMux I__5718 (
            .O(N__31773),
            .I(N__31769));
    InMux I__5717 (
            .O(N__31772),
            .I(N__31766));
    LocalMux I__5716 (
            .O(N__31769),
            .I(secclk_cnt_13));
    LocalMux I__5715 (
            .O(N__31766),
            .I(secclk_cnt_13));
    CascadeMux I__5714 (
            .O(N__31761),
            .I(N__31757));
    InMux I__5713 (
            .O(N__31760),
            .I(N__31754));
    InMux I__5712 (
            .O(N__31757),
            .I(N__31751));
    LocalMux I__5711 (
            .O(N__31754),
            .I(secclk_cnt_7));
    LocalMux I__5710 (
            .O(N__31751),
            .I(secclk_cnt_7));
    InMux I__5709 (
            .O(N__31746),
            .I(N__31742));
    InMux I__5708 (
            .O(N__31745),
            .I(N__31739));
    LocalMux I__5707 (
            .O(N__31742),
            .I(secclk_cnt_16));
    LocalMux I__5706 (
            .O(N__31739),
            .I(secclk_cnt_16));
    InMux I__5705 (
            .O(N__31734),
            .I(N__31731));
    LocalMux I__5704 (
            .O(N__31731),
            .I(n26_adj_1656));
    InMux I__5703 (
            .O(N__31728),
            .I(N__31724));
    InMux I__5702 (
            .O(N__31727),
            .I(N__31721));
    LocalMux I__5701 (
            .O(N__31724),
            .I(N__31718));
    LocalMux I__5700 (
            .O(N__31721),
            .I(N__31715));
    Span4Mux_v I__5699 (
            .O(N__31718),
            .I(N__31710));
    Span4Mux_h I__5698 (
            .O(N__31715),
            .I(N__31710));
    Odrv4 I__5697 (
            .O(N__31710),
            .I(n14_adj_1552));
    InMux I__5696 (
            .O(N__31707),
            .I(N__31704));
    LocalMux I__5695 (
            .O(N__31704),
            .I(\ADC_VDC.n11 ));
    InMux I__5694 (
            .O(N__31701),
            .I(N__31698));
    LocalMux I__5693 (
            .O(N__31698),
            .I(\ADC_VDC.n65 ));
    CascadeMux I__5692 (
            .O(N__31695),
            .I(N__31692));
    InMux I__5691 (
            .O(N__31692),
            .I(N__31689));
    LocalMux I__5690 (
            .O(N__31689),
            .I(\ADC_VDC.n21133 ));
    CEMux I__5689 (
            .O(N__31686),
            .I(N__31683));
    LocalMux I__5688 (
            .O(N__31683),
            .I(\ADC_VDC.n42_adj_1452 ));
    InMux I__5687 (
            .O(N__31680),
            .I(N__31677));
    LocalMux I__5686 (
            .O(N__31677),
            .I(N__31674));
    Odrv4 I__5685 (
            .O(N__31674),
            .I(\ADC_VDC.n20998 ));
    InMux I__5684 (
            .O(N__31671),
            .I(N__31668));
    LocalMux I__5683 (
            .O(N__31668),
            .I(\ADC_VDC.n11494 ));
    CascadeMux I__5682 (
            .O(N__31665),
            .I(\ADC_VDC.n11494_cascade_ ));
    CascadeMux I__5681 (
            .O(N__31662),
            .I(N__31658));
    InMux I__5680 (
            .O(N__31661),
            .I(N__31655));
    InMux I__5679 (
            .O(N__31658),
            .I(N__31652));
    LocalMux I__5678 (
            .O(N__31655),
            .I(N__31649));
    LocalMux I__5677 (
            .O(N__31652),
            .I(N__31646));
    Span4Mux_h I__5676 (
            .O(N__31649),
            .I(N__31643));
    Span4Mux_v I__5675 (
            .O(N__31646),
            .I(N__31640));
    Odrv4 I__5674 (
            .O(N__31643),
            .I(\ADC_VDC.n15 ));
    Odrv4 I__5673 (
            .O(N__31640),
            .I(\ADC_VDC.n15 ));
    CascadeMux I__5672 (
            .O(N__31635),
            .I(\ADC_VDC.n15_cascade_ ));
    InMux I__5671 (
            .O(N__31632),
            .I(N__31629));
    LocalMux I__5670 (
            .O(N__31629),
            .I(\ADC_VDC.n21185 ));
    InMux I__5669 (
            .O(N__31626),
            .I(N__31621));
    InMux I__5668 (
            .O(N__31625),
            .I(N__31614));
    CascadeMux I__5667 (
            .O(N__31624),
            .I(N__31611));
    LocalMux I__5666 (
            .O(N__31621),
            .I(N__31605));
    InMux I__5665 (
            .O(N__31620),
            .I(N__31602));
    CascadeMux I__5664 (
            .O(N__31619),
            .I(N__31597));
    CascadeMux I__5663 (
            .O(N__31618),
            .I(N__31594));
    CascadeMux I__5662 (
            .O(N__31617),
            .I(N__31591));
    LocalMux I__5661 (
            .O(N__31614),
            .I(N__31577));
    InMux I__5660 (
            .O(N__31611),
            .I(N__31570));
    InMux I__5659 (
            .O(N__31610),
            .I(N__31570));
    InMux I__5658 (
            .O(N__31609),
            .I(N__31570));
    InMux I__5657 (
            .O(N__31608),
            .I(N__31567));
    Span4Mux_v I__5656 (
            .O(N__31605),
            .I(N__31562));
    LocalMux I__5655 (
            .O(N__31602),
            .I(N__31562));
    InMux I__5654 (
            .O(N__31601),
            .I(N__31549));
    InMux I__5653 (
            .O(N__31600),
            .I(N__31549));
    InMux I__5652 (
            .O(N__31597),
            .I(N__31549));
    InMux I__5651 (
            .O(N__31594),
            .I(N__31549));
    InMux I__5650 (
            .O(N__31591),
            .I(N__31549));
    InMux I__5649 (
            .O(N__31590),
            .I(N__31549));
    InMux I__5648 (
            .O(N__31589),
            .I(N__31540));
    InMux I__5647 (
            .O(N__31588),
            .I(N__31540));
    InMux I__5646 (
            .O(N__31587),
            .I(N__31540));
    InMux I__5645 (
            .O(N__31586),
            .I(N__31540));
    InMux I__5644 (
            .O(N__31585),
            .I(N__31537));
    InMux I__5643 (
            .O(N__31584),
            .I(N__31526));
    InMux I__5642 (
            .O(N__31583),
            .I(N__31526));
    InMux I__5641 (
            .O(N__31582),
            .I(N__31526));
    InMux I__5640 (
            .O(N__31581),
            .I(N__31526));
    InMux I__5639 (
            .O(N__31580),
            .I(N__31526));
    Span4Mux_v I__5638 (
            .O(N__31577),
            .I(N__31521));
    LocalMux I__5637 (
            .O(N__31570),
            .I(N__31521));
    LocalMux I__5636 (
            .O(N__31567),
            .I(N__31518));
    Span4Mux_h I__5635 (
            .O(N__31562),
            .I(N__31513));
    LocalMux I__5634 (
            .O(N__31549),
            .I(N__31513));
    LocalMux I__5633 (
            .O(N__31540),
            .I(N__31502));
    LocalMux I__5632 (
            .O(N__31537),
            .I(N__31502));
    LocalMux I__5631 (
            .O(N__31526),
            .I(N__31502));
    Span4Mux_v I__5630 (
            .O(N__31521),
            .I(N__31502));
    Span4Mux_v I__5629 (
            .O(N__31518),
            .I(N__31502));
    Odrv4 I__5628 (
            .O(N__31513),
            .I(n11891));
    Odrv4 I__5627 (
            .O(N__31502),
            .I(n11891));
    CascadeMux I__5626 (
            .O(N__31497),
            .I(N__31494));
    InMux I__5625 (
            .O(N__31494),
            .I(N__31490));
    CascadeMux I__5624 (
            .O(N__31493),
            .I(N__31487));
    LocalMux I__5623 (
            .O(N__31490),
            .I(N__31484));
    InMux I__5622 (
            .O(N__31487),
            .I(N__31481));
    Span4Mux_v I__5621 (
            .O(N__31484),
            .I(N__31478));
    LocalMux I__5620 (
            .O(N__31481),
            .I(N__31475));
    Odrv4 I__5619 (
            .O(N__31478),
            .I(cmd_rdadcbuf_12));
    Odrv4 I__5618 (
            .O(N__31475),
            .I(cmd_rdadcbuf_12));
    InMux I__5617 (
            .O(N__31470),
            .I(N__31467));
    LocalMux I__5616 (
            .O(N__31467),
            .I(\ADC_VDC.n21203 ));
    CascadeMux I__5615 (
            .O(N__31464),
            .I(N__31461));
    InMux I__5614 (
            .O(N__31461),
            .I(N__31458));
    LocalMux I__5613 (
            .O(N__31458),
            .I(\SIG_DDS.tmp_buf_1 ));
    InMux I__5612 (
            .O(N__31455),
            .I(N__31452));
    LocalMux I__5611 (
            .O(N__31452),
            .I(N__31449));
    Span4Mux_v I__5610 (
            .O(N__31449),
            .I(N__31444));
    InMux I__5609 (
            .O(N__31448),
            .I(N__31439));
    InMux I__5608 (
            .O(N__31447),
            .I(N__31439));
    Odrv4 I__5607 (
            .O(N__31444),
            .I(buf_dds0_2));
    LocalMux I__5606 (
            .O(N__31439),
            .I(buf_dds0_2));
    CascadeMux I__5605 (
            .O(N__31434),
            .I(N__31431));
    InMux I__5604 (
            .O(N__31431),
            .I(N__31428));
    LocalMux I__5603 (
            .O(N__31428),
            .I(\SIG_DDS.tmp_buf_2 ));
    CascadeMux I__5602 (
            .O(N__31425),
            .I(N__31422));
    InMux I__5601 (
            .O(N__31422),
            .I(N__31419));
    LocalMux I__5600 (
            .O(N__31419),
            .I(\SIG_DDS.tmp_buf_3 ));
    CascadeMux I__5599 (
            .O(N__31416),
            .I(N__31413));
    InMux I__5598 (
            .O(N__31413),
            .I(N__31410));
    LocalMux I__5597 (
            .O(N__31410),
            .I(\SIG_DDS.tmp_buf_4 ));
    CascadeMux I__5596 (
            .O(N__31407),
            .I(N__31404));
    InMux I__5595 (
            .O(N__31404),
            .I(N__31401));
    LocalMux I__5594 (
            .O(N__31401),
            .I(\SIG_DDS.tmp_buf_5 ));
    CascadeMux I__5593 (
            .O(N__31398),
            .I(N__31395));
    InMux I__5592 (
            .O(N__31395),
            .I(N__31392));
    LocalMux I__5591 (
            .O(N__31392),
            .I(N__31389));
    Odrv4 I__5590 (
            .O(N__31389),
            .I(\ADC_VDC.n21007 ));
    CascadeMux I__5589 (
            .O(N__31386),
            .I(\ADC_VDC.n21007_cascade_ ));
    SRMux I__5588 (
            .O(N__31383),
            .I(N__31380));
    LocalMux I__5587 (
            .O(N__31380),
            .I(\ADC_VDC.n4 ));
    CascadeMux I__5586 (
            .O(N__31377),
            .I(N__31374));
    InMux I__5585 (
            .O(N__31374),
            .I(N__31371));
    LocalMux I__5584 (
            .O(N__31371),
            .I(\SIG_DDS.tmp_buf_10 ));
    InMux I__5583 (
            .O(N__31368),
            .I(N__31363));
    InMux I__5582 (
            .O(N__31367),
            .I(N__31360));
    InMux I__5581 (
            .O(N__31366),
            .I(N__31357));
    LocalMux I__5580 (
            .O(N__31363),
            .I(buf_dds0_11));
    LocalMux I__5579 (
            .O(N__31360),
            .I(buf_dds0_11));
    LocalMux I__5578 (
            .O(N__31357),
            .I(buf_dds0_11));
    CascadeMux I__5577 (
            .O(N__31350),
            .I(N__31347));
    InMux I__5576 (
            .O(N__31347),
            .I(N__31344));
    LocalMux I__5575 (
            .O(N__31344),
            .I(\SIG_DDS.tmp_buf_11 ));
    CascadeMux I__5574 (
            .O(N__31341),
            .I(N__31338));
    InMux I__5573 (
            .O(N__31338),
            .I(N__31335));
    LocalMux I__5572 (
            .O(N__31335),
            .I(\SIG_DDS.tmp_buf_12 ));
    CascadeMux I__5571 (
            .O(N__31332),
            .I(N__31329));
    InMux I__5570 (
            .O(N__31329),
            .I(N__31326));
    LocalMux I__5569 (
            .O(N__31326),
            .I(\SIG_DDS.tmp_buf_13 ));
    InMux I__5568 (
            .O(N__31323),
            .I(N__31320));
    LocalMux I__5567 (
            .O(N__31320),
            .I(N__31315));
    InMux I__5566 (
            .O(N__31319),
            .I(N__31312));
    InMux I__5565 (
            .O(N__31318),
            .I(N__31309));
    Span4Mux_v I__5564 (
            .O(N__31315),
            .I(N__31306));
    LocalMux I__5563 (
            .O(N__31312),
            .I(buf_dds0_14));
    LocalMux I__5562 (
            .O(N__31309),
            .I(buf_dds0_14));
    Odrv4 I__5561 (
            .O(N__31306),
            .I(buf_dds0_14));
    CascadeMux I__5560 (
            .O(N__31299),
            .I(N__31295));
    CascadeMux I__5559 (
            .O(N__31298),
            .I(N__31291));
    InMux I__5558 (
            .O(N__31295),
            .I(N__31288));
    CascadeMux I__5557 (
            .O(N__31294),
            .I(N__31285));
    InMux I__5556 (
            .O(N__31291),
            .I(N__31282));
    LocalMux I__5555 (
            .O(N__31288),
            .I(N__31279));
    InMux I__5554 (
            .O(N__31285),
            .I(N__31276));
    LocalMux I__5553 (
            .O(N__31282),
            .I(N__31273));
    Span4Mux_h I__5552 (
            .O(N__31279),
            .I(N__31270));
    LocalMux I__5551 (
            .O(N__31276),
            .I(buf_dds0_15));
    Odrv12 I__5550 (
            .O(N__31273),
            .I(buf_dds0_15));
    Odrv4 I__5549 (
            .O(N__31270),
            .I(buf_dds0_15));
    InMux I__5548 (
            .O(N__31263),
            .I(N__31260));
    LocalMux I__5547 (
            .O(N__31260),
            .I(\SIG_DDS.tmp_buf_14 ));
    InMux I__5546 (
            .O(N__31257),
            .I(N__31254));
    LocalMux I__5545 (
            .O(N__31254),
            .I(N__31249));
    InMux I__5544 (
            .O(N__31253),
            .I(N__31246));
    InMux I__5543 (
            .O(N__31252),
            .I(N__31243));
    Span4Mux_v I__5542 (
            .O(N__31249),
            .I(N__31238));
    LocalMux I__5541 (
            .O(N__31246),
            .I(N__31238));
    LocalMux I__5540 (
            .O(N__31243),
            .I(buf_dds0_9));
    Odrv4 I__5539 (
            .O(N__31238),
            .I(buf_dds0_9));
    CascadeMux I__5538 (
            .O(N__31233),
            .I(N__31230));
    InMux I__5537 (
            .O(N__31230),
            .I(N__31227));
    LocalMux I__5536 (
            .O(N__31227),
            .I(\SIG_DDS.tmp_buf_9 ));
    CascadeMux I__5535 (
            .O(N__31224),
            .I(N__31221));
    InMux I__5534 (
            .O(N__31221),
            .I(N__31218));
    LocalMux I__5533 (
            .O(N__31218),
            .I(N__31215));
    Odrv4 I__5532 (
            .O(N__31215),
            .I(\SIG_DDS.tmp_buf_8 ));
    CascadeMux I__5531 (
            .O(N__31212),
            .I(N__31209));
    InMux I__5530 (
            .O(N__31209),
            .I(N__31206));
    LocalMux I__5529 (
            .O(N__31206),
            .I(\SIG_DDS.tmp_buf_0 ));
    InMux I__5528 (
            .O(N__31203),
            .I(N__31200));
    LocalMux I__5527 (
            .O(N__31200),
            .I(N__31195));
    InMux I__5526 (
            .O(N__31199),
            .I(N__31190));
    InMux I__5525 (
            .O(N__31198),
            .I(N__31190));
    Odrv4 I__5524 (
            .O(N__31195),
            .I(buf_dds0_1));
    LocalMux I__5523 (
            .O(N__31190),
            .I(buf_dds0_1));
    CascadeMux I__5522 (
            .O(N__31185),
            .I(N__31181));
    InMux I__5521 (
            .O(N__31184),
            .I(N__31178));
    InMux I__5520 (
            .O(N__31181),
            .I(N__31175));
    LocalMux I__5519 (
            .O(N__31178),
            .I(N__31172));
    LocalMux I__5518 (
            .O(N__31175),
            .I(N__31166));
    Sp12to4 I__5517 (
            .O(N__31172),
            .I(N__31166));
    InMux I__5516 (
            .O(N__31171),
            .I(N__31163));
    Odrv12 I__5515 (
            .O(N__31166),
            .I(acadc_skipCount_15));
    LocalMux I__5514 (
            .O(N__31163),
            .I(acadc_skipCount_15));
    CascadeMux I__5513 (
            .O(N__31158),
            .I(N__31155));
    InMux I__5512 (
            .O(N__31155),
            .I(N__31151));
    InMux I__5511 (
            .O(N__31154),
            .I(N__31148));
    LocalMux I__5510 (
            .O(N__31151),
            .I(N__31145));
    LocalMux I__5509 (
            .O(N__31148),
            .I(n11570));
    Odrv12 I__5508 (
            .O(N__31145),
            .I(n11570));
    InMux I__5507 (
            .O(N__31140),
            .I(N__31137));
    LocalMux I__5506 (
            .O(N__31137),
            .I(N__31134));
    Sp12to4 I__5505 (
            .O(N__31134),
            .I(N__31131));
    Span12Mux_v I__5504 (
            .O(N__31131),
            .I(N__31128));
    Odrv12 I__5503 (
            .O(N__31128),
            .I(EIS_SYNCCLK));
    IoInMux I__5502 (
            .O(N__31125),
            .I(N__31122));
    LocalMux I__5501 (
            .O(N__31122),
            .I(N__31118));
    IoInMux I__5500 (
            .O(N__31121),
            .I(N__31115));
    Span4Mux_s2_v I__5499 (
            .O(N__31118),
            .I(N__31112));
    LocalMux I__5498 (
            .O(N__31115),
            .I(N__31109));
    Span4Mux_v I__5497 (
            .O(N__31112),
            .I(N__31106));
    IoSpan4Mux I__5496 (
            .O(N__31109),
            .I(N__31103));
    Span4Mux_v I__5495 (
            .O(N__31106),
            .I(N__31098));
    Span4Mux_s3_h I__5494 (
            .O(N__31103),
            .I(N__31098));
    Sp12to4 I__5493 (
            .O(N__31098),
            .I(N__31095));
    Odrv12 I__5492 (
            .O(N__31095),
            .I(IAC_CLK));
    InMux I__5491 (
            .O(N__31092),
            .I(N__31088));
    InMux I__5490 (
            .O(N__31091),
            .I(N__31085));
    LocalMux I__5489 (
            .O(N__31088),
            .I(N__31082));
    LocalMux I__5488 (
            .O(N__31085),
            .I(N__31078));
    Span4Mux_h I__5487 (
            .O(N__31082),
            .I(N__31075));
    InMux I__5486 (
            .O(N__31081),
            .I(N__31072));
    Span4Mux_h I__5485 (
            .O(N__31078),
            .I(N__31069));
    Odrv4 I__5484 (
            .O(N__31075),
            .I(buf_dds0_10));
    LocalMux I__5483 (
            .O(N__31072),
            .I(buf_dds0_10));
    Odrv4 I__5482 (
            .O(N__31069),
            .I(buf_dds0_10));
    CascadeMux I__5481 (
            .O(N__31062),
            .I(n21501_cascade_));
    InMux I__5480 (
            .O(N__31059),
            .I(N__31056));
    LocalMux I__5479 (
            .O(N__31056),
            .I(eis_state_2_N_392_0));
    InMux I__5478 (
            .O(N__31053),
            .I(N__31050));
    LocalMux I__5477 (
            .O(N__31050),
            .I(n22479));
    InMux I__5476 (
            .O(N__31047),
            .I(N__31040));
    InMux I__5475 (
            .O(N__31046),
            .I(N__31040));
    CascadeMux I__5474 (
            .O(N__31045),
            .I(N__31037));
    LocalMux I__5473 (
            .O(N__31040),
            .I(N__31034));
    InMux I__5472 (
            .O(N__31037),
            .I(N__31031));
    Span4Mux_v I__5471 (
            .O(N__31034),
            .I(N__31025));
    LocalMux I__5470 (
            .O(N__31031),
            .I(N__31022));
    InMux I__5469 (
            .O(N__31030),
            .I(N__31017));
    InMux I__5468 (
            .O(N__31029),
            .I(N__31017));
    InMux I__5467 (
            .O(N__31028),
            .I(N__31014));
    Span4Mux_h I__5466 (
            .O(N__31025),
            .I(N__31011));
    Span4Mux_h I__5465 (
            .O(N__31022),
            .I(N__31006));
    LocalMux I__5464 (
            .O(N__31017),
            .I(N__31006));
    LocalMux I__5463 (
            .O(N__31014),
            .I(eis_start));
    Odrv4 I__5462 (
            .O(N__31011),
            .I(eis_start));
    Odrv4 I__5461 (
            .O(N__31006),
            .I(eis_start));
    CascadeMux I__5460 (
            .O(N__30999),
            .I(n11_adj_1632_cascade_));
    CEMux I__5459 (
            .O(N__30996),
            .I(N__30992));
    CEMux I__5458 (
            .O(N__30995),
            .I(N__30989));
    LocalMux I__5457 (
            .O(N__30992),
            .I(n11908));
    LocalMux I__5456 (
            .O(N__30989),
            .I(n11908));
    CascadeMux I__5455 (
            .O(N__30984),
            .I(N__30976));
    CascadeMux I__5454 (
            .O(N__30983),
            .I(N__30973));
    CascadeMux I__5453 (
            .O(N__30982),
            .I(N__30970));
    CascadeMux I__5452 (
            .O(N__30981),
            .I(N__30959));
    CascadeMux I__5451 (
            .O(N__30980),
            .I(N__30956));
    InMux I__5450 (
            .O(N__30979),
            .I(N__30944));
    InMux I__5449 (
            .O(N__30976),
            .I(N__30944));
    InMux I__5448 (
            .O(N__30973),
            .I(N__30944));
    InMux I__5447 (
            .O(N__30970),
            .I(N__30944));
    InMux I__5446 (
            .O(N__30969),
            .I(N__30944));
    InMux I__5445 (
            .O(N__30968),
            .I(N__30937));
    InMux I__5444 (
            .O(N__30967),
            .I(N__30937));
    InMux I__5443 (
            .O(N__30966),
            .I(N__30937));
    InMux I__5442 (
            .O(N__30965),
            .I(N__30932));
    InMux I__5441 (
            .O(N__30964),
            .I(N__30932));
    InMux I__5440 (
            .O(N__30963),
            .I(N__30929));
    InMux I__5439 (
            .O(N__30962),
            .I(N__30920));
    InMux I__5438 (
            .O(N__30959),
            .I(N__30920));
    InMux I__5437 (
            .O(N__30956),
            .I(N__30920));
    InMux I__5436 (
            .O(N__30955),
            .I(N__30920));
    LocalMux I__5435 (
            .O(N__30944),
            .I(eis_state_0));
    LocalMux I__5434 (
            .O(N__30937),
            .I(eis_state_0));
    LocalMux I__5433 (
            .O(N__30932),
            .I(eis_state_0));
    LocalMux I__5432 (
            .O(N__30929),
            .I(eis_state_0));
    LocalMux I__5431 (
            .O(N__30920),
            .I(eis_state_0));
    InMux I__5430 (
            .O(N__30909),
            .I(N__30905));
    InMux I__5429 (
            .O(N__30908),
            .I(N__30902));
    LocalMux I__5428 (
            .O(N__30905),
            .I(n21041));
    LocalMux I__5427 (
            .O(N__30902),
            .I(n21041));
    InMux I__5426 (
            .O(N__30897),
            .I(N__30894));
    LocalMux I__5425 (
            .O(N__30894),
            .I(N__30890));
    InMux I__5424 (
            .O(N__30893),
            .I(N__30886));
    Span4Mux_h I__5423 (
            .O(N__30890),
            .I(N__30883));
    InMux I__5422 (
            .O(N__30889),
            .I(N__30880));
    LocalMux I__5421 (
            .O(N__30886),
            .I(buf_dds1_15));
    Odrv4 I__5420 (
            .O(N__30883),
            .I(buf_dds1_15));
    LocalMux I__5419 (
            .O(N__30880),
            .I(buf_dds1_15));
    InMux I__5418 (
            .O(N__30873),
            .I(N__30869));
    InMux I__5417 (
            .O(N__30872),
            .I(N__30866));
    LocalMux I__5416 (
            .O(N__30869),
            .I(N__30863));
    LocalMux I__5415 (
            .O(N__30866),
            .I(N__30857));
    Span4Mux_h I__5414 (
            .O(N__30863),
            .I(N__30857));
    InMux I__5413 (
            .O(N__30862),
            .I(N__30854));
    Odrv4 I__5412 (
            .O(N__30857),
            .I(buf_dds1_10));
    LocalMux I__5411 (
            .O(N__30854),
            .I(buf_dds1_10));
    CascadeMux I__5410 (
            .O(N__30849),
            .I(n22395_cascade_));
    CascadeMux I__5409 (
            .O(N__30846),
            .I(N__30842));
    InMux I__5408 (
            .O(N__30845),
            .I(N__30838));
    InMux I__5407 (
            .O(N__30842),
            .I(N__30835));
    InMux I__5406 (
            .O(N__30841),
            .I(N__30832));
    LocalMux I__5405 (
            .O(N__30838),
            .I(N__30827));
    LocalMux I__5404 (
            .O(N__30835),
            .I(N__30827));
    LocalMux I__5403 (
            .O(N__30832),
            .I(req_data_cnt_8));
    Odrv4 I__5402 (
            .O(N__30827),
            .I(req_data_cnt_8));
    IoInMux I__5401 (
            .O(N__30822),
            .I(N__30819));
    LocalMux I__5400 (
            .O(N__30819),
            .I(N__30816));
    Span4Mux_s3_h I__5399 (
            .O(N__30816),
            .I(N__30813));
    Span4Mux_h I__5398 (
            .O(N__30813),
            .I(N__30810));
    Span4Mux_h I__5397 (
            .O(N__30810),
            .I(N__30807));
    Sp12to4 I__5396 (
            .O(N__30807),
            .I(N__30802));
    InMux I__5395 (
            .O(N__30806),
            .I(N__30799));
    InMux I__5394 (
            .O(N__30805),
            .I(N__30796));
    Span12Mux_v I__5393 (
            .O(N__30802),
            .I(N__30793));
    LocalMux I__5392 (
            .O(N__30799),
            .I(N__30790));
    LocalMux I__5391 (
            .O(N__30796),
            .I(N__30787));
    Odrv12 I__5390 (
            .O(N__30793),
            .I(VAC_FLT0));
    Odrv4 I__5389 (
            .O(N__30790),
            .I(VAC_FLT0));
    Odrv4 I__5388 (
            .O(N__30787),
            .I(VAC_FLT0));
    CascadeMux I__5387 (
            .O(N__30780),
            .I(N__30775));
    InMux I__5386 (
            .O(N__30779),
            .I(N__30772));
    CascadeMux I__5385 (
            .O(N__30778),
            .I(N__30769));
    InMux I__5384 (
            .O(N__30775),
            .I(N__30766));
    LocalMux I__5383 (
            .O(N__30772),
            .I(N__30763));
    InMux I__5382 (
            .O(N__30769),
            .I(N__30760));
    LocalMux I__5381 (
            .O(N__30766),
            .I(N__30757));
    Span4Mux_h I__5380 (
            .O(N__30763),
            .I(N__30754));
    LocalMux I__5379 (
            .O(N__30760),
            .I(N__30749));
    Span4Mux_v I__5378 (
            .O(N__30757),
            .I(N__30749));
    Sp12to4 I__5377 (
            .O(N__30754),
            .I(N__30746));
    Sp12to4 I__5376 (
            .O(N__30749),
            .I(N__30741));
    Span12Mux_v I__5375 (
            .O(N__30746),
            .I(N__30741));
    Odrv12 I__5374 (
            .O(N__30741),
            .I(buf_adcdata_iac_22));
    CascadeMux I__5373 (
            .O(N__30738),
            .I(n22635_cascade_));
    InMux I__5372 (
            .O(N__30735),
            .I(N__30732));
    LocalMux I__5371 (
            .O(N__30732),
            .I(N__30729));
    Span4Mux_h I__5370 (
            .O(N__30729),
            .I(N__30726));
    Odrv4 I__5369 (
            .O(N__30726),
            .I(n21236));
    InMux I__5368 (
            .O(N__30723),
            .I(N__30718));
    CascadeMux I__5367 (
            .O(N__30722),
            .I(N__30715));
    InMux I__5366 (
            .O(N__30721),
            .I(N__30712));
    LocalMux I__5365 (
            .O(N__30718),
            .I(N__30709));
    InMux I__5364 (
            .O(N__30715),
            .I(N__30706));
    LocalMux I__5363 (
            .O(N__30712),
            .I(N__30703));
    Span4Mux_v I__5362 (
            .O(N__30709),
            .I(N__30700));
    LocalMux I__5361 (
            .O(N__30706),
            .I(N__30697));
    Span4Mux_h I__5360 (
            .O(N__30703),
            .I(N__30694));
    Sp12to4 I__5359 (
            .O(N__30700),
            .I(N__30689));
    Span12Mux_v I__5358 (
            .O(N__30697),
            .I(N__30689));
    Span4Mux_h I__5357 (
            .O(N__30694),
            .I(N__30686));
    Odrv12 I__5356 (
            .O(N__30689),
            .I(n14_adj_1578));
    Odrv4 I__5355 (
            .O(N__30686),
            .I(n14_adj_1578));
    CascadeMux I__5354 (
            .O(N__30681),
            .I(n2_cascade_));
    InMux I__5353 (
            .O(N__30678),
            .I(N__30674));
    CascadeMux I__5352 (
            .O(N__30677),
            .I(N__30671));
    LocalMux I__5351 (
            .O(N__30674),
            .I(N__30668));
    InMux I__5350 (
            .O(N__30671),
            .I(N__30665));
    Span4Mux_v I__5349 (
            .O(N__30668),
            .I(N__30662));
    LocalMux I__5348 (
            .O(N__30665),
            .I(N__30657));
    Span4Mux_v I__5347 (
            .O(N__30662),
            .I(N__30657));
    Sp12to4 I__5346 (
            .O(N__30657),
            .I(N__30654));
    Odrv12 I__5345 (
            .O(N__30654),
            .I(data_idxvec_4));
    CascadeMux I__5344 (
            .O(N__30651),
            .I(n26_adj_1635_cascade_));
    CascadeMux I__5343 (
            .O(N__30648),
            .I(n22443_cascade_));
    CascadeMux I__5342 (
            .O(N__30645),
            .I(n22446_cascade_));
    CascadeMux I__5341 (
            .O(N__30642),
            .I(n30_adj_1636_cascade_));
    InMux I__5340 (
            .O(N__30639),
            .I(N__30636));
    LocalMux I__5339 (
            .O(N__30636),
            .I(n19_adj_1634));
    CascadeMux I__5338 (
            .O(N__30633),
            .I(N__30630));
    InMux I__5337 (
            .O(N__30630),
            .I(N__30627));
    LocalMux I__5336 (
            .O(N__30627),
            .I(N__30624));
    Span4Mux_v I__5335 (
            .O(N__30624),
            .I(N__30621));
    Span4Mux_h I__5334 (
            .O(N__30621),
            .I(N__30617));
    InMux I__5333 (
            .O(N__30620),
            .I(N__30614));
    Odrv4 I__5332 (
            .O(N__30617),
            .I(buf_readRTD_4));
    LocalMux I__5331 (
            .O(N__30614),
            .I(buf_readRTD_4));
    InMux I__5330 (
            .O(N__30609),
            .I(N__30605));
    InMux I__5329 (
            .O(N__30608),
            .I(N__30602));
    LocalMux I__5328 (
            .O(N__30605),
            .I(N__30598));
    LocalMux I__5327 (
            .O(N__30602),
            .I(N__30595));
    InMux I__5326 (
            .O(N__30601),
            .I(N__30592));
    Span12Mux_h I__5325 (
            .O(N__30598),
            .I(N__30589));
    Span4Mux_v I__5324 (
            .O(N__30595),
            .I(N__30586));
    LocalMux I__5323 (
            .O(N__30592),
            .I(buf_adcdata_iac_12));
    Odrv12 I__5322 (
            .O(N__30589),
            .I(buf_adcdata_iac_12));
    Odrv4 I__5321 (
            .O(N__30586),
            .I(buf_adcdata_iac_12));
    CascadeMux I__5320 (
            .O(N__30579),
            .I(n22467_cascade_));
    InMux I__5319 (
            .O(N__30576),
            .I(N__30573));
    LocalMux I__5318 (
            .O(N__30573),
            .I(N__30570));
    Span4Mux_v I__5317 (
            .O(N__30570),
            .I(N__30567));
    Odrv4 I__5316 (
            .O(N__30567),
            .I(n16_adj_1633));
    InMux I__5315 (
            .O(N__30564),
            .I(N__30561));
    LocalMux I__5314 (
            .O(N__30561),
            .I(n22470));
    InMux I__5313 (
            .O(N__30558),
            .I(N__30555));
    LocalMux I__5312 (
            .O(N__30555),
            .I(N__30552));
    Span4Mux_h I__5311 (
            .O(N__30552),
            .I(N__30549));
    Odrv4 I__5310 (
            .O(N__30549),
            .I(n21329));
    IoInMux I__5309 (
            .O(N__30546),
            .I(N__30543));
    LocalMux I__5308 (
            .O(N__30543),
            .I(N__30539));
    InMux I__5307 (
            .O(N__30542),
            .I(N__30536));
    IoSpan4Mux I__5306 (
            .O(N__30539),
            .I(N__30533));
    LocalMux I__5305 (
            .O(N__30536),
            .I(N__30530));
    Span4Mux_s2_v I__5304 (
            .O(N__30533),
            .I(N__30527));
    Span4Mux_h I__5303 (
            .O(N__30530),
            .I(N__30523));
    Span4Mux_v I__5302 (
            .O(N__30527),
            .I(N__30520));
    InMux I__5301 (
            .O(N__30526),
            .I(N__30517));
    Span4Mux_v I__5300 (
            .O(N__30523),
            .I(N__30514));
    Odrv4 I__5299 (
            .O(N__30520),
            .I(IAC_FLT0));
    LocalMux I__5298 (
            .O(N__30517),
            .I(IAC_FLT0));
    Odrv4 I__5297 (
            .O(N__30514),
            .I(IAC_FLT0));
    InMux I__5296 (
            .O(N__30507),
            .I(N__30504));
    LocalMux I__5295 (
            .O(N__30504),
            .I(N__30501));
    Odrv4 I__5294 (
            .O(N__30501),
            .I(n22374));
    CascadeMux I__5293 (
            .O(N__30498),
            .I(N__30495));
    InMux I__5292 (
            .O(N__30495),
            .I(N__30492));
    LocalMux I__5291 (
            .O(N__30492),
            .I(N__30489));
    Odrv4 I__5290 (
            .O(N__30489),
            .I(n21240));
    InMux I__5289 (
            .O(N__30486),
            .I(N__30483));
    LocalMux I__5288 (
            .O(N__30483),
            .I(N__30480));
    Odrv4 I__5287 (
            .O(N__30480),
            .I(n22401));
    InMux I__5286 (
            .O(N__30477),
            .I(N__30474));
    LocalMux I__5285 (
            .O(N__30474),
            .I(N__30471));
    Span4Mux_h I__5284 (
            .O(N__30471),
            .I(N__30468));
    Odrv4 I__5283 (
            .O(N__30468),
            .I(n21122));
    CascadeMux I__5282 (
            .O(N__30465),
            .I(n21122_cascade_));
    CascadeMux I__5281 (
            .O(N__30462),
            .I(n12610_cascade_));
    InMux I__5280 (
            .O(N__30459),
            .I(N__30456));
    LocalMux I__5279 (
            .O(N__30456),
            .I(N__30453));
    Span4Mux_v I__5278 (
            .O(N__30453),
            .I(N__30450));
    Span4Mux_h I__5277 (
            .O(N__30450),
            .I(N__30447));
    Odrv4 I__5276 (
            .O(N__30447),
            .I(buf_data_iac_5));
    InMux I__5275 (
            .O(N__30444),
            .I(N__30441));
    LocalMux I__5274 (
            .O(N__30441),
            .I(N__30438));
    Odrv12 I__5273 (
            .O(N__30438),
            .I(n22_adj_1604));
    InMux I__5272 (
            .O(N__30435),
            .I(n19974));
    InMux I__5271 (
            .O(N__30432),
            .I(n19975));
    InMux I__5270 (
            .O(N__30429),
            .I(n19976));
    InMux I__5269 (
            .O(N__30426),
            .I(n19977));
    InMux I__5268 (
            .O(N__30423),
            .I(N__30419));
    InMux I__5267 (
            .O(N__30422),
            .I(N__30416));
    LocalMux I__5266 (
            .O(N__30419),
            .I(N__30413));
    LocalMux I__5265 (
            .O(N__30416),
            .I(secclk_cnt_21));
    Odrv4 I__5264 (
            .O(N__30413),
            .I(secclk_cnt_21));
    InMux I__5263 (
            .O(N__30408),
            .I(N__30404));
    InMux I__5262 (
            .O(N__30407),
            .I(N__30401));
    LocalMux I__5261 (
            .O(N__30404),
            .I(secclk_cnt_19));
    LocalMux I__5260 (
            .O(N__30401),
            .I(secclk_cnt_19));
    CascadeMux I__5259 (
            .O(N__30396),
            .I(N__30393));
    InMux I__5258 (
            .O(N__30393),
            .I(N__30389));
    InMux I__5257 (
            .O(N__30392),
            .I(N__30386));
    LocalMux I__5256 (
            .O(N__30389),
            .I(N__30383));
    LocalMux I__5255 (
            .O(N__30386),
            .I(secclk_cnt_12));
    Odrv4 I__5254 (
            .O(N__30383),
            .I(secclk_cnt_12));
    InMux I__5253 (
            .O(N__30378),
            .I(N__30374));
    InMux I__5252 (
            .O(N__30377),
            .I(N__30371));
    LocalMux I__5251 (
            .O(N__30374),
            .I(secclk_cnt_22));
    LocalMux I__5250 (
            .O(N__30371),
            .I(secclk_cnt_22));
    InMux I__5249 (
            .O(N__30366),
            .I(N__30363));
    LocalMux I__5248 (
            .O(N__30363),
            .I(N__30360));
    Span4Mux_h I__5247 (
            .O(N__30360),
            .I(N__30356));
    InMux I__5246 (
            .O(N__30359),
            .I(N__30353));
    Span4Mux_h I__5245 (
            .O(N__30356),
            .I(N__30348));
    LocalMux I__5244 (
            .O(N__30353),
            .I(N__30348));
    Odrv4 I__5243 (
            .O(N__30348),
            .I(n14_adj_1571));
    InMux I__5242 (
            .O(N__30345),
            .I(n19965));
    InMux I__5241 (
            .O(N__30342),
            .I(n19966));
    InMux I__5240 (
            .O(N__30339),
            .I(n19967));
    InMux I__5239 (
            .O(N__30336),
            .I(n19968));
    InMux I__5238 (
            .O(N__30333),
            .I(n19969));
    InMux I__5237 (
            .O(N__30330),
            .I(n19970));
    InMux I__5236 (
            .O(N__30327),
            .I(bfn_11_9_0_));
    InMux I__5235 (
            .O(N__30324),
            .I(n19972));
    InMux I__5234 (
            .O(N__30321),
            .I(n19973));
    InMux I__5233 (
            .O(N__30318),
            .I(n19956));
    InMux I__5232 (
            .O(N__30315),
            .I(n19957));
    InMux I__5231 (
            .O(N__30312),
            .I(n19958));
    InMux I__5230 (
            .O(N__30309),
            .I(n19959));
    InMux I__5229 (
            .O(N__30306),
            .I(n19960));
    InMux I__5228 (
            .O(N__30303),
            .I(n19961));
    InMux I__5227 (
            .O(N__30300),
            .I(n19962));
    InMux I__5226 (
            .O(N__30297),
            .I(bfn_11_8_0_));
    InMux I__5225 (
            .O(N__30294),
            .I(n19964));
    InMux I__5224 (
            .O(N__30291),
            .I(N__30288));
    LocalMux I__5223 (
            .O(N__30288),
            .I(\ADC_VDC.n22587 ));
    InMux I__5222 (
            .O(N__30285),
            .I(N__30282));
    LocalMux I__5221 (
            .O(N__30282),
            .I(\ADC_VDC.n10708 ));
    CascadeMux I__5220 (
            .O(N__30279),
            .I(N__30275));
    InMux I__5219 (
            .O(N__30278),
            .I(N__30271));
    InMux I__5218 (
            .O(N__30275),
            .I(N__30268));
    CascadeMux I__5217 (
            .O(N__30274),
            .I(N__30265));
    LocalMux I__5216 (
            .O(N__30271),
            .I(N__30262));
    LocalMux I__5215 (
            .O(N__30268),
            .I(N__30259));
    InMux I__5214 (
            .O(N__30265),
            .I(N__30256));
    Span4Mux_v I__5213 (
            .O(N__30262),
            .I(N__30251));
    Span4Mux_v I__5212 (
            .O(N__30259),
            .I(N__30251));
    LocalMux I__5211 (
            .O(N__30256),
            .I(cmd_rdadctmp_22_adj_1501));
    Odrv4 I__5210 (
            .O(N__30251),
            .I(cmd_rdadctmp_22_adj_1501));
    CascadeMux I__5209 (
            .O(N__30246),
            .I(\ADC_VDC.n10708_cascade_ ));
    CascadeMux I__5208 (
            .O(N__30243),
            .I(N__30240));
    InMux I__5207 (
            .O(N__30240),
            .I(N__30237));
    LocalMux I__5206 (
            .O(N__30237),
            .I(N__30233));
    InMux I__5205 (
            .O(N__30236),
            .I(N__30230));
    Span4Mux_v I__5204 (
            .O(N__30233),
            .I(N__30227));
    LocalMux I__5203 (
            .O(N__30230),
            .I(\ADC_VDC.cmd_rdadctmp_23 ));
    Odrv4 I__5202 (
            .O(N__30227),
            .I(\ADC_VDC.cmd_rdadctmp_23 ));
    SRMux I__5201 (
            .O(N__30222),
            .I(N__30219));
    LocalMux I__5200 (
            .O(N__30219),
            .I(N__30216));
    Span4Mux_v I__5199 (
            .O(N__30216),
            .I(N__30213));
    Odrv4 I__5198 (
            .O(N__30213),
            .I(\ADC_VDC.n5 ));
    InMux I__5197 (
            .O(N__30210),
            .I(N__30206));
    InMux I__5196 (
            .O(N__30209),
            .I(N__30203));
    LocalMux I__5195 (
            .O(N__30206),
            .I(\ADC_VDC.avg_cnt_9 ));
    LocalMux I__5194 (
            .O(N__30203),
            .I(\ADC_VDC.avg_cnt_9 ));
    InMux I__5193 (
            .O(N__30198),
            .I(N__30194));
    InMux I__5192 (
            .O(N__30197),
            .I(N__30191));
    LocalMux I__5191 (
            .O(N__30194),
            .I(\ADC_VDC.avg_cnt_8 ));
    LocalMux I__5190 (
            .O(N__30191),
            .I(\ADC_VDC.avg_cnt_8 ));
    CascadeMux I__5189 (
            .O(N__30186),
            .I(N__30182));
    InMux I__5188 (
            .O(N__30185),
            .I(N__30179));
    InMux I__5187 (
            .O(N__30182),
            .I(N__30176));
    LocalMux I__5186 (
            .O(N__30179),
            .I(\ADC_VDC.avg_cnt_6 ));
    LocalMux I__5185 (
            .O(N__30176),
            .I(\ADC_VDC.avg_cnt_6 ));
    InMux I__5184 (
            .O(N__30171),
            .I(N__30167));
    InMux I__5183 (
            .O(N__30170),
            .I(N__30164));
    LocalMux I__5182 (
            .O(N__30167),
            .I(\ADC_VDC.avg_cnt_3 ));
    LocalMux I__5181 (
            .O(N__30164),
            .I(\ADC_VDC.avg_cnt_3 ));
    InMux I__5180 (
            .O(N__30159),
            .I(N__30156));
    LocalMux I__5179 (
            .O(N__30156),
            .I(N__30153));
    Span4Mux_h I__5178 (
            .O(N__30153),
            .I(N__30150));
    Odrv4 I__5177 (
            .O(N__30150),
            .I(\ADC_VDC.n20 ));
    CEMux I__5176 (
            .O(N__30147),
            .I(N__30144));
    LocalMux I__5175 (
            .O(N__30144),
            .I(N__30140));
    CEMux I__5174 (
            .O(N__30143),
            .I(N__30137));
    Span4Mux_h I__5173 (
            .O(N__30140),
            .I(N__30132));
    LocalMux I__5172 (
            .O(N__30137),
            .I(N__30132));
    Span4Mux_v I__5171 (
            .O(N__30132),
            .I(N__30129));
    Span4Mux_v I__5170 (
            .O(N__30129),
            .I(N__30126));
    Odrv4 I__5169 (
            .O(N__30126),
            .I(\CLK_DDS.n13005 ));
    CEMux I__5168 (
            .O(N__30123),
            .I(N__30120));
    LocalMux I__5167 (
            .O(N__30120),
            .I(N__30117));
    Odrv12 I__5166 (
            .O(N__30117),
            .I(\CLK_DDS.n9_adj_1433 ));
    CascadeMux I__5165 (
            .O(N__30114),
            .I(N__30111));
    InMux I__5164 (
            .O(N__30111),
            .I(N__30090));
    InMux I__5163 (
            .O(N__30110),
            .I(N__30075));
    InMux I__5162 (
            .O(N__30109),
            .I(N__30075));
    InMux I__5161 (
            .O(N__30108),
            .I(N__30075));
    InMux I__5160 (
            .O(N__30107),
            .I(N__30075));
    InMux I__5159 (
            .O(N__30106),
            .I(N__30075));
    InMux I__5158 (
            .O(N__30105),
            .I(N__30075));
    InMux I__5157 (
            .O(N__30104),
            .I(N__30075));
    InMux I__5156 (
            .O(N__30103),
            .I(N__30069));
    InMux I__5155 (
            .O(N__30102),
            .I(N__30066));
    InMux I__5154 (
            .O(N__30101),
            .I(N__30049));
    InMux I__5153 (
            .O(N__30100),
            .I(N__30049));
    InMux I__5152 (
            .O(N__30099),
            .I(N__30049));
    InMux I__5151 (
            .O(N__30098),
            .I(N__30049));
    InMux I__5150 (
            .O(N__30097),
            .I(N__30049));
    InMux I__5149 (
            .O(N__30096),
            .I(N__30049));
    InMux I__5148 (
            .O(N__30095),
            .I(N__30049));
    InMux I__5147 (
            .O(N__30094),
            .I(N__30049));
    InMux I__5146 (
            .O(N__30093),
            .I(N__30046));
    LocalMux I__5145 (
            .O(N__30090),
            .I(N__30042));
    LocalMux I__5144 (
            .O(N__30075),
            .I(N__30039));
    InMux I__5143 (
            .O(N__30074),
            .I(N__30032));
    InMux I__5142 (
            .O(N__30073),
            .I(N__30032));
    InMux I__5141 (
            .O(N__30072),
            .I(N__30032));
    LocalMux I__5140 (
            .O(N__30069),
            .I(N__30026));
    LocalMux I__5139 (
            .O(N__30066),
            .I(N__30026));
    LocalMux I__5138 (
            .O(N__30049),
            .I(N__30023));
    LocalMux I__5137 (
            .O(N__30046),
            .I(N__30020));
    CascadeMux I__5136 (
            .O(N__30045),
            .I(N__30017));
    Span4Mux_v I__5135 (
            .O(N__30042),
            .I(N__30011));
    Span4Mux_v I__5134 (
            .O(N__30039),
            .I(N__30011));
    LocalMux I__5133 (
            .O(N__30032),
            .I(N__30008));
    CascadeMux I__5132 (
            .O(N__30031),
            .I(N__30004));
    Span4Mux_v I__5131 (
            .O(N__30026),
            .I(N__30001));
    Span4Mux_v I__5130 (
            .O(N__30023),
            .I(N__29998));
    Span4Mux_h I__5129 (
            .O(N__30020),
            .I(N__29995));
    InMux I__5128 (
            .O(N__30017),
            .I(N__29990));
    InMux I__5127 (
            .O(N__30016),
            .I(N__29990));
    Span4Mux_v I__5126 (
            .O(N__30011),
            .I(N__29987));
    Sp12to4 I__5125 (
            .O(N__30008),
            .I(N__29984));
    InMux I__5124 (
            .O(N__30007),
            .I(N__29981));
    InMux I__5123 (
            .O(N__30004),
            .I(N__29978));
    Span4Mux_h I__5122 (
            .O(N__30001),
            .I(N__29973));
    Span4Mux_h I__5121 (
            .O(N__29998),
            .I(N__29973));
    Span4Mux_h I__5120 (
            .O(N__29995),
            .I(N__29968));
    LocalMux I__5119 (
            .O(N__29990),
            .I(N__29968));
    Sp12to4 I__5118 (
            .O(N__29987),
            .I(N__29963));
    Span12Mux_v I__5117 (
            .O(N__29984),
            .I(N__29963));
    LocalMux I__5116 (
            .O(N__29981),
            .I(dds_state_2_adj_1494));
    LocalMux I__5115 (
            .O(N__29978),
            .I(dds_state_2_adj_1494));
    Odrv4 I__5114 (
            .O(N__29973),
            .I(dds_state_2_adj_1494));
    Odrv4 I__5113 (
            .O(N__29968),
            .I(dds_state_2_adj_1494));
    Odrv12 I__5112 (
            .O(N__29963),
            .I(dds_state_2_adj_1494));
    CascadeMux I__5111 (
            .O(N__29952),
            .I(N__29948));
    InMux I__5110 (
            .O(N__29951),
            .I(N__29943));
    InMux I__5109 (
            .O(N__29948),
            .I(N__29934));
    InMux I__5108 (
            .O(N__29947),
            .I(N__29934));
    InMux I__5107 (
            .O(N__29946),
            .I(N__29934));
    LocalMux I__5106 (
            .O(N__29943),
            .I(N__29931));
    InMux I__5105 (
            .O(N__29942),
            .I(N__29928));
    InMux I__5104 (
            .O(N__29941),
            .I(N__29925));
    LocalMux I__5103 (
            .O(N__29934),
            .I(N__29922));
    Span4Mux_h I__5102 (
            .O(N__29931),
            .I(N__29919));
    LocalMux I__5101 (
            .O(N__29928),
            .I(N__29914));
    LocalMux I__5100 (
            .O(N__29925),
            .I(N__29914));
    Span4Mux_v I__5099 (
            .O(N__29922),
            .I(N__29911));
    Span4Mux_h I__5098 (
            .O(N__29919),
            .I(N__29904));
    Span4Mux_v I__5097 (
            .O(N__29914),
            .I(N__29899));
    Span4Mux_h I__5096 (
            .O(N__29911),
            .I(N__29899));
    InMux I__5095 (
            .O(N__29910),
            .I(N__29894));
    InMux I__5094 (
            .O(N__29909),
            .I(N__29894));
    InMux I__5093 (
            .O(N__29908),
            .I(N__29889));
    InMux I__5092 (
            .O(N__29907),
            .I(N__29889));
    Odrv4 I__5091 (
            .O(N__29904),
            .I(dds_state_0_adj_1496));
    Odrv4 I__5090 (
            .O(N__29899),
            .I(dds_state_0_adj_1496));
    LocalMux I__5089 (
            .O(N__29894),
            .I(dds_state_0_adj_1496));
    LocalMux I__5088 (
            .O(N__29889),
            .I(dds_state_0_adj_1496));
    InMux I__5087 (
            .O(N__29880),
            .I(N__29855));
    InMux I__5086 (
            .O(N__29879),
            .I(N__29855));
    InMux I__5085 (
            .O(N__29878),
            .I(N__29855));
    InMux I__5084 (
            .O(N__29877),
            .I(N__29855));
    InMux I__5083 (
            .O(N__29876),
            .I(N__29855));
    InMux I__5082 (
            .O(N__29875),
            .I(N__29855));
    InMux I__5081 (
            .O(N__29874),
            .I(N__29855));
    InMux I__5080 (
            .O(N__29873),
            .I(N__29855));
    CascadeMux I__5079 (
            .O(N__29872),
            .I(N__29848));
    LocalMux I__5078 (
            .O(N__29855),
            .I(N__29841));
    InMux I__5077 (
            .O(N__29854),
            .I(N__29823));
    InMux I__5076 (
            .O(N__29853),
            .I(N__29823));
    InMux I__5075 (
            .O(N__29852),
            .I(N__29823));
    InMux I__5074 (
            .O(N__29851),
            .I(N__29823));
    InMux I__5073 (
            .O(N__29848),
            .I(N__29823));
    InMux I__5072 (
            .O(N__29847),
            .I(N__29823));
    InMux I__5071 (
            .O(N__29846),
            .I(N__29823));
    InMux I__5070 (
            .O(N__29845),
            .I(N__29823));
    SRMux I__5069 (
            .O(N__29844),
            .I(N__29816));
    Span4Mux_h I__5068 (
            .O(N__29841),
            .I(N__29813));
    InMux I__5067 (
            .O(N__29840),
            .I(N__29810));
    LocalMux I__5066 (
            .O(N__29823),
            .I(N__29807));
    InMux I__5065 (
            .O(N__29822),
            .I(N__29804));
    CEMux I__5064 (
            .O(N__29821),
            .I(N__29801));
    InMux I__5063 (
            .O(N__29820),
            .I(N__29798));
    InMux I__5062 (
            .O(N__29819),
            .I(N__29795));
    LocalMux I__5061 (
            .O(N__29816),
            .I(N__29787));
    Span4Mux_v I__5060 (
            .O(N__29813),
            .I(N__29782));
    LocalMux I__5059 (
            .O(N__29810),
            .I(N__29782));
    Span4Mux_v I__5058 (
            .O(N__29807),
            .I(N__29777));
    LocalMux I__5057 (
            .O(N__29804),
            .I(N__29777));
    LocalMux I__5056 (
            .O(N__29801),
            .I(N__29774));
    LocalMux I__5055 (
            .O(N__29798),
            .I(N__29771));
    LocalMux I__5054 (
            .O(N__29795),
            .I(N__29768));
    InMux I__5053 (
            .O(N__29794),
            .I(N__29760));
    InMux I__5052 (
            .O(N__29793),
            .I(N__29760));
    InMux I__5051 (
            .O(N__29792),
            .I(N__29760));
    InMux I__5050 (
            .O(N__29791),
            .I(N__29755));
    InMux I__5049 (
            .O(N__29790),
            .I(N__29755));
    Span4Mux_v I__5048 (
            .O(N__29787),
            .I(N__29750));
    Span4Mux_v I__5047 (
            .O(N__29782),
            .I(N__29750));
    Span4Mux_v I__5046 (
            .O(N__29777),
            .I(N__29747));
    Span4Mux_h I__5045 (
            .O(N__29774),
            .I(N__29742));
    Span4Mux_h I__5044 (
            .O(N__29771),
            .I(N__29742));
    Span4Mux_h I__5043 (
            .O(N__29768),
            .I(N__29739));
    InMux I__5042 (
            .O(N__29767),
            .I(N__29736));
    LocalMux I__5041 (
            .O(N__29760),
            .I(N__29731));
    LocalMux I__5040 (
            .O(N__29755),
            .I(N__29731));
    Odrv4 I__5039 (
            .O(N__29750),
            .I(dds_state_1_adj_1495));
    Odrv4 I__5038 (
            .O(N__29747),
            .I(dds_state_1_adj_1495));
    Odrv4 I__5037 (
            .O(N__29742),
            .I(dds_state_1_adj_1495));
    Odrv4 I__5036 (
            .O(N__29739),
            .I(dds_state_1_adj_1495));
    LocalMux I__5035 (
            .O(N__29736),
            .I(dds_state_1_adj_1495));
    Odrv12 I__5034 (
            .O(N__29731),
            .I(dds_state_1_adj_1495));
    CEMux I__5033 (
            .O(N__29718),
            .I(N__29715));
    LocalMux I__5032 (
            .O(N__29715),
            .I(N__29712));
    Span4Mux_v I__5031 (
            .O(N__29712),
            .I(N__29708));
    CEMux I__5030 (
            .O(N__29711),
            .I(N__29705));
    Span4Mux_h I__5029 (
            .O(N__29708),
            .I(N__29702));
    LocalMux I__5028 (
            .O(N__29705),
            .I(N__29699));
    Odrv4 I__5027 (
            .O(N__29702),
            .I(\CLK_DDS.n9 ));
    Odrv12 I__5026 (
            .O(N__29699),
            .I(\CLK_DDS.n9 ));
    InMux I__5025 (
            .O(N__29694),
            .I(bfn_11_7_0_));
    CascadeMux I__5024 (
            .O(N__29691),
            .I(\ADC_VDC.n7_cascade_ ));
    InMux I__5023 (
            .O(N__29688),
            .I(N__29683));
    InMux I__5022 (
            .O(N__29687),
            .I(N__29680));
    InMux I__5021 (
            .O(N__29686),
            .I(N__29677));
    LocalMux I__5020 (
            .O(N__29683),
            .I(\ADC_VDC.n21193 ));
    LocalMux I__5019 (
            .O(N__29680),
            .I(\ADC_VDC.n21193 ));
    LocalMux I__5018 (
            .O(N__29677),
            .I(\ADC_VDC.n21193 ));
    InMux I__5017 (
            .O(N__29670),
            .I(N__29667));
    LocalMux I__5016 (
            .O(N__29667),
            .I(N__29663));
    CascadeMux I__5015 (
            .O(N__29666),
            .I(N__29660));
    Span4Mux_h I__5014 (
            .O(N__29663),
            .I(N__29657));
    InMux I__5013 (
            .O(N__29660),
            .I(N__29654));
    Odrv4 I__5012 (
            .O(N__29657),
            .I(cmd_rdadcbuf_19));
    LocalMux I__5011 (
            .O(N__29654),
            .I(cmd_rdadcbuf_19));
    InMux I__5010 (
            .O(N__29649),
            .I(N__29646));
    LocalMux I__5009 (
            .O(N__29646),
            .I(N__29643));
    Span4Mux_h I__5008 (
            .O(N__29643),
            .I(N__29639));
    InMux I__5007 (
            .O(N__29642),
            .I(N__29636));
    Odrv4 I__5006 (
            .O(N__29639),
            .I(cmd_rdadcbuf_24));
    LocalMux I__5005 (
            .O(N__29636),
            .I(cmd_rdadcbuf_24));
    InMux I__5004 (
            .O(N__29631),
            .I(N__29628));
    LocalMux I__5003 (
            .O(N__29628),
            .I(N__29625));
    Span4Mux_v I__5002 (
            .O(N__29625),
            .I(N__29622));
    Span4Mux_v I__5001 (
            .O(N__29622),
            .I(N__29618));
    InMux I__5000 (
            .O(N__29621),
            .I(N__29615));
    Odrv4 I__4999 (
            .O(N__29618),
            .I(buf_adcdata_vdc_13));
    LocalMux I__4998 (
            .O(N__29615),
            .I(buf_adcdata_vdc_13));
    InMux I__4997 (
            .O(N__29610),
            .I(N__29607));
    LocalMux I__4996 (
            .O(N__29607),
            .I(N__29604));
    Span4Mux_h I__4995 (
            .O(N__29604),
            .I(N__29601));
    Span4Mux_v I__4994 (
            .O(N__29601),
            .I(N__29597));
    InMux I__4993 (
            .O(N__29600),
            .I(N__29594));
    Odrv4 I__4992 (
            .O(N__29597),
            .I(cmd_rdadcbuf_30));
    LocalMux I__4991 (
            .O(N__29594),
            .I(cmd_rdadcbuf_30));
    InMux I__4990 (
            .O(N__29589),
            .I(N__29586));
    LocalMux I__4989 (
            .O(N__29586),
            .I(N__29583));
    Span12Mux_h I__4988 (
            .O(N__29583),
            .I(N__29579));
    InMux I__4987 (
            .O(N__29582),
            .I(N__29576));
    Odrv12 I__4986 (
            .O(N__29579),
            .I(buf_adcdata_vdc_19));
    LocalMux I__4985 (
            .O(N__29576),
            .I(buf_adcdata_vdc_19));
    InMux I__4984 (
            .O(N__29571),
            .I(N__29568));
    LocalMux I__4983 (
            .O(N__29568),
            .I(N__29565));
    Span4Mux_h I__4982 (
            .O(N__29565),
            .I(N__29561));
    InMux I__4981 (
            .O(N__29564),
            .I(N__29558));
    Odrv4 I__4980 (
            .O(N__29561),
            .I(cmd_rdadcbuf_28));
    LocalMux I__4979 (
            .O(N__29558),
            .I(cmd_rdadcbuf_28));
    InMux I__4978 (
            .O(N__29553),
            .I(N__29550));
    LocalMux I__4977 (
            .O(N__29550),
            .I(N__29547));
    Span4Mux_h I__4976 (
            .O(N__29547),
            .I(N__29544));
    Span4Mux_v I__4975 (
            .O(N__29544),
            .I(N__29541));
    Sp12to4 I__4974 (
            .O(N__29541),
            .I(N__29537));
    InMux I__4973 (
            .O(N__29540),
            .I(N__29534));
    Odrv12 I__4972 (
            .O(N__29537),
            .I(buf_adcdata_vdc_17));
    LocalMux I__4971 (
            .O(N__29534),
            .I(buf_adcdata_vdc_17));
    InMux I__4970 (
            .O(N__29529),
            .I(N__29526));
    LocalMux I__4969 (
            .O(N__29526),
            .I(N__29523));
    Span4Mux_v I__4968 (
            .O(N__29523),
            .I(N__29520));
    Span4Mux_h I__4967 (
            .O(N__29520),
            .I(N__29516));
    InMux I__4966 (
            .O(N__29519),
            .I(N__29513));
    Odrv4 I__4965 (
            .O(N__29516),
            .I(cmd_rdadcbuf_32));
    LocalMux I__4964 (
            .O(N__29513),
            .I(cmd_rdadcbuf_32));
    InMux I__4963 (
            .O(N__29508),
            .I(N__29505));
    LocalMux I__4962 (
            .O(N__29505),
            .I(N__29502));
    Span4Mux_v I__4961 (
            .O(N__29502),
            .I(N__29498));
    CascadeMux I__4960 (
            .O(N__29501),
            .I(N__29495));
    Span4Mux_h I__4959 (
            .O(N__29498),
            .I(N__29492));
    InMux I__4958 (
            .O(N__29495),
            .I(N__29489));
    Odrv4 I__4957 (
            .O(N__29492),
            .I(buf_adcdata_vdc_21));
    LocalMux I__4956 (
            .O(N__29489),
            .I(buf_adcdata_vdc_21));
    InMux I__4955 (
            .O(N__29484),
            .I(N__29481));
    LocalMux I__4954 (
            .O(N__29481),
            .I(N__29478));
    Span4Mux_h I__4953 (
            .O(N__29478),
            .I(N__29475));
    Span4Mux_v I__4952 (
            .O(N__29475),
            .I(N__29471));
    InMux I__4951 (
            .O(N__29474),
            .I(N__29468));
    Odrv4 I__4950 (
            .O(N__29471),
            .I(cmd_rdadcbuf_31));
    LocalMux I__4949 (
            .O(N__29468),
            .I(cmd_rdadcbuf_31));
    InMux I__4948 (
            .O(N__29463),
            .I(N__29460));
    LocalMux I__4947 (
            .O(N__29460),
            .I(N__29457));
    Span4Mux_v I__4946 (
            .O(N__29457),
            .I(N__29453));
    InMux I__4945 (
            .O(N__29456),
            .I(N__29449));
    Span4Mux_h I__4944 (
            .O(N__29453),
            .I(N__29446));
    InMux I__4943 (
            .O(N__29452),
            .I(N__29443));
    LocalMux I__4942 (
            .O(N__29449),
            .I(N__29440));
    Span4Mux_v I__4941 (
            .O(N__29446),
            .I(N__29437));
    LocalMux I__4940 (
            .O(N__29443),
            .I(buf_dds1_4));
    Odrv4 I__4939 (
            .O(N__29440),
            .I(buf_dds1_4));
    Odrv4 I__4938 (
            .O(N__29437),
            .I(buf_dds1_4));
    CascadeMux I__4937 (
            .O(N__29430),
            .I(N__29425));
    CascadeMux I__4936 (
            .O(N__29429),
            .I(N__29422));
    CascadeMux I__4935 (
            .O(N__29428),
            .I(N__29419));
    InMux I__4934 (
            .O(N__29425),
            .I(N__29416));
    InMux I__4933 (
            .O(N__29422),
            .I(N__29413));
    InMux I__4932 (
            .O(N__29419),
            .I(N__29410));
    LocalMux I__4931 (
            .O(N__29416),
            .I(N__29407));
    LocalMux I__4930 (
            .O(N__29413),
            .I(N__29402));
    LocalMux I__4929 (
            .O(N__29410),
            .I(N__29402));
    Span4Mux_h I__4928 (
            .O(N__29407),
            .I(N__29399));
    Odrv4 I__4927 (
            .O(N__29402),
            .I(cmd_rdadctmp_20));
    Odrv4 I__4926 (
            .O(N__29399),
            .I(cmd_rdadctmp_20));
    CascadeMux I__4925 (
            .O(N__29394),
            .I(N__29387));
    InMux I__4924 (
            .O(N__29393),
            .I(N__29375));
    InMux I__4923 (
            .O(N__29392),
            .I(N__29375));
    CascadeMux I__4922 (
            .O(N__29391),
            .I(N__29369));
    CascadeMux I__4921 (
            .O(N__29390),
            .I(N__29366));
    InMux I__4920 (
            .O(N__29387),
            .I(N__29357));
    InMux I__4919 (
            .O(N__29386),
            .I(N__29357));
    InMux I__4918 (
            .O(N__29385),
            .I(N__29354));
    InMux I__4917 (
            .O(N__29384),
            .I(N__29349));
    InMux I__4916 (
            .O(N__29383),
            .I(N__29349));
    InMux I__4915 (
            .O(N__29382),
            .I(N__29344));
    InMux I__4914 (
            .O(N__29381),
            .I(N__29344));
    InMux I__4913 (
            .O(N__29380),
            .I(N__29341));
    LocalMux I__4912 (
            .O(N__29375),
            .I(N__29338));
    CascadeMux I__4911 (
            .O(N__29374),
            .I(N__29329));
    InMux I__4910 (
            .O(N__29373),
            .I(N__29320));
    InMux I__4909 (
            .O(N__29372),
            .I(N__29313));
    InMux I__4908 (
            .O(N__29369),
            .I(N__29313));
    InMux I__4907 (
            .O(N__29366),
            .I(N__29313));
    InMux I__4906 (
            .O(N__29365),
            .I(N__29308));
    InMux I__4905 (
            .O(N__29364),
            .I(N__29308));
    InMux I__4904 (
            .O(N__29363),
            .I(N__29303));
    InMux I__4903 (
            .O(N__29362),
            .I(N__29303));
    LocalMux I__4902 (
            .O(N__29357),
            .I(N__29298));
    LocalMux I__4901 (
            .O(N__29354),
            .I(N__29298));
    LocalMux I__4900 (
            .O(N__29349),
            .I(N__29295));
    LocalMux I__4899 (
            .O(N__29344),
            .I(N__29292));
    LocalMux I__4898 (
            .O(N__29341),
            .I(N__29287));
    Span4Mux_v I__4897 (
            .O(N__29338),
            .I(N__29287));
    InMux I__4896 (
            .O(N__29337),
            .I(N__29284));
    InMux I__4895 (
            .O(N__29336),
            .I(N__29277));
    InMux I__4894 (
            .O(N__29335),
            .I(N__29277));
    InMux I__4893 (
            .O(N__29334),
            .I(N__29277));
    InMux I__4892 (
            .O(N__29333),
            .I(N__29272));
    InMux I__4891 (
            .O(N__29332),
            .I(N__29272));
    InMux I__4890 (
            .O(N__29329),
            .I(N__29263));
    InMux I__4889 (
            .O(N__29328),
            .I(N__29263));
    InMux I__4888 (
            .O(N__29327),
            .I(N__29263));
    InMux I__4887 (
            .O(N__29326),
            .I(N__29263));
    InMux I__4886 (
            .O(N__29325),
            .I(N__29256));
    InMux I__4885 (
            .O(N__29324),
            .I(N__29256));
    InMux I__4884 (
            .O(N__29323),
            .I(N__29256));
    LocalMux I__4883 (
            .O(N__29320),
            .I(N__29249));
    LocalMux I__4882 (
            .O(N__29313),
            .I(N__29249));
    LocalMux I__4881 (
            .O(N__29308),
            .I(N__29249));
    LocalMux I__4880 (
            .O(N__29303),
            .I(N__29246));
    Span4Mux_h I__4879 (
            .O(N__29298),
            .I(N__29241));
    Span4Mux_v I__4878 (
            .O(N__29295),
            .I(N__29241));
    Span4Mux_h I__4877 (
            .O(N__29292),
            .I(N__29236));
    Span4Mux_v I__4876 (
            .O(N__29287),
            .I(N__29236));
    LocalMux I__4875 (
            .O(N__29284),
            .I(n12771));
    LocalMux I__4874 (
            .O(N__29277),
            .I(n12771));
    LocalMux I__4873 (
            .O(N__29272),
            .I(n12771));
    LocalMux I__4872 (
            .O(N__29263),
            .I(n12771));
    LocalMux I__4871 (
            .O(N__29256),
            .I(n12771));
    Odrv4 I__4870 (
            .O(N__29249),
            .I(n12771));
    Odrv12 I__4869 (
            .O(N__29246),
            .I(n12771));
    Odrv4 I__4868 (
            .O(N__29241),
            .I(n12771));
    Odrv4 I__4867 (
            .O(N__29236),
            .I(n12771));
    CascadeMux I__4866 (
            .O(N__29217),
            .I(N__29214));
    InMux I__4865 (
            .O(N__29214),
            .I(N__29210));
    InMux I__4864 (
            .O(N__29213),
            .I(N__29207));
    LocalMux I__4863 (
            .O(N__29210),
            .I(cmd_rdadctmp_31));
    LocalMux I__4862 (
            .O(N__29207),
            .I(cmd_rdadctmp_31));
    CascadeMux I__4861 (
            .O(N__29202),
            .I(N__29198));
    InMux I__4860 (
            .O(N__29201),
            .I(N__29195));
    InMux I__4859 (
            .O(N__29198),
            .I(N__29192));
    LocalMux I__4858 (
            .O(N__29195),
            .I(N__29189));
    LocalMux I__4857 (
            .O(N__29192),
            .I(N__29185));
    Span12Mux_h I__4856 (
            .O(N__29189),
            .I(N__29182));
    InMux I__4855 (
            .O(N__29188),
            .I(N__29179));
    Span4Mux_v I__4854 (
            .O(N__29185),
            .I(N__29176));
    Span12Mux_v I__4853 (
            .O(N__29182),
            .I(N__29173));
    LocalMux I__4852 (
            .O(N__29179),
            .I(buf_adcdata_iac_23));
    Odrv4 I__4851 (
            .O(N__29176),
            .I(buf_adcdata_iac_23));
    Odrv12 I__4850 (
            .O(N__29173),
            .I(buf_adcdata_iac_23));
    CEMux I__4849 (
            .O(N__29166),
            .I(N__29163));
    LocalMux I__4848 (
            .O(N__29163),
            .I(N__29160));
    Span4Mux_v I__4847 (
            .O(N__29160),
            .I(N__29157));
    Odrv4 I__4846 (
            .O(N__29157),
            .I(\ADC_VDC.n16 ));
    CascadeMux I__4845 (
            .O(N__29154),
            .I(\ADC_VDC.n21593_cascade_ ));
    CascadeMux I__4844 (
            .O(N__29151),
            .I(\ADC_VDC.n21590_cascade_ ));
    InMux I__4843 (
            .O(N__29148),
            .I(N__29145));
    LocalMux I__4842 (
            .O(N__29145),
            .I(\ADC_VDC.n22590 ));
    CascadeMux I__4841 (
            .O(N__29142),
            .I(N__29131));
    CascadeMux I__4840 (
            .O(N__29141),
            .I(N__29128));
    CascadeMux I__4839 (
            .O(N__29140),
            .I(N__29125));
    CascadeMux I__4838 (
            .O(N__29139),
            .I(N__29122));
    CascadeMux I__4837 (
            .O(N__29138),
            .I(N__29119));
    InMux I__4836 (
            .O(N__29137),
            .I(N__29097));
    InMux I__4835 (
            .O(N__29136),
            .I(N__29097));
    InMux I__4834 (
            .O(N__29135),
            .I(N__29097));
    InMux I__4833 (
            .O(N__29134),
            .I(N__29097));
    InMux I__4832 (
            .O(N__29131),
            .I(N__29097));
    InMux I__4831 (
            .O(N__29128),
            .I(N__29097));
    InMux I__4830 (
            .O(N__29125),
            .I(N__29097));
    InMux I__4829 (
            .O(N__29122),
            .I(N__29097));
    InMux I__4828 (
            .O(N__29119),
            .I(N__29094));
    CascadeMux I__4827 (
            .O(N__29118),
            .I(N__29088));
    CascadeMux I__4826 (
            .O(N__29117),
            .I(N__29085));
    CascadeMux I__4825 (
            .O(N__29116),
            .I(N__29077));
    CascadeMux I__4824 (
            .O(N__29115),
            .I(N__29074));
    CascadeMux I__4823 (
            .O(N__29114),
            .I(N__29071));
    LocalMux I__4822 (
            .O(N__29097),
            .I(N__29067));
    LocalMux I__4821 (
            .O(N__29094),
            .I(N__29064));
    InMux I__4820 (
            .O(N__29093),
            .I(N__29047));
    InMux I__4819 (
            .O(N__29092),
            .I(N__29047));
    InMux I__4818 (
            .O(N__29091),
            .I(N__29047));
    InMux I__4817 (
            .O(N__29088),
            .I(N__29047));
    InMux I__4816 (
            .O(N__29085),
            .I(N__29047));
    InMux I__4815 (
            .O(N__29084),
            .I(N__29047));
    InMux I__4814 (
            .O(N__29083),
            .I(N__29047));
    InMux I__4813 (
            .O(N__29082),
            .I(N__29047));
    InMux I__4812 (
            .O(N__29081),
            .I(N__29034));
    InMux I__4811 (
            .O(N__29080),
            .I(N__29034));
    InMux I__4810 (
            .O(N__29077),
            .I(N__29034));
    InMux I__4809 (
            .O(N__29074),
            .I(N__29034));
    InMux I__4808 (
            .O(N__29071),
            .I(N__29034));
    InMux I__4807 (
            .O(N__29070),
            .I(N__29034));
    Span4Mux_h I__4806 (
            .O(N__29067),
            .I(N__29031));
    Span4Mux_h I__4805 (
            .O(N__29064),
            .I(N__29028));
    LocalMux I__4804 (
            .O(N__29047),
            .I(N__29023));
    LocalMux I__4803 (
            .O(N__29034),
            .I(N__29023));
    Sp12to4 I__4802 (
            .O(N__29031),
            .I(N__29020));
    Span4Mux_v I__4801 (
            .O(N__29028),
            .I(N__29017));
    Span4Mux_h I__4800 (
            .O(N__29023),
            .I(N__29014));
    Odrv12 I__4799 (
            .O(N__29020),
            .I(n13324));
    Odrv4 I__4798 (
            .O(N__29017),
            .I(n13324));
    Odrv4 I__4797 (
            .O(N__29014),
            .I(n13324));
    IoInMux I__4796 (
            .O(N__29007),
            .I(N__29004));
    LocalMux I__4795 (
            .O(N__29004),
            .I(N__29001));
    Span4Mux_s1_h I__4794 (
            .O(N__29001),
            .I(N__28998));
    Sp12to4 I__4793 (
            .O(N__28998),
            .I(N__28995));
    Span12Mux_s5_v I__4792 (
            .O(N__28995),
            .I(N__28991));
    InMux I__4791 (
            .O(N__28994),
            .I(N__28987));
    Span12Mux_h I__4790 (
            .O(N__28991),
            .I(N__28984));
    InMux I__4789 (
            .O(N__28990),
            .I(N__28981));
    LocalMux I__4788 (
            .O(N__28987),
            .I(N__28978));
    Odrv12 I__4787 (
            .O(N__28984),
            .I(VAC_FLT1));
    LocalMux I__4786 (
            .O(N__28981),
            .I(VAC_FLT1));
    Odrv4 I__4785 (
            .O(N__28978),
            .I(VAC_FLT1));
    CascadeMux I__4784 (
            .O(N__28971),
            .I(N__28968));
    InMux I__4783 (
            .O(N__28968),
            .I(N__28965));
    LocalMux I__4782 (
            .O(N__28965),
            .I(N__28962));
    Span4Mux_h I__4781 (
            .O(N__28962),
            .I(N__28957));
    InMux I__4780 (
            .O(N__28961),
            .I(N__28952));
    InMux I__4779 (
            .O(N__28960),
            .I(N__28952));
    Odrv4 I__4778 (
            .O(N__28957),
            .I(cmd_rdadctmp_29));
    LocalMux I__4777 (
            .O(N__28952),
            .I(cmd_rdadctmp_29));
    InMux I__4776 (
            .O(N__28947),
            .I(N__28944));
    LocalMux I__4775 (
            .O(N__28944),
            .I(N__28941));
    Span4Mux_h I__4774 (
            .O(N__28941),
            .I(N__28937));
    InMux I__4773 (
            .O(N__28940),
            .I(N__28934));
    Sp12to4 I__4772 (
            .O(N__28937),
            .I(N__28930));
    LocalMux I__4771 (
            .O(N__28934),
            .I(N__28927));
    InMux I__4770 (
            .O(N__28933),
            .I(N__28924));
    Span12Mux_v I__4769 (
            .O(N__28930),
            .I(N__28921));
    Span4Mux_v I__4768 (
            .O(N__28927),
            .I(N__28918));
    LocalMux I__4767 (
            .O(N__28924),
            .I(buf_adcdata_iac_21));
    Odrv12 I__4766 (
            .O(N__28921),
            .I(buf_adcdata_iac_21));
    Odrv4 I__4765 (
            .O(N__28918),
            .I(buf_adcdata_iac_21));
    CascadeMux I__4764 (
            .O(N__28911),
            .I(N__28908));
    InMux I__4763 (
            .O(N__28908),
            .I(N__28904));
    CascadeMux I__4762 (
            .O(N__28907),
            .I(N__28901));
    LocalMux I__4761 (
            .O(N__28904),
            .I(N__28897));
    InMux I__4760 (
            .O(N__28901),
            .I(N__28892));
    InMux I__4759 (
            .O(N__28900),
            .I(N__28892));
    Odrv4 I__4758 (
            .O(N__28897),
            .I(cmd_rdadctmp_28));
    LocalMux I__4757 (
            .O(N__28892),
            .I(cmd_rdadctmp_28));
    CascadeMux I__4756 (
            .O(N__28887),
            .I(N__28883));
    CascadeMux I__4755 (
            .O(N__28886),
            .I(N__28880));
    InMux I__4754 (
            .O(N__28883),
            .I(N__28876));
    InMux I__4753 (
            .O(N__28880),
            .I(N__28873));
    InMux I__4752 (
            .O(N__28879),
            .I(N__28870));
    LocalMux I__4751 (
            .O(N__28876),
            .I(cmd_rdadctmp_25));
    LocalMux I__4750 (
            .O(N__28873),
            .I(cmd_rdadctmp_25));
    LocalMux I__4749 (
            .O(N__28870),
            .I(cmd_rdadctmp_25));
    InMux I__4748 (
            .O(N__28863),
            .I(N__28859));
    InMux I__4747 (
            .O(N__28862),
            .I(N__28856));
    LocalMux I__4746 (
            .O(N__28859),
            .I(n17728));
    LocalMux I__4745 (
            .O(N__28856),
            .I(n17728));
    CascadeMux I__4744 (
            .O(N__28851),
            .I(n11_cascade_));
    InMux I__4743 (
            .O(N__28848),
            .I(N__28843));
    InMux I__4742 (
            .O(N__28847),
            .I(N__28840));
    InMux I__4741 (
            .O(N__28846),
            .I(N__28836));
    LocalMux I__4740 (
            .O(N__28843),
            .I(N__28833));
    LocalMux I__4739 (
            .O(N__28840),
            .I(N__28830));
    InMux I__4738 (
            .O(N__28839),
            .I(N__28827));
    LocalMux I__4737 (
            .O(N__28836),
            .I(N__28823));
    Span4Mux_h I__4736 (
            .O(N__28833),
            .I(N__28816));
    Span4Mux_v I__4735 (
            .O(N__28830),
            .I(N__28816));
    LocalMux I__4734 (
            .O(N__28827),
            .I(N__28816));
    InMux I__4733 (
            .O(N__28826),
            .I(N__28813));
    Odrv4 I__4732 (
            .O(N__28823),
            .I(acadc_dtrig_v));
    Odrv4 I__4731 (
            .O(N__28816),
            .I(acadc_dtrig_v));
    LocalMux I__4730 (
            .O(N__28813),
            .I(acadc_dtrig_v));
    InMux I__4729 (
            .O(N__28806),
            .I(N__28803));
    LocalMux I__4728 (
            .O(N__28803),
            .I(N__28798));
    InMux I__4727 (
            .O(N__28802),
            .I(N__28795));
    InMux I__4726 (
            .O(N__28801),
            .I(N__28792));
    Span4Mux_v I__4725 (
            .O(N__28798),
            .I(N__28787));
    LocalMux I__4724 (
            .O(N__28795),
            .I(N__28787));
    LocalMux I__4723 (
            .O(N__28792),
            .I(N__28782));
    Span4Mux_h I__4722 (
            .O(N__28787),
            .I(N__28779));
    InMux I__4721 (
            .O(N__28786),
            .I(N__28774));
    InMux I__4720 (
            .O(N__28785),
            .I(N__28774));
    Span4Mux_v I__4719 (
            .O(N__28782),
            .I(N__28771));
    Odrv4 I__4718 (
            .O(N__28779),
            .I(acadc_dtrig_i));
    LocalMux I__4717 (
            .O(N__28774),
            .I(acadc_dtrig_i));
    Odrv4 I__4716 (
            .O(N__28771),
            .I(acadc_dtrig_i));
    InMux I__4715 (
            .O(N__28764),
            .I(N__28761));
    LocalMux I__4714 (
            .O(N__28761),
            .I(eis_state_2_N_392_1));
    CascadeMux I__4713 (
            .O(N__28758),
            .I(eis_state_2_N_392_1_cascade_));
    CascadeMux I__4712 (
            .O(N__28755),
            .I(n2_adj_1696_cascade_));
    InMux I__4711 (
            .O(N__28752),
            .I(N__28749));
    LocalMux I__4710 (
            .O(N__28749),
            .I(n22437));
    InMux I__4709 (
            .O(N__28746),
            .I(N__28742));
    InMux I__4708 (
            .O(N__28745),
            .I(N__28739));
    LocalMux I__4707 (
            .O(N__28742),
            .I(N__28735));
    LocalMux I__4706 (
            .O(N__28739),
            .I(N__28732));
    InMux I__4705 (
            .O(N__28738),
            .I(N__28729));
    Odrv4 I__4704 (
            .O(N__28735),
            .I(cmd_rdadctmp_23));
    Odrv4 I__4703 (
            .O(N__28732),
            .I(cmd_rdadctmp_23));
    LocalMux I__4702 (
            .O(N__28729),
            .I(cmd_rdadctmp_23));
    InMux I__4701 (
            .O(N__28722),
            .I(N__28719));
    LocalMux I__4700 (
            .O(N__28719),
            .I(n22371));
    CascadeMux I__4699 (
            .O(N__28716),
            .I(n12_adj_1454_cascade_));
    InMux I__4698 (
            .O(N__28713),
            .I(N__28710));
    LocalMux I__4697 (
            .O(N__28710),
            .I(N__28705));
    InMux I__4696 (
            .O(N__28709),
            .I(N__28702));
    InMux I__4695 (
            .O(N__28708),
            .I(N__28699));
    Span4Mux_v I__4694 (
            .O(N__28705),
            .I(N__28692));
    LocalMux I__4693 (
            .O(N__28702),
            .I(N__28692));
    LocalMux I__4692 (
            .O(N__28699),
            .I(N__28689));
    InMux I__4691 (
            .O(N__28698),
            .I(N__28686));
    InMux I__4690 (
            .O(N__28697),
            .I(N__28683));
    Span4Mux_h I__4689 (
            .O(N__28692),
            .I(N__28680));
    Span4Mux_v I__4688 (
            .O(N__28689),
            .I(N__28677));
    LocalMux I__4687 (
            .O(N__28686),
            .I(N__28674));
    LocalMux I__4686 (
            .O(N__28683),
            .I(acadc_trig));
    Odrv4 I__4685 (
            .O(N__28680),
            .I(acadc_trig));
    Odrv4 I__4684 (
            .O(N__28677),
            .I(acadc_trig));
    Odrv12 I__4683 (
            .O(N__28674),
            .I(acadc_trig));
    CascadeMux I__4682 (
            .O(N__28665),
            .I(N__28661));
    InMux I__4681 (
            .O(N__28664),
            .I(N__28658));
    InMux I__4680 (
            .O(N__28661),
            .I(N__28655));
    LocalMux I__4679 (
            .O(N__28658),
            .I(n21053));
    LocalMux I__4678 (
            .O(N__28655),
            .I(n21053));
    CascadeMux I__4677 (
            .O(N__28650),
            .I(n21042_cascade_));
    CascadeMux I__4676 (
            .O(N__28647),
            .I(n21030_cascade_));
    InMux I__4675 (
            .O(N__28644),
            .I(N__28640));
    InMux I__4674 (
            .O(N__28643),
            .I(N__28637));
    LocalMux I__4673 (
            .O(N__28640),
            .I(eis_end));
    LocalMux I__4672 (
            .O(N__28637),
            .I(eis_end));
    SRMux I__4671 (
            .O(N__28632),
            .I(N__28628));
    SRMux I__4670 (
            .O(N__28631),
            .I(N__28623));
    LocalMux I__4669 (
            .O(N__28628),
            .I(N__28618));
    SRMux I__4668 (
            .O(N__28627),
            .I(N__28615));
    SRMux I__4667 (
            .O(N__28626),
            .I(N__28611));
    LocalMux I__4666 (
            .O(N__28623),
            .I(N__28607));
    SRMux I__4665 (
            .O(N__28622),
            .I(N__28604));
    SRMux I__4664 (
            .O(N__28621),
            .I(N__28599));
    Span4Mux_h I__4663 (
            .O(N__28618),
            .I(N__28596));
    LocalMux I__4662 (
            .O(N__28615),
            .I(N__28593));
    SRMux I__4661 (
            .O(N__28614),
            .I(N__28590));
    LocalMux I__4660 (
            .O(N__28611),
            .I(N__28587));
    SRMux I__4659 (
            .O(N__28610),
            .I(N__28584));
    Span4Mux_v I__4658 (
            .O(N__28607),
            .I(N__28579));
    LocalMux I__4657 (
            .O(N__28604),
            .I(N__28579));
    SRMux I__4656 (
            .O(N__28603),
            .I(N__28576));
    SRMux I__4655 (
            .O(N__28602),
            .I(N__28572));
    LocalMux I__4654 (
            .O(N__28599),
            .I(N__28568));
    Span4Mux_v I__4653 (
            .O(N__28596),
            .I(N__28563));
    Span4Mux_h I__4652 (
            .O(N__28593),
            .I(N__28563));
    LocalMux I__4651 (
            .O(N__28590),
            .I(N__28560));
    Span4Mux_v I__4650 (
            .O(N__28587),
            .I(N__28555));
    LocalMux I__4649 (
            .O(N__28584),
            .I(N__28555));
    Span4Mux_v I__4648 (
            .O(N__28579),
            .I(N__28550));
    LocalMux I__4647 (
            .O(N__28576),
            .I(N__28550));
    SRMux I__4646 (
            .O(N__28575),
            .I(N__28547));
    LocalMux I__4645 (
            .O(N__28572),
            .I(N__28544));
    SRMux I__4644 (
            .O(N__28571),
            .I(N__28541));
    Span4Mux_h I__4643 (
            .O(N__28568),
            .I(N__28538));
    Span4Mux_v I__4642 (
            .O(N__28563),
            .I(N__28533));
    Span4Mux_h I__4641 (
            .O(N__28560),
            .I(N__28533));
    Span4Mux_v I__4640 (
            .O(N__28555),
            .I(N__28528));
    Span4Mux_v I__4639 (
            .O(N__28550),
            .I(N__28528));
    LocalMux I__4638 (
            .O(N__28547),
            .I(N__28525));
    Span4Mux_v I__4637 (
            .O(N__28544),
            .I(N__28520));
    LocalMux I__4636 (
            .O(N__28541),
            .I(N__28520));
    Span4Mux_v I__4635 (
            .O(N__28538),
            .I(N__28511));
    Span4Mux_v I__4634 (
            .O(N__28533),
            .I(N__28511));
    Span4Mux_h I__4633 (
            .O(N__28528),
            .I(N__28511));
    Span4Mux_h I__4632 (
            .O(N__28525),
            .I(N__28511));
    Sp12to4 I__4631 (
            .O(N__28520),
            .I(N__28508));
    Span4Mux_h I__4630 (
            .O(N__28511),
            .I(N__28505));
    Span12Mux_v I__4629 (
            .O(N__28508),
            .I(N__28502));
    Span4Mux_h I__4628 (
            .O(N__28505),
            .I(N__28499));
    Odrv12 I__4627 (
            .O(N__28502),
            .I(iac_raw_buf_N_774));
    Odrv4 I__4626 (
            .O(N__28499),
            .I(iac_raw_buf_N_774));
    InMux I__4625 (
            .O(N__28494),
            .I(N__28491));
    LocalMux I__4624 (
            .O(N__28491),
            .I(n21334));
    InMux I__4623 (
            .O(N__28488),
            .I(N__28485));
    LocalMux I__4622 (
            .O(N__28485),
            .I(n22512));
    InMux I__4621 (
            .O(N__28482),
            .I(N__28478));
    InMux I__4620 (
            .O(N__28481),
            .I(N__28475));
    LocalMux I__4619 (
            .O(N__28478),
            .I(N__28472));
    LocalMux I__4618 (
            .O(N__28475),
            .I(data_idxvec_15));
    Odrv4 I__4617 (
            .O(N__28472),
            .I(data_idxvec_15));
    InMux I__4616 (
            .O(N__28467),
            .I(N__28464));
    LocalMux I__4615 (
            .O(N__28464),
            .I(N__28461));
    Span4Mux_h I__4614 (
            .O(N__28461),
            .I(N__28458));
    Span4Mux_h I__4613 (
            .O(N__28458),
            .I(N__28455));
    Sp12to4 I__4612 (
            .O(N__28455),
            .I(N__28452));
    Span12Mux_v I__4611 (
            .O(N__28452),
            .I(N__28449));
    Odrv12 I__4610 (
            .O(N__28449),
            .I(buf_data_iac_23));
    CascadeMux I__4609 (
            .O(N__28446),
            .I(n26_adj_1659_cascade_));
    CascadeMux I__4608 (
            .O(N__28443),
            .I(n21324_cascade_));
    InMux I__4607 (
            .O(N__28440),
            .I(N__28437));
    LocalMux I__4606 (
            .O(N__28437),
            .I(N__28434));
    Span4Mux_h I__4605 (
            .O(N__28434),
            .I(N__28429));
    InMux I__4604 (
            .O(N__28433),
            .I(N__28426));
    CascadeMux I__4603 (
            .O(N__28432),
            .I(N__28423));
    Span4Mux_h I__4602 (
            .O(N__28429),
            .I(N__28418));
    LocalMux I__4601 (
            .O(N__28426),
            .I(N__28418));
    InMux I__4600 (
            .O(N__28423),
            .I(N__28415));
    Span4Mux_h I__4599 (
            .O(N__28418),
            .I(N__28412));
    LocalMux I__4598 (
            .O(N__28415),
            .I(buf_adcdata_vac_15));
    Odrv4 I__4597 (
            .O(N__28412),
            .I(buf_adcdata_vac_15));
    InMux I__4596 (
            .O(N__28407),
            .I(N__28404));
    LocalMux I__4595 (
            .O(N__28404),
            .I(N__28400));
    InMux I__4594 (
            .O(N__28403),
            .I(N__28397));
    Span4Mux_v I__4593 (
            .O(N__28400),
            .I(N__28392));
    LocalMux I__4592 (
            .O(N__28397),
            .I(N__28392));
    Odrv4 I__4591 (
            .O(N__28392),
            .I(buf_adcdata_vdc_15));
    InMux I__4590 (
            .O(N__28389),
            .I(N__28386));
    LocalMux I__4589 (
            .O(N__28386),
            .I(N__28383));
    Span4Mux_h I__4588 (
            .O(N__28383),
            .I(N__28380));
    Odrv4 I__4587 (
            .O(N__28380),
            .I(n19_adj_1621));
    CascadeMux I__4586 (
            .O(N__28377),
            .I(N__28374));
    InMux I__4585 (
            .O(N__28374),
            .I(N__28371));
    LocalMux I__4584 (
            .O(N__28371),
            .I(N__28368));
    Odrv12 I__4583 (
            .O(N__28368),
            .I(n23_adj_1658));
    InMux I__4582 (
            .O(N__28365),
            .I(N__28362));
    LocalMux I__4581 (
            .O(N__28362),
            .I(n21323));
    InMux I__4580 (
            .O(N__28359),
            .I(N__28356));
    LocalMux I__4579 (
            .O(N__28356),
            .I(N__28353));
    Span4Mux_h I__4578 (
            .O(N__28353),
            .I(N__28350));
    Odrv4 I__4577 (
            .O(N__28350),
            .I(n19_adj_1652));
    CascadeMux I__4576 (
            .O(N__28347),
            .I(N__28344));
    InMux I__4575 (
            .O(N__28344),
            .I(N__28341));
    LocalMux I__4574 (
            .O(N__28341),
            .I(N__28338));
    Span4Mux_v I__4573 (
            .O(N__28338),
            .I(N__28334));
    CascadeMux I__4572 (
            .O(N__28337),
            .I(N__28331));
    Span4Mux_h I__4571 (
            .O(N__28334),
            .I(N__28328));
    InMux I__4570 (
            .O(N__28331),
            .I(N__28325));
    Odrv4 I__4569 (
            .O(N__28328),
            .I(buf_readRTD_1));
    LocalMux I__4568 (
            .O(N__28325),
            .I(buf_readRTD_1));
    InMux I__4567 (
            .O(N__28320),
            .I(N__28317));
    LocalMux I__4566 (
            .O(N__28317),
            .I(N__28314));
    Sp12to4 I__4565 (
            .O(N__28314),
            .I(N__28309));
    CascadeMux I__4564 (
            .O(N__28313),
            .I(N__28306));
    InMux I__4563 (
            .O(N__28312),
            .I(N__28303));
    Span12Mux_v I__4562 (
            .O(N__28309),
            .I(N__28300));
    InMux I__4561 (
            .O(N__28306),
            .I(N__28297));
    LocalMux I__4560 (
            .O(N__28303),
            .I(N__28292));
    Span12Mux_h I__4559 (
            .O(N__28300),
            .I(N__28292));
    LocalMux I__4558 (
            .O(N__28297),
            .I(buf_adcdata_vac_13));
    Odrv12 I__4557 (
            .O(N__28292),
            .I(buf_adcdata_vac_13));
    InMux I__4556 (
            .O(N__28287),
            .I(N__28284));
    LocalMux I__4555 (
            .O(N__28284),
            .I(N__28280));
    InMux I__4554 (
            .O(N__28283),
            .I(N__28277));
    Odrv12 I__4553 (
            .O(N__28280),
            .I(buf_readRTD_5));
    LocalMux I__4552 (
            .O(N__28277),
            .I(buf_readRTD_5));
    CascadeMux I__4551 (
            .O(N__28272),
            .I(n19_adj_1629_cascade_));
    InMux I__4550 (
            .O(N__28269),
            .I(N__28262));
    InMux I__4549 (
            .O(N__28268),
            .I(N__28257));
    InMux I__4548 (
            .O(N__28267),
            .I(N__28257));
    InMux I__4547 (
            .O(N__28266),
            .I(N__28251));
    InMux I__4546 (
            .O(N__28265),
            .I(N__28248));
    LocalMux I__4545 (
            .O(N__28262),
            .I(N__28241));
    LocalMux I__4544 (
            .O(N__28257),
            .I(N__28234));
    InMux I__4543 (
            .O(N__28256),
            .I(N__28227));
    InMux I__4542 (
            .O(N__28255),
            .I(N__28227));
    InMux I__4541 (
            .O(N__28254),
            .I(N__28227));
    LocalMux I__4540 (
            .O(N__28251),
            .I(N__28224));
    LocalMux I__4539 (
            .O(N__28248),
            .I(N__28221));
    InMux I__4538 (
            .O(N__28247),
            .I(N__28216));
    InMux I__4537 (
            .O(N__28246),
            .I(N__28216));
    InMux I__4536 (
            .O(N__28245),
            .I(N__28205));
    InMux I__4535 (
            .O(N__28244),
            .I(N__28205));
    Span4Mux_h I__4534 (
            .O(N__28241),
            .I(N__28202));
    InMux I__4533 (
            .O(N__28240),
            .I(N__28195));
    InMux I__4532 (
            .O(N__28239),
            .I(N__28195));
    InMux I__4531 (
            .O(N__28238),
            .I(N__28195));
    InMux I__4530 (
            .O(N__28237),
            .I(N__28192));
    Span4Mux_v I__4529 (
            .O(N__28234),
            .I(N__28180));
    LocalMux I__4528 (
            .O(N__28227),
            .I(N__28180));
    Span4Mux_h I__4527 (
            .O(N__28224),
            .I(N__28173));
    Span4Mux_v I__4526 (
            .O(N__28221),
            .I(N__28173));
    LocalMux I__4525 (
            .O(N__28216),
            .I(N__28173));
    InMux I__4524 (
            .O(N__28215),
            .I(N__28160));
    InMux I__4523 (
            .O(N__28214),
            .I(N__28160));
    InMux I__4522 (
            .O(N__28213),
            .I(N__28160));
    InMux I__4521 (
            .O(N__28212),
            .I(N__28160));
    InMux I__4520 (
            .O(N__28211),
            .I(N__28160));
    InMux I__4519 (
            .O(N__28210),
            .I(N__28160));
    LocalMux I__4518 (
            .O(N__28205),
            .I(N__28157));
    Span4Mux_v I__4517 (
            .O(N__28202),
            .I(N__28150));
    LocalMux I__4516 (
            .O(N__28195),
            .I(N__28150));
    LocalMux I__4515 (
            .O(N__28192),
            .I(N__28150));
    InMux I__4514 (
            .O(N__28191),
            .I(N__28145));
    InMux I__4513 (
            .O(N__28190),
            .I(N__28145));
    InMux I__4512 (
            .O(N__28189),
            .I(N__28138));
    InMux I__4511 (
            .O(N__28188),
            .I(N__28138));
    InMux I__4510 (
            .O(N__28187),
            .I(N__28138));
    InMux I__4509 (
            .O(N__28186),
            .I(N__28133));
    InMux I__4508 (
            .O(N__28185),
            .I(N__28133));
    Span4Mux_v I__4507 (
            .O(N__28180),
            .I(N__28127));
    Span4Mux_h I__4506 (
            .O(N__28173),
            .I(N__28122));
    LocalMux I__4505 (
            .O(N__28160),
            .I(N__28122));
    Span4Mux_v I__4504 (
            .O(N__28157),
            .I(N__28117));
    Span4Mux_h I__4503 (
            .O(N__28150),
            .I(N__28117));
    LocalMux I__4502 (
            .O(N__28145),
            .I(N__28112));
    LocalMux I__4501 (
            .O(N__28138),
            .I(N__28112));
    LocalMux I__4500 (
            .O(N__28133),
            .I(N__28109));
    InMux I__4499 (
            .O(N__28132),
            .I(N__28102));
    InMux I__4498 (
            .O(N__28131),
            .I(N__28102));
    InMux I__4497 (
            .O(N__28130),
            .I(N__28102));
    Odrv4 I__4496 (
            .O(N__28127),
            .I(n12850));
    Odrv4 I__4495 (
            .O(N__28122),
            .I(n12850));
    Odrv4 I__4494 (
            .O(N__28117),
            .I(n12850));
    Odrv12 I__4493 (
            .O(N__28112),
            .I(n12850));
    Odrv4 I__4492 (
            .O(N__28109),
            .I(n12850));
    LocalMux I__4491 (
            .O(N__28102),
            .I(n12850));
    InMux I__4490 (
            .O(N__28089),
            .I(N__28085));
    InMux I__4489 (
            .O(N__28088),
            .I(N__28082));
    LocalMux I__4488 (
            .O(N__28085),
            .I(N__28079));
    LocalMux I__4487 (
            .O(N__28082),
            .I(N__28075));
    Span4Mux_v I__4486 (
            .O(N__28079),
            .I(N__28072));
    InMux I__4485 (
            .O(N__28078),
            .I(N__28069));
    Odrv12 I__4484 (
            .O(N__28075),
            .I(cmd_rdadctmp_21_adj_1471));
    Odrv4 I__4483 (
            .O(N__28072),
            .I(cmd_rdadctmp_21_adj_1471));
    LocalMux I__4482 (
            .O(N__28069),
            .I(cmd_rdadctmp_21_adj_1471));
    CascadeMux I__4481 (
            .O(N__28062),
            .I(N__28059));
    InMux I__4480 (
            .O(N__28059),
            .I(N__28056));
    LocalMux I__4479 (
            .O(N__28056),
            .I(N__28053));
    Odrv4 I__4478 (
            .O(N__28053),
            .I(n8));
    InMux I__4477 (
            .O(N__28050),
            .I(N__28047));
    LocalMux I__4476 (
            .O(N__28047),
            .I(N__28043));
    InMux I__4475 (
            .O(N__28046),
            .I(N__28040));
    Span4Mux_v I__4474 (
            .O(N__28043),
            .I(N__28035));
    LocalMux I__4473 (
            .O(N__28040),
            .I(N__28035));
    Span4Mux_v I__4472 (
            .O(N__28035),
            .I(N__28031));
    InMux I__4471 (
            .O(N__28034),
            .I(N__28028));
    Odrv4 I__4470 (
            .O(N__28031),
            .I(n10695));
    LocalMux I__4469 (
            .O(N__28028),
            .I(n10695));
    InMux I__4468 (
            .O(N__28023),
            .I(N__28020));
    LocalMux I__4467 (
            .O(N__28020),
            .I(N__28016));
    CascadeMux I__4466 (
            .O(N__28019),
            .I(N__28013));
    Span4Mux_v I__4465 (
            .O(N__28016),
            .I(N__28010));
    InMux I__4464 (
            .O(N__28013),
            .I(N__28007));
    Odrv4 I__4463 (
            .O(N__28010),
            .I(buf_adcdata_vdc_12));
    LocalMux I__4462 (
            .O(N__28007),
            .I(buf_adcdata_vdc_12));
    InMux I__4461 (
            .O(N__28002),
            .I(N__27992));
    InMux I__4460 (
            .O(N__28001),
            .I(N__27992));
    InMux I__4459 (
            .O(N__28000),
            .I(N__27985));
    InMux I__4458 (
            .O(N__27999),
            .I(N__27982));
    InMux I__4457 (
            .O(N__27998),
            .I(N__27968));
    InMux I__4456 (
            .O(N__27997),
            .I(N__27968));
    LocalMux I__4455 (
            .O(N__27992),
            .I(N__27961));
    InMux I__4454 (
            .O(N__27991),
            .I(N__27952));
    InMux I__4453 (
            .O(N__27990),
            .I(N__27952));
    InMux I__4452 (
            .O(N__27989),
            .I(N__27952));
    InMux I__4451 (
            .O(N__27988),
            .I(N__27952));
    LocalMux I__4450 (
            .O(N__27985),
            .I(N__27947));
    LocalMux I__4449 (
            .O(N__27982),
            .I(N__27947));
    InMux I__4448 (
            .O(N__27981),
            .I(N__27940));
    InMux I__4447 (
            .O(N__27980),
            .I(N__27940));
    InMux I__4446 (
            .O(N__27979),
            .I(N__27940));
    InMux I__4445 (
            .O(N__27978),
            .I(N__27937));
    InMux I__4444 (
            .O(N__27977),
            .I(N__27928));
    InMux I__4443 (
            .O(N__27976),
            .I(N__27928));
    InMux I__4442 (
            .O(N__27975),
            .I(N__27928));
    InMux I__4441 (
            .O(N__27974),
            .I(N__27928));
    InMux I__4440 (
            .O(N__27973),
            .I(N__27925));
    LocalMux I__4439 (
            .O(N__27968),
            .I(N__27922));
    InMux I__4438 (
            .O(N__27967),
            .I(N__27917));
    InMux I__4437 (
            .O(N__27966),
            .I(N__27917));
    InMux I__4436 (
            .O(N__27965),
            .I(N__27914));
    CascadeMux I__4435 (
            .O(N__27964),
            .I(N__27911));
    Span4Mux_v I__4434 (
            .O(N__27961),
            .I(N__27906));
    LocalMux I__4433 (
            .O(N__27952),
            .I(N__27906));
    Span4Mux_v I__4432 (
            .O(N__27947),
            .I(N__27899));
    LocalMux I__4431 (
            .O(N__27940),
            .I(N__27899));
    LocalMux I__4430 (
            .O(N__27937),
            .I(N__27899));
    LocalMux I__4429 (
            .O(N__27928),
            .I(N__27894));
    LocalMux I__4428 (
            .O(N__27925),
            .I(N__27894));
    Span4Mux_v I__4427 (
            .O(N__27922),
            .I(N__27887));
    LocalMux I__4426 (
            .O(N__27917),
            .I(N__27887));
    LocalMux I__4425 (
            .O(N__27914),
            .I(N__27887));
    InMux I__4424 (
            .O(N__27911),
            .I(N__27884));
    Span4Mux_v I__4423 (
            .O(N__27906),
            .I(N__27880));
    Span4Mux_h I__4422 (
            .O(N__27899),
            .I(N__27877));
    Span4Mux_v I__4421 (
            .O(N__27894),
            .I(N__27870));
    Span4Mux_h I__4420 (
            .O(N__27887),
            .I(N__27870));
    LocalMux I__4419 (
            .O(N__27884),
            .I(N__27870));
    InMux I__4418 (
            .O(N__27883),
            .I(N__27867));
    Odrv4 I__4417 (
            .O(N__27880),
            .I(n21076));
    Odrv4 I__4416 (
            .O(N__27877),
            .I(n21076));
    Odrv4 I__4415 (
            .O(N__27870),
            .I(n21076));
    LocalMux I__4414 (
            .O(N__27867),
            .I(n21076));
    CascadeMux I__4413 (
            .O(N__27858),
            .I(N__27852));
    CascadeMux I__4412 (
            .O(N__27857),
            .I(N__27844));
    CascadeMux I__4411 (
            .O(N__27856),
            .I(N__27836));
    CascadeMux I__4410 (
            .O(N__27855),
            .I(N__27828));
    InMux I__4409 (
            .O(N__27852),
            .I(N__27817));
    InMux I__4408 (
            .O(N__27851),
            .I(N__27812));
    InMux I__4407 (
            .O(N__27850),
            .I(N__27812));
    InMux I__4406 (
            .O(N__27849),
            .I(N__27807));
    InMux I__4405 (
            .O(N__27848),
            .I(N__27807));
    CascadeMux I__4404 (
            .O(N__27847),
            .I(N__27797));
    InMux I__4403 (
            .O(N__27844),
            .I(N__27787));
    InMux I__4402 (
            .O(N__27843),
            .I(N__27784));
    InMux I__4401 (
            .O(N__27842),
            .I(N__27779));
    InMux I__4400 (
            .O(N__27841),
            .I(N__27779));
    InMux I__4399 (
            .O(N__27840),
            .I(N__27773));
    InMux I__4398 (
            .O(N__27839),
            .I(N__27773));
    InMux I__4397 (
            .O(N__27836),
            .I(N__27760));
    InMux I__4396 (
            .O(N__27835),
            .I(N__27760));
    InMux I__4395 (
            .O(N__27834),
            .I(N__27760));
    InMux I__4394 (
            .O(N__27833),
            .I(N__27760));
    InMux I__4393 (
            .O(N__27832),
            .I(N__27760));
    InMux I__4392 (
            .O(N__27831),
            .I(N__27760));
    InMux I__4391 (
            .O(N__27828),
            .I(N__27752));
    InMux I__4390 (
            .O(N__27827),
            .I(N__27747));
    InMux I__4389 (
            .O(N__27826),
            .I(N__27747));
    InMux I__4388 (
            .O(N__27825),
            .I(N__27742));
    InMux I__4387 (
            .O(N__27824),
            .I(N__27742));
    InMux I__4386 (
            .O(N__27823),
            .I(N__27733));
    InMux I__4385 (
            .O(N__27822),
            .I(N__27733));
    InMux I__4384 (
            .O(N__27821),
            .I(N__27733));
    InMux I__4383 (
            .O(N__27820),
            .I(N__27733));
    LocalMux I__4382 (
            .O(N__27817),
            .I(N__27726));
    LocalMux I__4381 (
            .O(N__27812),
            .I(N__27726));
    LocalMux I__4380 (
            .O(N__27807),
            .I(N__27726));
    InMux I__4379 (
            .O(N__27806),
            .I(N__27708));
    InMux I__4378 (
            .O(N__27805),
            .I(N__27708));
    InMux I__4377 (
            .O(N__27804),
            .I(N__27708));
    InMux I__4376 (
            .O(N__27803),
            .I(N__27708));
    InMux I__4375 (
            .O(N__27802),
            .I(N__27708));
    InMux I__4374 (
            .O(N__27801),
            .I(N__27708));
    InMux I__4373 (
            .O(N__27800),
            .I(N__27705));
    InMux I__4372 (
            .O(N__27797),
            .I(N__27700));
    InMux I__4371 (
            .O(N__27796),
            .I(N__27700));
    InMux I__4370 (
            .O(N__27795),
            .I(N__27687));
    InMux I__4369 (
            .O(N__27794),
            .I(N__27687));
    InMux I__4368 (
            .O(N__27793),
            .I(N__27687));
    InMux I__4367 (
            .O(N__27792),
            .I(N__27687));
    InMux I__4366 (
            .O(N__27791),
            .I(N__27687));
    InMux I__4365 (
            .O(N__27790),
            .I(N__27687));
    LocalMux I__4364 (
            .O(N__27787),
            .I(N__27684));
    LocalMux I__4363 (
            .O(N__27784),
            .I(N__27679));
    LocalMux I__4362 (
            .O(N__27779),
            .I(N__27679));
    InMux I__4361 (
            .O(N__27778),
            .I(N__27676));
    LocalMux I__4360 (
            .O(N__27773),
            .I(N__27671));
    LocalMux I__4359 (
            .O(N__27760),
            .I(N__27671));
    CascadeMux I__4358 (
            .O(N__27759),
            .I(N__27665));
    CascadeMux I__4357 (
            .O(N__27758),
            .I(N__27662));
    CascadeMux I__4356 (
            .O(N__27757),
            .I(N__27659));
    CascadeMux I__4355 (
            .O(N__27756),
            .I(N__27652));
    CascadeMux I__4354 (
            .O(N__27755),
            .I(N__27647));
    LocalMux I__4353 (
            .O(N__27752),
            .I(N__27639));
    LocalMux I__4352 (
            .O(N__27747),
            .I(N__27639));
    LocalMux I__4351 (
            .O(N__27742),
            .I(N__27632));
    LocalMux I__4350 (
            .O(N__27733),
            .I(N__27632));
    Span4Mux_v I__4349 (
            .O(N__27726),
            .I(N__27632));
    InMux I__4348 (
            .O(N__27725),
            .I(N__27621));
    InMux I__4347 (
            .O(N__27724),
            .I(N__27621));
    InMux I__4346 (
            .O(N__27723),
            .I(N__27621));
    InMux I__4345 (
            .O(N__27722),
            .I(N__27616));
    InMux I__4344 (
            .O(N__27721),
            .I(N__27616));
    LocalMux I__4343 (
            .O(N__27708),
            .I(N__27613));
    LocalMux I__4342 (
            .O(N__27705),
            .I(N__27610));
    LocalMux I__4341 (
            .O(N__27700),
            .I(N__27601));
    LocalMux I__4340 (
            .O(N__27687),
            .I(N__27601));
    Span4Mux_h I__4339 (
            .O(N__27684),
            .I(N__27601));
    Span4Mux_v I__4338 (
            .O(N__27679),
            .I(N__27601));
    LocalMux I__4337 (
            .O(N__27676),
            .I(N__27596));
    Span4Mux_v I__4336 (
            .O(N__27671),
            .I(N__27596));
    InMux I__4335 (
            .O(N__27670),
            .I(N__27589));
    InMux I__4334 (
            .O(N__27669),
            .I(N__27589));
    InMux I__4333 (
            .O(N__27668),
            .I(N__27589));
    InMux I__4332 (
            .O(N__27665),
            .I(N__27574));
    InMux I__4331 (
            .O(N__27662),
            .I(N__27574));
    InMux I__4330 (
            .O(N__27659),
            .I(N__27574));
    InMux I__4329 (
            .O(N__27658),
            .I(N__27574));
    InMux I__4328 (
            .O(N__27657),
            .I(N__27574));
    InMux I__4327 (
            .O(N__27656),
            .I(N__27574));
    InMux I__4326 (
            .O(N__27655),
            .I(N__27574));
    InMux I__4325 (
            .O(N__27652),
            .I(N__27571));
    InMux I__4324 (
            .O(N__27651),
            .I(N__27566));
    InMux I__4323 (
            .O(N__27650),
            .I(N__27566));
    InMux I__4322 (
            .O(N__27647),
            .I(N__27557));
    InMux I__4321 (
            .O(N__27646),
            .I(N__27557));
    InMux I__4320 (
            .O(N__27645),
            .I(N__27557));
    InMux I__4319 (
            .O(N__27644),
            .I(N__27557));
    Span4Mux_v I__4318 (
            .O(N__27639),
            .I(N__27552));
    Span4Mux_v I__4317 (
            .O(N__27632),
            .I(N__27552));
    InMux I__4316 (
            .O(N__27631),
            .I(N__27543));
    InMux I__4315 (
            .O(N__27630),
            .I(N__27543));
    InMux I__4314 (
            .O(N__27629),
            .I(N__27543));
    InMux I__4313 (
            .O(N__27628),
            .I(N__27543));
    LocalMux I__4312 (
            .O(N__27621),
            .I(N__27526));
    LocalMux I__4311 (
            .O(N__27616),
            .I(N__27526));
    Span4Mux_v I__4310 (
            .O(N__27613),
            .I(N__27526));
    Span4Mux_v I__4309 (
            .O(N__27610),
            .I(N__27526));
    Span4Mux_h I__4308 (
            .O(N__27601),
            .I(N__27526));
    Span4Mux_h I__4307 (
            .O(N__27596),
            .I(N__27526));
    LocalMux I__4306 (
            .O(N__27589),
            .I(N__27526));
    LocalMux I__4305 (
            .O(N__27574),
            .I(N__27526));
    LocalMux I__4304 (
            .O(N__27571),
            .I(adc_state_0_adj_1460));
    LocalMux I__4303 (
            .O(N__27566),
            .I(adc_state_0_adj_1460));
    LocalMux I__4302 (
            .O(N__27557),
            .I(adc_state_0_adj_1460));
    Odrv4 I__4301 (
            .O(N__27552),
            .I(adc_state_0_adj_1460));
    LocalMux I__4300 (
            .O(N__27543),
            .I(adc_state_0_adj_1460));
    Odrv4 I__4299 (
            .O(N__27526),
            .I(adc_state_0_adj_1460));
    CascadeMux I__4298 (
            .O(N__27513),
            .I(N__27509));
    InMux I__4297 (
            .O(N__27512),
            .I(N__27504));
    InMux I__4296 (
            .O(N__27509),
            .I(N__27504));
    LocalMux I__4295 (
            .O(N__27504),
            .I(N__27501));
    Span4Mux_v I__4294 (
            .O(N__27501),
            .I(N__27497));
    InMux I__4293 (
            .O(N__27500),
            .I(N__27494));
    Span4Mux_v I__4292 (
            .O(N__27497),
            .I(N__27489));
    LocalMux I__4291 (
            .O(N__27494),
            .I(N__27489));
    Odrv4 I__4290 (
            .O(N__27489),
            .I(cmd_rdadctmp_20_adj_1472));
    InMux I__4289 (
            .O(N__27486),
            .I(N__27483));
    LocalMux I__4288 (
            .O(N__27483),
            .I(N__27478));
    InMux I__4287 (
            .O(N__27482),
            .I(N__27473));
    InMux I__4286 (
            .O(N__27481),
            .I(N__27473));
    Span12Mux_v I__4285 (
            .O(N__27478),
            .I(N__27470));
    LocalMux I__4284 (
            .O(N__27473),
            .I(buf_adcdata_vac_12));
    Odrv12 I__4283 (
            .O(N__27470),
            .I(buf_adcdata_vac_12));
    CascadeMux I__4282 (
            .O(N__27465),
            .I(N__27462));
    InMux I__4281 (
            .O(N__27462),
            .I(N__27459));
    LocalMux I__4280 (
            .O(N__27459),
            .I(N__27455));
    InMux I__4279 (
            .O(N__27458),
            .I(N__27452));
    Span4Mux_v I__4278 (
            .O(N__27455),
            .I(N__27449));
    LocalMux I__4277 (
            .O(N__27452),
            .I(N__27446));
    Span4Mux_v I__4276 (
            .O(N__27449),
            .I(N__27442));
    Span4Mux_v I__4275 (
            .O(N__27446),
            .I(N__27439));
    InMux I__4274 (
            .O(N__27445),
            .I(N__27436));
    Odrv4 I__4273 (
            .O(N__27442),
            .I(cmd_rdadctmp_19_adj_1473));
    Odrv4 I__4272 (
            .O(N__27439),
            .I(cmd_rdadctmp_19_adj_1473));
    LocalMux I__4271 (
            .O(N__27436),
            .I(cmd_rdadctmp_19_adj_1473));
    InMux I__4270 (
            .O(N__27429),
            .I(N__27426));
    LocalMux I__4269 (
            .O(N__27426),
            .I(N__27422));
    InMux I__4268 (
            .O(N__27425),
            .I(N__27418));
    Span4Mux_v I__4267 (
            .O(N__27422),
            .I(N__27415));
    CascadeMux I__4266 (
            .O(N__27421),
            .I(N__27412));
    LocalMux I__4265 (
            .O(N__27418),
            .I(N__27409));
    Sp12to4 I__4264 (
            .O(N__27415),
            .I(N__27406));
    InMux I__4263 (
            .O(N__27412),
            .I(N__27403));
    Span4Mux_h I__4262 (
            .O(N__27409),
            .I(N__27400));
    Span12Mux_h I__4261 (
            .O(N__27406),
            .I(N__27397));
    LocalMux I__4260 (
            .O(N__27403),
            .I(buf_adcdata_vac_21));
    Odrv4 I__4259 (
            .O(N__27400),
            .I(buf_adcdata_vac_21));
    Odrv12 I__4258 (
            .O(N__27397),
            .I(buf_adcdata_vac_21));
    IoInMux I__4257 (
            .O(N__27390),
            .I(N__27387));
    LocalMux I__4256 (
            .O(N__27387),
            .I(N__27384));
    IoSpan4Mux I__4255 (
            .O(N__27384),
            .I(N__27380));
    InMux I__4254 (
            .O(N__27383),
            .I(N__27377));
    Sp12to4 I__4253 (
            .O(N__27380),
            .I(N__27374));
    LocalMux I__4252 (
            .O(N__27377),
            .I(N__27370));
    Span12Mux_h I__4251 (
            .O(N__27374),
            .I(N__27367));
    InMux I__4250 (
            .O(N__27373),
            .I(N__27364));
    Span4Mux_v I__4249 (
            .O(N__27370),
            .I(N__27361));
    Odrv12 I__4248 (
            .O(N__27367),
            .I(VAC_OSR1));
    LocalMux I__4247 (
            .O(N__27364),
            .I(VAC_OSR1));
    Odrv4 I__4246 (
            .O(N__27361),
            .I(VAC_OSR1));
    InMux I__4245 (
            .O(N__27354),
            .I(N__27351));
    LocalMux I__4244 (
            .O(N__27351),
            .I(N__27347));
    CascadeMux I__4243 (
            .O(N__27350),
            .I(N__27344));
    Span4Mux_v I__4242 (
            .O(N__27347),
            .I(N__27341));
    InMux I__4241 (
            .O(N__27344),
            .I(N__27338));
    Odrv4 I__4240 (
            .O(N__27341),
            .I(buf_adcdata_vdc_10));
    LocalMux I__4239 (
            .O(N__27338),
            .I(buf_adcdata_vdc_10));
    InMux I__4238 (
            .O(N__27333),
            .I(N__27330));
    LocalMux I__4237 (
            .O(N__27330),
            .I(N__27326));
    InMux I__4236 (
            .O(N__27329),
            .I(N__27322));
    Span4Mux_v I__4235 (
            .O(N__27326),
            .I(N__27319));
    CascadeMux I__4234 (
            .O(N__27325),
            .I(N__27316));
    LocalMux I__4233 (
            .O(N__27322),
            .I(N__27313));
    Span4Mux_v I__4232 (
            .O(N__27319),
            .I(N__27310));
    InMux I__4231 (
            .O(N__27316),
            .I(N__27307));
    Span4Mux_h I__4230 (
            .O(N__27313),
            .I(N__27304));
    Sp12to4 I__4229 (
            .O(N__27310),
            .I(N__27301));
    LocalMux I__4228 (
            .O(N__27307),
            .I(buf_adcdata_vac_10));
    Odrv4 I__4227 (
            .O(N__27304),
            .I(buf_adcdata_vac_10));
    Odrv12 I__4226 (
            .O(N__27301),
            .I(buf_adcdata_vac_10));
    InMux I__4225 (
            .O(N__27294),
            .I(N__27290));
    CascadeMux I__4224 (
            .O(N__27293),
            .I(N__27287));
    LocalMux I__4223 (
            .O(N__27290),
            .I(N__27284));
    InMux I__4222 (
            .O(N__27287),
            .I(N__27281));
    Span4Mux_v I__4221 (
            .O(N__27284),
            .I(N__27276));
    LocalMux I__4220 (
            .O(N__27281),
            .I(N__27276));
    Odrv4 I__4219 (
            .O(N__27276),
            .I(buf_adcdata_vdc_0));
    InMux I__4218 (
            .O(N__27273),
            .I(N__27269));
    InMux I__4217 (
            .O(N__27272),
            .I(N__27266));
    LocalMux I__4216 (
            .O(N__27269),
            .I(N__27263));
    LocalMux I__4215 (
            .O(N__27266),
            .I(N__27260));
    Span12Mux_s11_h I__4214 (
            .O(N__27263),
            .I(N__27256));
    Span4Mux_v I__4213 (
            .O(N__27260),
            .I(N__27253));
    InMux I__4212 (
            .O(N__27259),
            .I(N__27250));
    Span12Mux_h I__4211 (
            .O(N__27256),
            .I(N__27247));
    Span4Mux_h I__4210 (
            .O(N__27253),
            .I(N__27244));
    LocalMux I__4209 (
            .O(N__27250),
            .I(buf_adcdata_vac_0));
    Odrv12 I__4208 (
            .O(N__27247),
            .I(buf_adcdata_vac_0));
    Odrv4 I__4207 (
            .O(N__27244),
            .I(buf_adcdata_vac_0));
    InMux I__4206 (
            .O(N__27237),
            .I(N__27234));
    LocalMux I__4205 (
            .O(N__27234),
            .I(N__27231));
    Span4Mux_v I__4204 (
            .O(N__27231),
            .I(N__27227));
    InMux I__4203 (
            .O(N__27230),
            .I(N__27224));
    Sp12to4 I__4202 (
            .O(N__27227),
            .I(N__27220));
    LocalMux I__4201 (
            .O(N__27224),
            .I(N__27217));
    InMux I__4200 (
            .O(N__27223),
            .I(N__27214));
    Span12Mux_h I__4199 (
            .O(N__27220),
            .I(N__27211));
    Span4Mux_h I__4198 (
            .O(N__27217),
            .I(N__27208));
    LocalMux I__4197 (
            .O(N__27214),
            .I(buf_adcdata_iac_0));
    Odrv12 I__4196 (
            .O(N__27211),
            .I(buf_adcdata_iac_0));
    Odrv4 I__4195 (
            .O(N__27208),
            .I(buf_adcdata_iac_0));
    CascadeMux I__4194 (
            .O(N__27201),
            .I(n19_adj_1534_cascade_));
    InMux I__4193 (
            .O(N__27198),
            .I(N__27195));
    LocalMux I__4192 (
            .O(N__27195),
            .I(N__27192));
    Odrv12 I__4191 (
            .O(N__27192),
            .I(buf_control_7));
    IoInMux I__4190 (
            .O(N__27189),
            .I(N__27186));
    LocalMux I__4189 (
            .O(N__27186),
            .I(N__27183));
    Span4Mux_s3_v I__4188 (
            .O(N__27183),
            .I(N__27180));
    Sp12to4 I__4187 (
            .O(N__27180),
            .I(N__27176));
    CascadeMux I__4186 (
            .O(N__27179),
            .I(N__27173));
    Span12Mux_h I__4185 (
            .O(N__27176),
            .I(N__27170));
    InMux I__4184 (
            .O(N__27173),
            .I(N__27167));
    Odrv12 I__4183 (
            .O(N__27170),
            .I(DDS_SCK1));
    LocalMux I__4182 (
            .O(N__27167),
            .I(DDS_SCK1));
    CascadeMux I__4181 (
            .O(N__27162),
            .I(N__27159));
    InMux I__4180 (
            .O(N__27159),
            .I(N__27156));
    LocalMux I__4179 (
            .O(N__27156),
            .I(N__27153));
    Span4Mux_h I__4178 (
            .O(N__27153),
            .I(N__27150));
    Span4Mux_h I__4177 (
            .O(N__27150),
            .I(N__27146));
    InMux I__4176 (
            .O(N__27149),
            .I(N__27143));
    Odrv4 I__4175 (
            .O(N__27146),
            .I(buf_readRTD_15));
    LocalMux I__4174 (
            .O(N__27143),
            .I(buf_readRTD_15));
    CascadeMux I__4173 (
            .O(N__27138),
            .I(N__27134));
    InMux I__4172 (
            .O(N__27137),
            .I(N__27131));
    InMux I__4171 (
            .O(N__27134),
            .I(N__27128));
    LocalMux I__4170 (
            .O(N__27131),
            .I(buf_adcdata_vdc_23));
    LocalMux I__4169 (
            .O(N__27128),
            .I(buf_adcdata_vdc_23));
    CascadeMux I__4168 (
            .O(N__27123),
            .I(n22593_cascade_));
    InMux I__4167 (
            .O(N__27120),
            .I(N__27117));
    LocalMux I__4166 (
            .O(N__27117),
            .I(N__27114));
    Span4Mux_h I__4165 (
            .O(N__27114),
            .I(N__27110));
    InMux I__4164 (
            .O(N__27113),
            .I(N__27107));
    Sp12to4 I__4163 (
            .O(N__27110),
            .I(N__27104));
    LocalMux I__4162 (
            .O(N__27107),
            .I(N__27101));
    Span12Mux_v I__4161 (
            .O(N__27104),
            .I(N__27097));
    Span4Mux_h I__4160 (
            .O(N__27101),
            .I(N__27094));
    InMux I__4159 (
            .O(N__27100),
            .I(N__27091));
    Span12Mux_h I__4158 (
            .O(N__27097),
            .I(N__27088));
    Span4Mux_h I__4157 (
            .O(N__27094),
            .I(N__27085));
    LocalMux I__4156 (
            .O(N__27091),
            .I(buf_adcdata_vac_23));
    Odrv12 I__4155 (
            .O(N__27088),
            .I(buf_adcdata_vac_23));
    Odrv4 I__4154 (
            .O(N__27085),
            .I(buf_adcdata_vac_23));
    CascadeMux I__4153 (
            .O(N__27078),
            .I(N__27074));
    CascadeMux I__4152 (
            .O(N__27077),
            .I(N__27071));
    InMux I__4151 (
            .O(N__27074),
            .I(N__27067));
    InMux I__4150 (
            .O(N__27071),
            .I(N__27064));
    CascadeMux I__4149 (
            .O(N__27070),
            .I(N__27061));
    LocalMux I__4148 (
            .O(N__27067),
            .I(N__27057));
    LocalMux I__4147 (
            .O(N__27064),
            .I(N__27054));
    InMux I__4146 (
            .O(N__27061),
            .I(N__27050));
    InMux I__4145 (
            .O(N__27060),
            .I(N__27047));
    Span4Mux_h I__4144 (
            .O(N__27057),
            .I(N__27044));
    Span4Mux_v I__4143 (
            .O(N__27054),
            .I(N__27041));
    InMux I__4142 (
            .O(N__27053),
            .I(N__27038));
    LocalMux I__4141 (
            .O(N__27050),
            .I(N__27033));
    LocalMux I__4140 (
            .O(N__27047),
            .I(N__27033));
    Odrv4 I__4139 (
            .O(N__27044),
            .I(buf_cfgRTD_6));
    Odrv4 I__4138 (
            .O(N__27041),
            .I(buf_cfgRTD_6));
    LocalMux I__4137 (
            .O(N__27038),
            .I(buf_cfgRTD_6));
    Odrv12 I__4136 (
            .O(N__27033),
            .I(buf_cfgRTD_6));
    CascadeMux I__4135 (
            .O(N__27024),
            .I(N__27021));
    InMux I__4134 (
            .O(N__27021),
            .I(N__27018));
    LocalMux I__4133 (
            .O(N__27018),
            .I(N__27011));
    InMux I__4132 (
            .O(N__27017),
            .I(N__27006));
    InMux I__4131 (
            .O(N__27016),
            .I(N__27006));
    InMux I__4130 (
            .O(N__27015),
            .I(N__27001));
    InMux I__4129 (
            .O(N__27014),
            .I(N__27001));
    Span4Mux_v I__4128 (
            .O(N__27011),
            .I(N__26998));
    LocalMux I__4127 (
            .O(N__27006),
            .I(N__26995));
    LocalMux I__4126 (
            .O(N__27001),
            .I(N__26992));
    Odrv4 I__4125 (
            .O(N__26998),
            .I(buf_cfgRTD_7));
    Odrv4 I__4124 (
            .O(N__26995),
            .I(buf_cfgRTD_7));
    Odrv4 I__4123 (
            .O(N__26992),
            .I(buf_cfgRTD_7));
    CascadeMux I__4122 (
            .O(N__26985),
            .I(N__26982));
    InMux I__4121 (
            .O(N__26982),
            .I(N__26979));
    LocalMux I__4120 (
            .O(N__26979),
            .I(n30_adj_1499));
    InMux I__4119 (
            .O(N__26976),
            .I(N__26972));
    InMux I__4118 (
            .O(N__26975),
            .I(N__26969));
    LocalMux I__4117 (
            .O(N__26972),
            .I(\ADC_VDC.avg_cnt_10 ));
    LocalMux I__4116 (
            .O(N__26969),
            .I(\ADC_VDC.avg_cnt_10 ));
    InMux I__4115 (
            .O(N__26964),
            .I(\ADC_VDC.n19886 ));
    InMux I__4114 (
            .O(N__26961),
            .I(\ADC_VDC.n19887 ));
    InMux I__4113 (
            .O(N__26958),
            .I(N__26954));
    InMux I__4112 (
            .O(N__26957),
            .I(N__26951));
    LocalMux I__4111 (
            .O(N__26954),
            .I(\ADC_VDC.avg_cnt_11 ));
    LocalMux I__4110 (
            .O(N__26951),
            .I(\ADC_VDC.avg_cnt_11 ));
    CEMux I__4109 (
            .O(N__26946),
            .I(N__26942));
    CEMux I__4108 (
            .O(N__26945),
            .I(N__26937));
    LocalMux I__4107 (
            .O(N__26942),
            .I(N__26934));
    CEMux I__4106 (
            .O(N__26941),
            .I(N__26931));
    CEMux I__4105 (
            .O(N__26940),
            .I(N__26926));
    LocalMux I__4104 (
            .O(N__26937),
            .I(N__26923));
    Span4Mux_v I__4103 (
            .O(N__26934),
            .I(N__26918));
    LocalMux I__4102 (
            .O(N__26931),
            .I(N__26918));
    CEMux I__4101 (
            .O(N__26930),
            .I(N__26915));
    CEMux I__4100 (
            .O(N__26929),
            .I(N__26912));
    LocalMux I__4099 (
            .O(N__26926),
            .I(N__26909));
    Span4Mux_v I__4098 (
            .O(N__26923),
            .I(N__26901));
    Span4Mux_v I__4097 (
            .O(N__26918),
            .I(N__26901));
    LocalMux I__4096 (
            .O(N__26915),
            .I(N__26901));
    LocalMux I__4095 (
            .O(N__26912),
            .I(N__26897));
    Span4Mux_v I__4094 (
            .O(N__26909),
            .I(N__26894));
    CEMux I__4093 (
            .O(N__26908),
            .I(N__26891));
    Span4Mux_v I__4092 (
            .O(N__26901),
            .I(N__26888));
    InMux I__4091 (
            .O(N__26900),
            .I(N__26885));
    Span4Mux_v I__4090 (
            .O(N__26897),
            .I(N__26880));
    Span4Mux_h I__4089 (
            .O(N__26894),
            .I(N__26880));
    LocalMux I__4088 (
            .O(N__26891),
            .I(N__26873));
    Span4Mux_h I__4087 (
            .O(N__26888),
            .I(N__26873));
    LocalMux I__4086 (
            .O(N__26885),
            .I(N__26873));
    Odrv4 I__4085 (
            .O(N__26880),
            .I(\ADC_VDC.n13463 ));
    Odrv4 I__4084 (
            .O(N__26873),
            .I(\ADC_VDC.n13463 ));
    SRMux I__4083 (
            .O(N__26868),
            .I(N__26865));
    LocalMux I__4082 (
            .O(N__26865),
            .I(N__26860));
    SRMux I__4081 (
            .O(N__26864),
            .I(N__26857));
    SRMux I__4080 (
            .O(N__26863),
            .I(N__26850));
    Span4Mux_h I__4079 (
            .O(N__26860),
            .I(N__26845));
    LocalMux I__4078 (
            .O(N__26857),
            .I(N__26845));
    SRMux I__4077 (
            .O(N__26856),
            .I(N__26842));
    SRMux I__4076 (
            .O(N__26855),
            .I(N__26839));
    SRMux I__4075 (
            .O(N__26854),
            .I(N__26836));
    SRMux I__4074 (
            .O(N__26853),
            .I(N__26833));
    LocalMux I__4073 (
            .O(N__26850),
            .I(N__26830));
    Span4Mux_v I__4072 (
            .O(N__26845),
            .I(N__26827));
    LocalMux I__4071 (
            .O(N__26842),
            .I(N__26824));
    LocalMux I__4070 (
            .O(N__26839),
            .I(N__26819));
    LocalMux I__4069 (
            .O(N__26836),
            .I(N__26819));
    LocalMux I__4068 (
            .O(N__26833),
            .I(N__26816));
    Span4Mux_v I__4067 (
            .O(N__26830),
            .I(N__26813));
    Span4Mux_h I__4066 (
            .O(N__26827),
            .I(N__26810));
    Span4Mux_v I__4065 (
            .O(N__26824),
            .I(N__26805));
    Span4Mux_v I__4064 (
            .O(N__26819),
            .I(N__26805));
    Odrv12 I__4063 (
            .O(N__26816),
            .I(\ADC_VDC.n15175 ));
    Odrv4 I__4062 (
            .O(N__26813),
            .I(\ADC_VDC.n15175 ));
    Odrv4 I__4061 (
            .O(N__26810),
            .I(\ADC_VDC.n15175 ));
    Odrv4 I__4060 (
            .O(N__26805),
            .I(\ADC_VDC.n15175 ));
    InMux I__4059 (
            .O(N__26796),
            .I(N__26793));
    LocalMux I__4058 (
            .O(N__26793),
            .I(N__26789));
    InMux I__4057 (
            .O(N__26792),
            .I(N__26786));
    Odrv4 I__4056 (
            .O(N__26789),
            .I(cmd_rdadcbuf_23));
    LocalMux I__4055 (
            .O(N__26786),
            .I(cmd_rdadcbuf_23));
    InMux I__4054 (
            .O(N__26781),
            .I(N__26778));
    LocalMux I__4053 (
            .O(N__26778),
            .I(N__26774));
    InMux I__4052 (
            .O(N__26777),
            .I(N__26771));
    Odrv4 I__4051 (
            .O(N__26774),
            .I(cmd_rdadcbuf_18));
    LocalMux I__4050 (
            .O(N__26771),
            .I(cmd_rdadcbuf_18));
    InMux I__4049 (
            .O(N__26766),
            .I(N__26763));
    LocalMux I__4048 (
            .O(N__26763),
            .I(N__26760));
    Span12Mux_v I__4047 (
            .O(N__26760),
            .I(N__26756));
    InMux I__4046 (
            .O(N__26759),
            .I(N__26753));
    Odrv12 I__4045 (
            .O(N__26756),
            .I(buf_adcdata_vdc_7));
    LocalMux I__4044 (
            .O(N__26753),
            .I(buf_adcdata_vdc_7));
    CascadeMux I__4043 (
            .O(N__26748),
            .I(n11891_cascade_));
    InMux I__4042 (
            .O(N__26745),
            .I(N__26742));
    LocalMux I__4041 (
            .O(N__26742),
            .I(N__26739));
    Span4Mux_h I__4040 (
            .O(N__26739),
            .I(N__26735));
    InMux I__4039 (
            .O(N__26738),
            .I(N__26732));
    Odrv4 I__4038 (
            .O(N__26735),
            .I(cmd_rdadcbuf_26));
    LocalMux I__4037 (
            .O(N__26732),
            .I(cmd_rdadcbuf_26));
    InMux I__4036 (
            .O(N__26727),
            .I(N__26724));
    LocalMux I__4035 (
            .O(N__26724),
            .I(N__26721));
    Span4Mux_v I__4034 (
            .O(N__26721),
            .I(N__26717));
    InMux I__4033 (
            .O(N__26720),
            .I(N__26714));
    Odrv4 I__4032 (
            .O(N__26717),
            .I(cmd_rdadcbuf_25));
    LocalMux I__4031 (
            .O(N__26714),
            .I(cmd_rdadcbuf_25));
    InMux I__4030 (
            .O(N__26709),
            .I(N__26706));
    LocalMux I__4029 (
            .O(N__26706),
            .I(N__26702));
    InMux I__4028 (
            .O(N__26705),
            .I(N__26699));
    Odrv12 I__4027 (
            .O(N__26702),
            .I(cmd_rdadcbuf_22));
    LocalMux I__4026 (
            .O(N__26699),
            .I(cmd_rdadcbuf_22));
    InMux I__4025 (
            .O(N__26694),
            .I(N__26691));
    LocalMux I__4024 (
            .O(N__26691),
            .I(N__26687));
    InMux I__4023 (
            .O(N__26690),
            .I(N__26684));
    Span4Mux_v I__4022 (
            .O(N__26687),
            .I(N__26681));
    LocalMux I__4021 (
            .O(N__26684),
            .I(\ADC_VDC.avg_cnt_1 ));
    Odrv4 I__4020 (
            .O(N__26681),
            .I(\ADC_VDC.avg_cnt_1 ));
    InMux I__4019 (
            .O(N__26676),
            .I(\ADC_VDC.n19877 ));
    CascadeMux I__4018 (
            .O(N__26673),
            .I(N__26670));
    InMux I__4017 (
            .O(N__26670),
            .I(N__26666));
    InMux I__4016 (
            .O(N__26669),
            .I(N__26663));
    LocalMux I__4015 (
            .O(N__26666),
            .I(N__26660));
    LocalMux I__4014 (
            .O(N__26663),
            .I(\ADC_VDC.avg_cnt_2 ));
    Odrv4 I__4013 (
            .O(N__26660),
            .I(\ADC_VDC.avg_cnt_2 ));
    InMux I__4012 (
            .O(N__26655),
            .I(\ADC_VDC.n19878 ));
    InMux I__4011 (
            .O(N__26652),
            .I(\ADC_VDC.n19879 ));
    InMux I__4010 (
            .O(N__26649),
            .I(N__26645));
    InMux I__4009 (
            .O(N__26648),
            .I(N__26642));
    LocalMux I__4008 (
            .O(N__26645),
            .I(N__26639));
    LocalMux I__4007 (
            .O(N__26642),
            .I(\ADC_VDC.avg_cnt_4 ));
    Odrv4 I__4006 (
            .O(N__26639),
            .I(\ADC_VDC.avg_cnt_4 ));
    InMux I__4005 (
            .O(N__26634),
            .I(\ADC_VDC.n19880 ));
    CascadeMux I__4004 (
            .O(N__26631),
            .I(N__26627));
    InMux I__4003 (
            .O(N__26630),
            .I(N__26624));
    InMux I__4002 (
            .O(N__26627),
            .I(N__26621));
    LocalMux I__4001 (
            .O(N__26624),
            .I(\ADC_VDC.avg_cnt_5 ));
    LocalMux I__4000 (
            .O(N__26621),
            .I(\ADC_VDC.avg_cnt_5 ));
    InMux I__3999 (
            .O(N__26616),
            .I(\ADC_VDC.n19881 ));
    InMux I__3998 (
            .O(N__26613),
            .I(\ADC_VDC.n19882 ));
    InMux I__3997 (
            .O(N__26610),
            .I(N__26606));
    InMux I__3996 (
            .O(N__26609),
            .I(N__26603));
    LocalMux I__3995 (
            .O(N__26606),
            .I(N__26600));
    LocalMux I__3994 (
            .O(N__26603),
            .I(\ADC_VDC.avg_cnt_7 ));
    Odrv4 I__3993 (
            .O(N__26600),
            .I(\ADC_VDC.avg_cnt_7 ));
    InMux I__3992 (
            .O(N__26595),
            .I(\ADC_VDC.n19883 ));
    InMux I__3991 (
            .O(N__26592),
            .I(bfn_10_7_0_));
    InMux I__3990 (
            .O(N__26589),
            .I(\ADC_VDC.n19885 ));
    CascadeMux I__3989 (
            .O(N__26586),
            .I(N__26581));
    InMux I__3988 (
            .O(N__26585),
            .I(N__26578));
    InMux I__3987 (
            .O(N__26584),
            .I(N__26575));
    InMux I__3986 (
            .O(N__26581),
            .I(N__26572));
    LocalMux I__3985 (
            .O(N__26578),
            .I(cmd_rdadctmp_30));
    LocalMux I__3984 (
            .O(N__26575),
            .I(cmd_rdadctmp_30));
    LocalMux I__3983 (
            .O(N__26572),
            .I(cmd_rdadctmp_30));
    InMux I__3982 (
            .O(N__26565),
            .I(N__26562));
    LocalMux I__3981 (
            .O(N__26562),
            .I(N__26559));
    Span4Mux_v I__3980 (
            .O(N__26559),
            .I(N__26556));
    Odrv4 I__3979 (
            .O(N__26556),
            .I(\ADC_VDC.n18780 ));
    CascadeMux I__3978 (
            .O(N__26553),
            .I(\ADC_VDC.n18783_cascade_ ));
    CEMux I__3977 (
            .O(N__26550),
            .I(N__26547));
    LocalMux I__3976 (
            .O(N__26547),
            .I(\ADC_VDC.n16_adj_1450 ));
    InMux I__3975 (
            .O(N__26544),
            .I(N__26541));
    LocalMux I__3974 (
            .O(N__26541),
            .I(\ADC_VDC.n18 ));
    CascadeMux I__3973 (
            .O(N__26538),
            .I(\ADC_VDC.n18_cascade_ ));
    InMux I__3972 (
            .O(N__26535),
            .I(N__26532));
    LocalMux I__3971 (
            .O(N__26532),
            .I(N__26529));
    Span4Mux_h I__3970 (
            .O(N__26529),
            .I(N__26526));
    Sp12to4 I__3969 (
            .O(N__26526),
            .I(N__26523));
    Span12Mux_v I__3968 (
            .O(N__26523),
            .I(N__26520));
    Odrv12 I__3967 (
            .O(N__26520),
            .I(THERMOSTAT));
    InMux I__3966 (
            .O(N__26517),
            .I(N__26513));
    InMux I__3965 (
            .O(N__26516),
            .I(N__26510));
    LocalMux I__3964 (
            .O(N__26513),
            .I(\ADC_VDC.avg_cnt_0 ));
    LocalMux I__3963 (
            .O(N__26510),
            .I(\ADC_VDC.avg_cnt_0 ));
    InMux I__3962 (
            .O(N__26505),
            .I(bfn_10_6_0_));
    IoInMux I__3961 (
            .O(N__26502),
            .I(N__26499));
    LocalMux I__3960 (
            .O(N__26499),
            .I(N__26496));
    IoSpan4Mux I__3959 (
            .O(N__26496),
            .I(N__26493));
    Span4Mux_s1_v I__3958 (
            .O(N__26493),
            .I(N__26490));
    Span4Mux_v I__3957 (
            .O(N__26490),
            .I(N__26487));
    Span4Mux_v I__3956 (
            .O(N__26487),
            .I(N__26482));
    InMux I__3955 (
            .O(N__26486),
            .I(N__26477));
    InMux I__3954 (
            .O(N__26485),
            .I(N__26477));
    Odrv4 I__3953 (
            .O(N__26482),
            .I(IAC_FLT1));
    LocalMux I__3952 (
            .O(N__26477),
            .I(IAC_FLT1));
    InMux I__3951 (
            .O(N__26472),
            .I(N__26469));
    LocalMux I__3950 (
            .O(N__26469),
            .I(N__26466));
    Span12Mux_v I__3949 (
            .O(N__26466),
            .I(N__26462));
    CascadeMux I__3948 (
            .O(N__26465),
            .I(N__26458));
    Span12Mux_h I__3947 (
            .O(N__26462),
            .I(N__26455));
    InMux I__3946 (
            .O(N__26461),
            .I(N__26450));
    InMux I__3945 (
            .O(N__26458),
            .I(N__26450));
    Odrv12 I__3944 (
            .O(N__26455),
            .I(buf_adcdata_iac_19));
    LocalMux I__3943 (
            .O(N__26450),
            .I(buf_adcdata_iac_19));
    CascadeMux I__3942 (
            .O(N__26445),
            .I(n22605_cascade_));
    InMux I__3941 (
            .O(N__26442),
            .I(N__26438));
    InMux I__3940 (
            .O(N__26441),
            .I(N__26435));
    LocalMux I__3939 (
            .O(N__26438),
            .I(N__26432));
    LocalMux I__3938 (
            .O(N__26435),
            .I(N__26426));
    Span4Mux_v I__3937 (
            .O(N__26432),
            .I(N__26426));
    InMux I__3936 (
            .O(N__26431),
            .I(N__26423));
    Odrv4 I__3935 (
            .O(N__26426),
            .I(buf_dds1_11));
    LocalMux I__3934 (
            .O(N__26423),
            .I(buf_dds1_11));
    InMux I__3933 (
            .O(N__26418),
            .I(N__26415));
    LocalMux I__3932 (
            .O(N__26415),
            .I(N__26412));
    Odrv12 I__3931 (
            .O(N__26412),
            .I(n22608));
    InMux I__3930 (
            .O(N__26409),
            .I(N__26405));
    CascadeMux I__3929 (
            .O(N__26408),
            .I(N__26402));
    LocalMux I__3928 (
            .O(N__26405),
            .I(N__26398));
    InMux I__3927 (
            .O(N__26402),
            .I(N__26395));
    InMux I__3926 (
            .O(N__26401),
            .I(N__26392));
    Odrv4 I__3925 (
            .O(N__26398),
            .I(cmd_rdadctmp_27));
    LocalMux I__3924 (
            .O(N__26395),
            .I(cmd_rdadctmp_27));
    LocalMux I__3923 (
            .O(N__26392),
            .I(cmd_rdadctmp_27));
    InMux I__3922 (
            .O(N__26385),
            .I(N__26380));
    InMux I__3921 (
            .O(N__26384),
            .I(N__26375));
    InMux I__3920 (
            .O(N__26383),
            .I(N__26375));
    LocalMux I__3919 (
            .O(N__26380),
            .I(cmd_rdadctmp_19));
    LocalMux I__3918 (
            .O(N__26375),
            .I(cmd_rdadctmp_19));
    CascadeMux I__3917 (
            .O(N__26370),
            .I(N__26366));
    InMux I__3916 (
            .O(N__26369),
            .I(N__26358));
    InMux I__3915 (
            .O(N__26366),
            .I(N__26358));
    InMux I__3914 (
            .O(N__26365),
            .I(N__26358));
    LocalMux I__3913 (
            .O(N__26358),
            .I(cmd_rdadctmp_24));
    CascadeMux I__3912 (
            .O(N__26355),
            .I(N__26351));
    CascadeMux I__3911 (
            .O(N__26354),
            .I(N__26348));
    InMux I__3910 (
            .O(N__26351),
            .I(N__26342));
    InMux I__3909 (
            .O(N__26348),
            .I(N__26342));
    CascadeMux I__3908 (
            .O(N__26347),
            .I(N__26339));
    LocalMux I__3907 (
            .O(N__26342),
            .I(N__26336));
    InMux I__3906 (
            .O(N__26339),
            .I(N__26333));
    Odrv4 I__3905 (
            .O(N__26336),
            .I(cmd_rdadctmp_22_adj_1470));
    LocalMux I__3904 (
            .O(N__26333),
            .I(cmd_rdadctmp_22_adj_1470));
    CascadeMux I__3903 (
            .O(N__26328),
            .I(N__26324));
    InMux I__3902 (
            .O(N__26327),
            .I(N__26316));
    InMux I__3901 (
            .O(N__26324),
            .I(N__26316));
    InMux I__3900 (
            .O(N__26323),
            .I(N__26316));
    LocalMux I__3899 (
            .O(N__26316),
            .I(cmd_rdadctmp_23_adj_1469));
    InMux I__3898 (
            .O(N__26313),
            .I(N__26310));
    LocalMux I__3897 (
            .O(N__26310),
            .I(N__26307));
    Span4Mux_v I__3896 (
            .O(N__26307),
            .I(N__26304));
    Odrv4 I__3895 (
            .O(N__26304),
            .I(n69));
    CascadeMux I__3894 (
            .O(N__26301),
            .I(N__26297));
    CascadeMux I__3893 (
            .O(N__26300),
            .I(N__26294));
    InMux I__3892 (
            .O(N__26297),
            .I(N__26291));
    InMux I__3891 (
            .O(N__26294),
            .I(N__26288));
    LocalMux I__3890 (
            .O(N__26291),
            .I(N__26285));
    LocalMux I__3889 (
            .O(N__26288),
            .I(N__26282));
    Span4Mux_v I__3888 (
            .O(N__26285),
            .I(N__26278));
    Span4Mux_v I__3887 (
            .O(N__26282),
            .I(N__26275));
    InMux I__3886 (
            .O(N__26281),
            .I(N__26272));
    Odrv4 I__3885 (
            .O(N__26278),
            .I(cmd_rdadctmp_15));
    Odrv4 I__3884 (
            .O(N__26275),
            .I(cmd_rdadctmp_15));
    LocalMux I__3883 (
            .O(N__26272),
            .I(cmd_rdadctmp_15));
    InMux I__3882 (
            .O(N__26265),
            .I(N__26260));
    InMux I__3881 (
            .O(N__26264),
            .I(N__26255));
    InMux I__3880 (
            .O(N__26263),
            .I(N__26255));
    LocalMux I__3879 (
            .O(N__26260),
            .I(buf_dds1_2));
    LocalMux I__3878 (
            .O(N__26255),
            .I(buf_dds1_2));
    InMux I__3877 (
            .O(N__26250),
            .I(N__26247));
    LocalMux I__3876 (
            .O(N__26247),
            .I(N__26244));
    Span4Mux_v I__3875 (
            .O(N__26244),
            .I(N__26241));
    Odrv4 I__3874 (
            .O(N__26241),
            .I(n22476));
    InMux I__3873 (
            .O(N__26238),
            .I(N__26235));
    LocalMux I__3872 (
            .O(N__26235),
            .I(N__26231));
    CascadeMux I__3871 (
            .O(N__26234),
            .I(N__26228));
    Span4Mux_h I__3870 (
            .O(N__26231),
            .I(N__26225));
    InMux I__3869 (
            .O(N__26228),
            .I(N__26222));
    Sp12to4 I__3868 (
            .O(N__26225),
            .I(N__26216));
    LocalMux I__3867 (
            .O(N__26222),
            .I(N__26216));
    InMux I__3866 (
            .O(N__26221),
            .I(N__26213));
    Odrv12 I__3865 (
            .O(N__26216),
            .I(cmd_rdadctmp_16_adj_1476));
    LocalMux I__3864 (
            .O(N__26213),
            .I(cmd_rdadctmp_16_adj_1476));
    CascadeMux I__3863 (
            .O(N__26208),
            .I(N__26204));
    CascadeMux I__3862 (
            .O(N__26207),
            .I(N__26201));
    InMux I__3861 (
            .O(N__26204),
            .I(N__26198));
    InMux I__3860 (
            .O(N__26201),
            .I(N__26195));
    LocalMux I__3859 (
            .O(N__26198),
            .I(N__26189));
    LocalMux I__3858 (
            .O(N__26195),
            .I(N__26189));
    InMux I__3857 (
            .O(N__26194),
            .I(N__26186));
    Odrv12 I__3856 (
            .O(N__26189),
            .I(cmd_rdadctmp_25_adj_1467));
    LocalMux I__3855 (
            .O(N__26186),
            .I(cmd_rdadctmp_25_adj_1467));
    InMux I__3854 (
            .O(N__26181),
            .I(N__26178));
    LocalMux I__3853 (
            .O(N__26178),
            .I(N__26175));
    Span4Mux_h I__3852 (
            .O(N__26175),
            .I(N__26170));
    InMux I__3851 (
            .O(N__26174),
            .I(N__26165));
    InMux I__3850 (
            .O(N__26173),
            .I(N__26165));
    Odrv4 I__3849 (
            .O(N__26170),
            .I(cmd_rdadctmp_24_adj_1468));
    LocalMux I__3848 (
            .O(N__26165),
            .I(cmd_rdadctmp_24_adj_1468));
    CEMux I__3847 (
            .O(N__26160),
            .I(N__26157));
    LocalMux I__3846 (
            .O(N__26157),
            .I(N__26153));
    CEMux I__3845 (
            .O(N__26156),
            .I(N__26150));
    Span4Mux_v I__3844 (
            .O(N__26153),
            .I(N__26147));
    LocalMux I__3843 (
            .O(N__26150),
            .I(N__26142));
    Span4Mux_v I__3842 (
            .O(N__26147),
            .I(N__26142));
    Odrv4 I__3841 (
            .O(N__26142),
            .I(n12493));
    InMux I__3840 (
            .O(N__26139),
            .I(N__26136));
    LocalMux I__3839 (
            .O(N__26136),
            .I(N__26133));
    Span4Mux_h I__3838 (
            .O(N__26133),
            .I(N__26130));
    Odrv4 I__3837 (
            .O(N__26130),
            .I(n21705));
    CascadeMux I__3836 (
            .O(N__26127),
            .I(N__26123));
    CascadeMux I__3835 (
            .O(N__26126),
            .I(N__26119));
    InMux I__3834 (
            .O(N__26123),
            .I(N__26116));
    InMux I__3833 (
            .O(N__26122),
            .I(N__26113));
    InMux I__3832 (
            .O(N__26119),
            .I(N__26110));
    LocalMux I__3831 (
            .O(N__26116),
            .I(N__26107));
    LocalMux I__3830 (
            .O(N__26113),
            .I(cmd_rdadctmp_18_adj_1474));
    LocalMux I__3829 (
            .O(N__26110),
            .I(cmd_rdadctmp_18_adj_1474));
    Odrv12 I__3828 (
            .O(N__26107),
            .I(cmd_rdadctmp_18_adj_1474));
    IoInMux I__3827 (
            .O(N__26100),
            .I(N__26097));
    LocalMux I__3826 (
            .O(N__26097),
            .I(N__26094));
    IoSpan4Mux I__3825 (
            .O(N__26094),
            .I(N__26091));
    IoSpan4Mux I__3824 (
            .O(N__26091),
            .I(N__26087));
    InMux I__3823 (
            .O(N__26090),
            .I(N__26084));
    Sp12to4 I__3822 (
            .O(N__26087),
            .I(N__26081));
    LocalMux I__3821 (
            .O(N__26084),
            .I(N__26077));
    Span12Mux_s6_v I__3820 (
            .O(N__26081),
            .I(N__26074));
    InMux I__3819 (
            .O(N__26080),
            .I(N__26071));
    Span4Mux_v I__3818 (
            .O(N__26077),
            .I(N__26068));
    Odrv12 I__3817 (
            .O(N__26074),
            .I(IAC_OSR1));
    LocalMux I__3816 (
            .O(N__26071),
            .I(IAC_OSR1));
    Odrv4 I__3815 (
            .O(N__26068),
            .I(IAC_OSR1));
    CascadeMux I__3814 (
            .O(N__26061),
            .I(N__26057));
    InMux I__3813 (
            .O(N__26060),
            .I(N__26054));
    InMux I__3812 (
            .O(N__26057),
            .I(N__26051));
    LocalMux I__3811 (
            .O(N__26054),
            .I(N__26048));
    LocalMux I__3810 (
            .O(N__26051),
            .I(data_idxvec_11));
    Odrv4 I__3809 (
            .O(N__26048),
            .I(data_idxvec_11));
    CascadeMux I__3808 (
            .O(N__26043),
            .I(n26_adj_1678_cascade_));
    InMux I__3807 (
            .O(N__26040),
            .I(N__26037));
    LocalMux I__3806 (
            .O(N__26037),
            .I(n22509));
    InMux I__3805 (
            .O(N__26034),
            .I(bfn_9_12_0_));
    InMux I__3804 (
            .O(N__26031),
            .I(n19821));
    InMux I__3803 (
            .O(N__26028),
            .I(n19822));
    InMux I__3802 (
            .O(N__26025),
            .I(n19823));
    InMux I__3801 (
            .O(N__26022),
            .I(n19824));
    InMux I__3800 (
            .O(N__26019),
            .I(n19825));
    InMux I__3799 (
            .O(N__26016),
            .I(n19826));
    InMux I__3798 (
            .O(N__26013),
            .I(n19827));
    CascadeMux I__3797 (
            .O(N__26010),
            .I(N__26007));
    InMux I__3796 (
            .O(N__26007),
            .I(N__26004));
    LocalMux I__3795 (
            .O(N__26004),
            .I(N__26000));
    InMux I__3794 (
            .O(N__26003),
            .I(N__25997));
    Span4Mux_v I__3793 (
            .O(N__26000),
            .I(N__25993));
    LocalMux I__3792 (
            .O(N__25997),
            .I(N__25990));
    InMux I__3791 (
            .O(N__25996),
            .I(N__25987));
    Odrv4 I__3790 (
            .O(N__25993),
            .I(cmd_rdadctmp_27_adj_1465));
    Odrv4 I__3789 (
            .O(N__25990),
            .I(cmd_rdadctmp_27_adj_1465));
    LocalMux I__3788 (
            .O(N__25987),
            .I(cmd_rdadctmp_27_adj_1465));
    InMux I__3787 (
            .O(N__25980),
            .I(N__25977));
    LocalMux I__3786 (
            .O(N__25977),
            .I(N__25974));
    Span4Mux_h I__3785 (
            .O(N__25974),
            .I(N__25971));
    Span4Mux_v I__3784 (
            .O(N__25971),
            .I(N__25966));
    InMux I__3783 (
            .O(N__25970),
            .I(N__25963));
    InMux I__3782 (
            .O(N__25969),
            .I(N__25960));
    Sp12to4 I__3781 (
            .O(N__25966),
            .I(N__25957));
    LocalMux I__3780 (
            .O(N__25963),
            .I(N__25954));
    LocalMux I__3779 (
            .O(N__25960),
            .I(buf_adcdata_vac_19));
    Odrv12 I__3778 (
            .O(N__25957),
            .I(buf_adcdata_vac_19));
    Odrv12 I__3777 (
            .O(N__25954),
            .I(buf_adcdata_vac_19));
    CascadeMux I__3776 (
            .O(N__25947),
            .I(N__25943));
    InMux I__3775 (
            .O(N__25946),
            .I(N__25939));
    InMux I__3774 (
            .O(N__25943),
            .I(N__25934));
    InMux I__3773 (
            .O(N__25942),
            .I(N__25934));
    LocalMux I__3772 (
            .O(N__25939),
            .I(N__25929));
    LocalMux I__3771 (
            .O(N__25934),
            .I(N__25929));
    Span4Mux_v I__3770 (
            .O(N__25929),
            .I(N__25924));
    InMux I__3769 (
            .O(N__25928),
            .I(N__25919));
    InMux I__3768 (
            .O(N__25927),
            .I(N__25919));
    Odrv4 I__3767 (
            .O(N__25924),
            .I(buf_cfgRTD_3));
    LocalMux I__3766 (
            .O(N__25919),
            .I(buf_cfgRTD_3));
    CascadeMux I__3765 (
            .O(N__25914),
            .I(N__25911));
    InMux I__3764 (
            .O(N__25911),
            .I(N__25908));
    LocalMux I__3763 (
            .O(N__25908),
            .I(N__25904));
    InMux I__3762 (
            .O(N__25907),
            .I(N__25901));
    Odrv12 I__3761 (
            .O(N__25904),
            .I(buf_readRTD_11));
    LocalMux I__3760 (
            .O(N__25901),
            .I(buf_readRTD_11));
    InMux I__3759 (
            .O(N__25896),
            .I(N__25893));
    LocalMux I__3758 (
            .O(N__25893),
            .I(N__25890));
    Odrv12 I__3757 (
            .O(N__25890),
            .I(n22473));
    InMux I__3756 (
            .O(N__25887),
            .I(bfn_9_11_0_));
    InMux I__3755 (
            .O(N__25884),
            .I(n19813));
    InMux I__3754 (
            .O(N__25881),
            .I(n19814));
    InMux I__3753 (
            .O(N__25878),
            .I(n19815));
    InMux I__3752 (
            .O(N__25875),
            .I(n19816));
    InMux I__3751 (
            .O(N__25872),
            .I(n19817));
    InMux I__3750 (
            .O(N__25869),
            .I(n19818));
    InMux I__3749 (
            .O(N__25866),
            .I(n19819));
    InMux I__3748 (
            .O(N__25863),
            .I(N__25858));
    InMux I__3747 (
            .O(N__25862),
            .I(N__25855));
    InMux I__3746 (
            .O(N__25861),
            .I(N__25852));
    LocalMux I__3745 (
            .O(N__25858),
            .I(cmd_rdadcbuf_34));
    LocalMux I__3744 (
            .O(N__25855),
            .I(cmd_rdadcbuf_34));
    LocalMux I__3743 (
            .O(N__25852),
            .I(cmd_rdadcbuf_34));
    CascadeMux I__3742 (
            .O(N__25845),
            .I(\ADC_VDC.n18780_cascade_ ));
    CascadeMux I__3741 (
            .O(N__25842),
            .I(N__25839));
    InMux I__3740 (
            .O(N__25839),
            .I(N__25836));
    LocalMux I__3739 (
            .O(N__25836),
            .I(\ADC_VDC.n4_adj_1451 ));
    CEMux I__3738 (
            .O(N__25833),
            .I(N__25830));
    LocalMux I__3737 (
            .O(N__25830),
            .I(N__25827));
    Odrv4 I__3736 (
            .O(N__25827),
            .I(\ADC_VDC.n13503 ));
    InMux I__3735 (
            .O(N__25824),
            .I(N__25821));
    LocalMux I__3734 (
            .O(N__25821),
            .I(N__25818));
    Span4Mux_h I__3733 (
            .O(N__25818),
            .I(N__25814));
    InMux I__3732 (
            .O(N__25817),
            .I(N__25811));
    Odrv4 I__3731 (
            .O(N__25814),
            .I(buf_readRTD_8));
    LocalMux I__3730 (
            .O(N__25811),
            .I(buf_readRTD_8));
    InMux I__3729 (
            .O(N__25806),
            .I(N__25803));
    LocalMux I__3728 (
            .O(N__25803),
            .I(N__25800));
    Span4Mux_v I__3727 (
            .O(N__25800),
            .I(N__25796));
    CascadeMux I__3726 (
            .O(N__25799),
            .I(N__25793));
    Span4Mux_v I__3725 (
            .O(N__25796),
            .I(N__25790));
    InMux I__3724 (
            .O(N__25793),
            .I(N__25787));
    Odrv4 I__3723 (
            .O(N__25790),
            .I(buf_adcdata_vdc_16));
    LocalMux I__3722 (
            .O(N__25787),
            .I(buf_adcdata_vdc_16));
    InMux I__3721 (
            .O(N__25782),
            .I(N__25779));
    LocalMux I__3720 (
            .O(N__25779),
            .I(N__25775));
    InMux I__3719 (
            .O(N__25778),
            .I(N__25772));
    Span4Mux_v I__3718 (
            .O(N__25775),
            .I(N__25769));
    LocalMux I__3717 (
            .O(N__25772),
            .I(N__25766));
    Span4Mux_h I__3716 (
            .O(N__25769),
            .I(N__25763));
    Span4Mux_h I__3715 (
            .O(N__25766),
            .I(N__25759));
    Span4Mux_h I__3714 (
            .O(N__25763),
            .I(N__25756));
    InMux I__3713 (
            .O(N__25762),
            .I(N__25753));
    Span4Mux_v I__3712 (
            .O(N__25759),
            .I(N__25748));
    Span4Mux_h I__3711 (
            .O(N__25756),
            .I(N__25748));
    LocalMux I__3710 (
            .O(N__25753),
            .I(buf_adcdata_vac_16));
    Odrv4 I__3709 (
            .O(N__25748),
            .I(buf_adcdata_vac_16));
    CascadeMux I__3708 (
            .O(N__25743),
            .I(n22575_cascade_));
    CascadeMux I__3707 (
            .O(N__25740),
            .I(N__25736));
    InMux I__3706 (
            .O(N__25739),
            .I(N__25732));
    InMux I__3705 (
            .O(N__25736),
            .I(N__25729));
    InMux I__3704 (
            .O(N__25735),
            .I(N__25726));
    LocalMux I__3703 (
            .O(N__25732),
            .I(N__25723));
    LocalMux I__3702 (
            .O(N__25729),
            .I(N__25720));
    LocalMux I__3701 (
            .O(N__25726),
            .I(N__25717));
    Span12Mux_h I__3700 (
            .O(N__25723),
            .I(N__25712));
    Span4Mux_h I__3699 (
            .O(N__25720),
            .I(N__25709));
    Span4Mux_h I__3698 (
            .O(N__25717),
            .I(N__25706));
    InMux I__3697 (
            .O(N__25716),
            .I(N__25701));
    InMux I__3696 (
            .O(N__25715),
            .I(N__25701));
    Odrv12 I__3695 (
            .O(N__25712),
            .I(buf_cfgRTD_0));
    Odrv4 I__3694 (
            .O(N__25709),
            .I(buf_cfgRTD_0));
    Odrv4 I__3693 (
            .O(N__25706),
            .I(buf_cfgRTD_0));
    LocalMux I__3692 (
            .O(N__25701),
            .I(buf_cfgRTD_0));
    CascadeMux I__3691 (
            .O(N__25692),
            .I(n10902_cascade_));
    CascadeMux I__3690 (
            .O(N__25689),
            .I(n12624_cascade_));
    CascadeMux I__3689 (
            .O(N__25686),
            .I(N__25683));
    InMux I__3688 (
            .O(N__25683),
            .I(N__25680));
    LocalMux I__3687 (
            .O(N__25680),
            .I(N__25677));
    Span4Mux_v I__3686 (
            .O(N__25677),
            .I(N__25673));
    CascadeMux I__3685 (
            .O(N__25676),
            .I(N__25670));
    Span4Mux_h I__3684 (
            .O(N__25673),
            .I(N__25667));
    InMux I__3683 (
            .O(N__25670),
            .I(N__25664));
    Odrv4 I__3682 (
            .O(N__25667),
            .I(buf_adcdata_vdc_22));
    LocalMux I__3681 (
            .O(N__25664),
            .I(buf_adcdata_vdc_22));
    InMux I__3680 (
            .O(N__25659),
            .I(N__25655));
    InMux I__3679 (
            .O(N__25658),
            .I(N__25652));
    LocalMux I__3678 (
            .O(N__25655),
            .I(cmd_rdadcbuf_13));
    LocalMux I__3677 (
            .O(N__25652),
            .I(cmd_rdadcbuf_13));
    InMux I__3676 (
            .O(N__25647),
            .I(N__25644));
    LocalMux I__3675 (
            .O(N__25644),
            .I(N__25640));
    CascadeMux I__3674 (
            .O(N__25643),
            .I(N__25637));
    Span4Mux_h I__3673 (
            .O(N__25640),
            .I(N__25634));
    InMux I__3672 (
            .O(N__25637),
            .I(N__25631));
    Sp12to4 I__3671 (
            .O(N__25634),
            .I(N__25628));
    LocalMux I__3670 (
            .O(N__25631),
            .I(N__25625));
    Odrv12 I__3669 (
            .O(N__25628),
            .I(buf_adcdata_vdc_2));
    Odrv4 I__3668 (
            .O(N__25625),
            .I(buf_adcdata_vdc_2));
    InMux I__3667 (
            .O(N__25620),
            .I(N__25616));
    InMux I__3666 (
            .O(N__25619),
            .I(N__25613));
    LocalMux I__3665 (
            .O(N__25616),
            .I(cmd_rdadcbuf_15));
    LocalMux I__3664 (
            .O(N__25613),
            .I(cmd_rdadcbuf_15));
    InMux I__3663 (
            .O(N__25608),
            .I(N__25605));
    LocalMux I__3662 (
            .O(N__25605),
            .I(N__25601));
    CascadeMux I__3661 (
            .O(N__25604),
            .I(N__25598));
    Span4Mux_v I__3660 (
            .O(N__25601),
            .I(N__25595));
    InMux I__3659 (
            .O(N__25598),
            .I(N__25592));
    Odrv4 I__3658 (
            .O(N__25595),
            .I(buf_adcdata_vdc_4));
    LocalMux I__3657 (
            .O(N__25592),
            .I(buf_adcdata_vdc_4));
    InMux I__3656 (
            .O(N__25587),
            .I(N__25583));
    InMux I__3655 (
            .O(N__25586),
            .I(N__25580));
    LocalMux I__3654 (
            .O(N__25583),
            .I(cmd_rdadcbuf_16));
    LocalMux I__3653 (
            .O(N__25580),
            .I(cmd_rdadcbuf_16));
    InMux I__3652 (
            .O(N__25575),
            .I(N__25572));
    LocalMux I__3651 (
            .O(N__25572),
            .I(N__25568));
    CascadeMux I__3650 (
            .O(N__25571),
            .I(N__25565));
    Span4Mux_v I__3649 (
            .O(N__25568),
            .I(N__25562));
    InMux I__3648 (
            .O(N__25565),
            .I(N__25559));
    Odrv4 I__3647 (
            .O(N__25562),
            .I(buf_adcdata_vdc_5));
    LocalMux I__3646 (
            .O(N__25559),
            .I(buf_adcdata_vdc_5));
    CascadeMux I__3645 (
            .O(N__25554),
            .I(N__25550));
    InMux I__3644 (
            .O(N__25553),
            .I(N__25546));
    InMux I__3643 (
            .O(N__25550),
            .I(N__25543));
    InMux I__3642 (
            .O(N__25549),
            .I(N__25540));
    LocalMux I__3641 (
            .O(N__25546),
            .I(N__25535));
    LocalMux I__3640 (
            .O(N__25543),
            .I(N__25535));
    LocalMux I__3639 (
            .O(N__25540),
            .I(cmd_rdadctmp_20_adj_1503));
    Odrv4 I__3638 (
            .O(N__25535),
            .I(cmd_rdadctmp_20_adj_1503));
    InMux I__3637 (
            .O(N__25530),
            .I(N__25526));
    CascadeMux I__3636 (
            .O(N__25529),
            .I(N__25522));
    LocalMux I__3635 (
            .O(N__25526),
            .I(N__25519));
    InMux I__3634 (
            .O(N__25525),
            .I(N__25516));
    InMux I__3633 (
            .O(N__25522),
            .I(N__25513));
    Odrv12 I__3632 (
            .O(N__25519),
            .I(cmd_rdadctmp_21_adj_1502));
    LocalMux I__3631 (
            .O(N__25516),
            .I(cmd_rdadctmp_21_adj_1502));
    LocalMux I__3630 (
            .O(N__25513),
            .I(cmd_rdadctmp_21_adj_1502));
    InMux I__3629 (
            .O(N__25506),
            .I(N__25503));
    LocalMux I__3628 (
            .O(N__25503),
            .I(\ADC_VDC.cmd_rdadcbuf_35_N_1296_34 ));
    InMux I__3627 (
            .O(N__25500),
            .I(N__25497));
    LocalMux I__3626 (
            .O(N__25497),
            .I(N__25494));
    Odrv4 I__3625 (
            .O(N__25494),
            .I(\ADC_VDC.n19 ));
    CascadeMux I__3624 (
            .O(N__25491),
            .I(\ADC_VDC.n21_cascade_ ));
    CascadeMux I__3623 (
            .O(N__25488),
            .I(N__25483));
    InMux I__3622 (
            .O(N__25487),
            .I(N__25478));
    InMux I__3621 (
            .O(N__25486),
            .I(N__25478));
    InMux I__3620 (
            .O(N__25483),
            .I(N__25475));
    LocalMux I__3619 (
            .O(N__25478),
            .I(cmd_rdadctmp_14_adj_1509));
    LocalMux I__3618 (
            .O(N__25475),
            .I(cmd_rdadctmp_14_adj_1509));
    CascadeMux I__3617 (
            .O(N__25470),
            .I(N__25465));
    InMux I__3616 (
            .O(N__25469),
            .I(N__25462));
    InMux I__3615 (
            .O(N__25468),
            .I(N__25459));
    InMux I__3614 (
            .O(N__25465),
            .I(N__25456));
    LocalMux I__3613 (
            .O(N__25462),
            .I(cmd_rdadctmp_15_adj_1508));
    LocalMux I__3612 (
            .O(N__25459),
            .I(cmd_rdadctmp_15_adj_1508));
    LocalMux I__3611 (
            .O(N__25456),
            .I(cmd_rdadctmp_15_adj_1508));
    InMux I__3610 (
            .O(N__25449),
            .I(N__25445));
    InMux I__3609 (
            .O(N__25448),
            .I(N__25442));
    LocalMux I__3608 (
            .O(N__25445),
            .I(cmd_rdadcbuf_20));
    LocalMux I__3607 (
            .O(N__25442),
            .I(cmd_rdadcbuf_20));
    InMux I__3606 (
            .O(N__25437),
            .I(N__25434));
    LocalMux I__3605 (
            .O(N__25434),
            .I(N__25431));
    Span4Mux_v I__3604 (
            .O(N__25431),
            .I(N__25427));
    InMux I__3603 (
            .O(N__25430),
            .I(N__25424));
    Odrv4 I__3602 (
            .O(N__25427),
            .I(buf_adcdata_vdc_9));
    LocalMux I__3601 (
            .O(N__25424),
            .I(buf_adcdata_vdc_9));
    InMux I__3600 (
            .O(N__25419),
            .I(N__25415));
    InMux I__3599 (
            .O(N__25418),
            .I(N__25412));
    LocalMux I__3598 (
            .O(N__25415),
            .I(N__25409));
    LocalMux I__3597 (
            .O(N__25412),
            .I(cmd_rdadcbuf_17));
    Odrv4 I__3596 (
            .O(N__25409),
            .I(cmd_rdadcbuf_17));
    InMux I__3595 (
            .O(N__25404),
            .I(N__25401));
    LocalMux I__3594 (
            .O(N__25401),
            .I(N__25398));
    Span4Mux_h I__3593 (
            .O(N__25398),
            .I(N__25394));
    CascadeMux I__3592 (
            .O(N__25397),
            .I(N__25391));
    Span4Mux_v I__3591 (
            .O(N__25394),
            .I(N__25388));
    InMux I__3590 (
            .O(N__25391),
            .I(N__25385));
    Odrv4 I__3589 (
            .O(N__25388),
            .I(buf_adcdata_vdc_6));
    LocalMux I__3588 (
            .O(N__25385),
            .I(buf_adcdata_vdc_6));
    InMux I__3587 (
            .O(N__25380),
            .I(N__25376));
    InMux I__3586 (
            .O(N__25379),
            .I(N__25373));
    LocalMux I__3585 (
            .O(N__25376),
            .I(cmd_rdadcbuf_11));
    LocalMux I__3584 (
            .O(N__25373),
            .I(cmd_rdadcbuf_11));
    InMux I__3583 (
            .O(N__25368),
            .I(N__25365));
    LocalMux I__3582 (
            .O(N__25365),
            .I(N__25360));
    InMux I__3581 (
            .O(N__25364),
            .I(N__25357));
    InMux I__3580 (
            .O(N__25363),
            .I(N__25354));
    Span4Mux_v I__3579 (
            .O(N__25360),
            .I(N__25351));
    LocalMux I__3578 (
            .O(N__25357),
            .I(buf_dds1_5));
    LocalMux I__3577 (
            .O(N__25354),
            .I(buf_dds1_5));
    Odrv4 I__3576 (
            .O(N__25351),
            .I(buf_dds1_5));
    InMux I__3575 (
            .O(N__25344),
            .I(N__25340));
    InMux I__3574 (
            .O(N__25343),
            .I(N__25337));
    LocalMux I__3573 (
            .O(N__25340),
            .I(cmd_rdadcbuf_21));
    LocalMux I__3572 (
            .O(N__25337),
            .I(cmd_rdadcbuf_21));
    InMux I__3571 (
            .O(N__25332),
            .I(N__25329));
    LocalMux I__3570 (
            .O(N__25329),
            .I(N__25325));
    InMux I__3569 (
            .O(N__25328),
            .I(N__25322));
    Odrv4 I__3568 (
            .O(N__25325),
            .I(cmd_rdadcbuf_33));
    LocalMux I__3567 (
            .O(N__25322),
            .I(cmd_rdadcbuf_33));
    InMux I__3566 (
            .O(N__25317),
            .I(N__25310));
    InMux I__3565 (
            .O(N__25316),
            .I(N__25310));
    InMux I__3564 (
            .O(N__25315),
            .I(N__25307));
    LocalMux I__3563 (
            .O(N__25310),
            .I(cmd_rdadctmp_4_adj_1519));
    LocalMux I__3562 (
            .O(N__25307),
            .I(cmd_rdadctmp_4_adj_1519));
    CascadeMux I__3561 (
            .O(N__25302),
            .I(N__25297));
    InMux I__3560 (
            .O(N__25301),
            .I(N__25294));
    InMux I__3559 (
            .O(N__25300),
            .I(N__25291));
    InMux I__3558 (
            .O(N__25297),
            .I(N__25288));
    LocalMux I__3557 (
            .O(N__25294),
            .I(cmd_rdadctmp_5_adj_1518));
    LocalMux I__3556 (
            .O(N__25291),
            .I(cmd_rdadctmp_5_adj_1518));
    LocalMux I__3555 (
            .O(N__25288),
            .I(cmd_rdadctmp_5_adj_1518));
    CascadeMux I__3554 (
            .O(N__25281),
            .I(N__25278));
    InMux I__3553 (
            .O(N__25278),
            .I(N__25273));
    InMux I__3552 (
            .O(N__25277),
            .I(N__25270));
    InMux I__3551 (
            .O(N__25276),
            .I(N__25267));
    LocalMux I__3550 (
            .O(N__25273),
            .I(cmd_rdadctmp_7_adj_1516));
    LocalMux I__3549 (
            .O(N__25270),
            .I(cmd_rdadctmp_7_adj_1516));
    LocalMux I__3548 (
            .O(N__25267),
            .I(cmd_rdadctmp_7_adj_1516));
    InMux I__3547 (
            .O(N__25260),
            .I(N__25255));
    InMux I__3546 (
            .O(N__25259),
            .I(N__25252));
    InMux I__3545 (
            .O(N__25258),
            .I(N__25249));
    LocalMux I__3544 (
            .O(N__25255),
            .I(N__25246));
    LocalMux I__3543 (
            .O(N__25252),
            .I(cmd_rdadctmp_19_adj_1504));
    LocalMux I__3542 (
            .O(N__25249),
            .I(cmd_rdadctmp_19_adj_1504));
    Odrv4 I__3541 (
            .O(N__25246),
            .I(cmd_rdadctmp_19_adj_1504));
    CascadeMux I__3540 (
            .O(N__25239),
            .I(N__25235));
    CascadeMux I__3539 (
            .O(N__25238),
            .I(N__25231));
    InMux I__3538 (
            .O(N__25235),
            .I(N__25228));
    InMux I__3537 (
            .O(N__25234),
            .I(N__25225));
    InMux I__3536 (
            .O(N__25231),
            .I(N__25222));
    LocalMux I__3535 (
            .O(N__25228),
            .I(cmd_rdadctmp_8_adj_1515));
    LocalMux I__3534 (
            .O(N__25225),
            .I(cmd_rdadctmp_8_adj_1515));
    LocalMux I__3533 (
            .O(N__25222),
            .I(cmd_rdadctmp_8_adj_1515));
    CascadeMux I__3532 (
            .O(N__25215),
            .I(N__25210));
    InMux I__3531 (
            .O(N__25214),
            .I(N__25207));
    InMux I__3530 (
            .O(N__25213),
            .I(N__25204));
    InMux I__3529 (
            .O(N__25210),
            .I(N__25201));
    LocalMux I__3528 (
            .O(N__25207),
            .I(cmd_rdadctmp_9_adj_1514));
    LocalMux I__3527 (
            .O(N__25204),
            .I(cmd_rdadctmp_9_adj_1514));
    LocalMux I__3526 (
            .O(N__25201),
            .I(cmd_rdadctmp_9_adj_1514));
    CascadeMux I__3525 (
            .O(N__25194),
            .I(N__25190));
    CascadeMux I__3524 (
            .O(N__25193),
            .I(N__25186));
    InMux I__3523 (
            .O(N__25190),
            .I(N__25183));
    InMux I__3522 (
            .O(N__25189),
            .I(N__25180));
    InMux I__3521 (
            .O(N__25186),
            .I(N__25177));
    LocalMux I__3520 (
            .O(N__25183),
            .I(N__25174));
    LocalMux I__3519 (
            .O(N__25180),
            .I(cmd_rdadctmp_10_adj_1513));
    LocalMux I__3518 (
            .O(N__25177),
            .I(cmd_rdadctmp_10_adj_1513));
    Odrv4 I__3517 (
            .O(N__25174),
            .I(cmd_rdadctmp_10_adj_1513));
    CascadeMux I__3516 (
            .O(N__25167),
            .I(N__25162));
    InMux I__3515 (
            .O(N__25166),
            .I(N__25157));
    InMux I__3514 (
            .O(N__25165),
            .I(N__25157));
    InMux I__3513 (
            .O(N__25162),
            .I(N__25154));
    LocalMux I__3512 (
            .O(N__25157),
            .I(cmd_rdadctmp_11_adj_1512));
    LocalMux I__3511 (
            .O(N__25154),
            .I(cmd_rdadctmp_11_adj_1512));
    InMux I__3510 (
            .O(N__25149),
            .I(N__25142));
    InMux I__3509 (
            .O(N__25148),
            .I(N__25142));
    InMux I__3508 (
            .O(N__25147),
            .I(N__25139));
    LocalMux I__3507 (
            .O(N__25142),
            .I(cmd_rdadctmp_12_adj_1511));
    LocalMux I__3506 (
            .O(N__25139),
            .I(cmd_rdadctmp_12_adj_1511));
    CascadeMux I__3505 (
            .O(N__25134),
            .I(N__25130));
    CascadeMux I__3504 (
            .O(N__25133),
            .I(N__25127));
    InMux I__3503 (
            .O(N__25130),
            .I(N__25121));
    InMux I__3502 (
            .O(N__25127),
            .I(N__25121));
    CascadeMux I__3501 (
            .O(N__25126),
            .I(N__25118));
    LocalMux I__3500 (
            .O(N__25121),
            .I(N__25115));
    InMux I__3499 (
            .O(N__25118),
            .I(N__25112));
    Odrv4 I__3498 (
            .O(N__25115),
            .I(cmd_rdadctmp_13_adj_1510));
    LocalMux I__3497 (
            .O(N__25112),
            .I(cmd_rdadctmp_13_adj_1510));
    InMux I__3496 (
            .O(N__25107),
            .I(N__25104));
    LocalMux I__3495 (
            .O(N__25104),
            .I(N__25101));
    Span4Mux_v I__3494 (
            .O(N__25101),
            .I(N__25097));
    InMux I__3493 (
            .O(N__25100),
            .I(N__25094));
    Odrv4 I__3492 (
            .O(N__25097),
            .I(cmd_rdadcbuf_27));
    LocalMux I__3491 (
            .O(N__25094),
            .I(cmd_rdadcbuf_27));
    CascadeMux I__3490 (
            .O(N__25089),
            .I(\ADC_VDC.n10309_cascade_ ));
    CEMux I__3489 (
            .O(N__25086),
            .I(N__25083));
    LocalMux I__3488 (
            .O(N__25083),
            .I(N__25080));
    Span4Mux_v I__3487 (
            .O(N__25080),
            .I(N__25077));
    Odrv4 I__3486 (
            .O(N__25077),
            .I(\ADC_VDC.n13276 ));
    CascadeMux I__3485 (
            .O(N__25074),
            .I(N__25069));
    CascadeMux I__3484 (
            .O(N__25073),
            .I(N__25066));
    CascadeMux I__3483 (
            .O(N__25072),
            .I(N__25063));
    InMux I__3482 (
            .O(N__25069),
            .I(N__25060));
    InMux I__3481 (
            .O(N__25066),
            .I(N__25057));
    InMux I__3480 (
            .O(N__25063),
            .I(N__25054));
    LocalMux I__3479 (
            .O(N__25060),
            .I(cmd_rdadctmp_1_adj_1522));
    LocalMux I__3478 (
            .O(N__25057),
            .I(cmd_rdadctmp_1_adj_1522));
    LocalMux I__3477 (
            .O(N__25054),
            .I(cmd_rdadctmp_1_adj_1522));
    CascadeMux I__3476 (
            .O(N__25047),
            .I(N__25042));
    InMux I__3475 (
            .O(N__25046),
            .I(N__25037));
    InMux I__3474 (
            .O(N__25045),
            .I(N__25037));
    InMux I__3473 (
            .O(N__25042),
            .I(N__25034));
    LocalMux I__3472 (
            .O(N__25037),
            .I(cmd_rdadctmp_2_adj_1521));
    LocalMux I__3471 (
            .O(N__25034),
            .I(cmd_rdadctmp_2_adj_1521));
    CascadeMux I__3470 (
            .O(N__25029),
            .I(N__25024));
    InMux I__3469 (
            .O(N__25028),
            .I(N__25019));
    InMux I__3468 (
            .O(N__25027),
            .I(N__25019));
    InMux I__3467 (
            .O(N__25024),
            .I(N__25016));
    LocalMux I__3466 (
            .O(N__25019),
            .I(cmd_rdadctmp_3_adj_1520));
    LocalMux I__3465 (
            .O(N__25016),
            .I(cmd_rdadctmp_3_adj_1520));
    CascadeMux I__3464 (
            .O(N__25011),
            .I(\ADC_IAC.n21159_cascade_ ));
    CEMux I__3463 (
            .O(N__25008),
            .I(N__25005));
    LocalMux I__3462 (
            .O(N__25005),
            .I(N__25002));
    Odrv12 I__3461 (
            .O(N__25002),
            .I(\ADC_IAC.n21160 ));
    InMux I__3460 (
            .O(N__24999),
            .I(N__24993));
    InMux I__3459 (
            .O(N__24998),
            .I(N__24993));
    LocalMux I__3458 (
            .O(N__24993),
            .I(cmd_rdadctmp_1));
    CascadeMux I__3457 (
            .O(N__24990),
            .I(N__24986));
    InMux I__3456 (
            .O(N__24989),
            .I(N__24983));
    InMux I__3455 (
            .O(N__24986),
            .I(N__24980));
    LocalMux I__3454 (
            .O(N__24983),
            .I(cmd_rdadctmp_2));
    LocalMux I__3453 (
            .O(N__24980),
            .I(cmd_rdadctmp_2));
    CascadeMux I__3452 (
            .O(N__24975),
            .I(N__24972));
    InMux I__3451 (
            .O(N__24972),
            .I(N__24969));
    LocalMux I__3450 (
            .O(N__24969),
            .I(N__24966));
    Span4Mux_v I__3449 (
            .O(N__24966),
            .I(N__24963));
    Sp12to4 I__3448 (
            .O(N__24963),
            .I(N__24960));
    Span12Mux_h I__3447 (
            .O(N__24960),
            .I(N__24957));
    Odrv12 I__3446 (
            .O(N__24957),
            .I(IAC_MISO));
    CascadeMux I__3445 (
            .O(N__24954),
            .I(N__24951));
    InMux I__3444 (
            .O(N__24951),
            .I(N__24945));
    InMux I__3443 (
            .O(N__24950),
            .I(N__24945));
    LocalMux I__3442 (
            .O(N__24945),
            .I(cmd_rdadctmp_0));
    CascadeMux I__3441 (
            .O(N__24942),
            .I(N__24936));
    InMux I__3440 (
            .O(N__24941),
            .I(N__24932));
    CascadeMux I__3439 (
            .O(N__24940),
            .I(N__24929));
    InMux I__3438 (
            .O(N__24939),
            .I(N__24919));
    InMux I__3437 (
            .O(N__24936),
            .I(N__24919));
    InMux I__3436 (
            .O(N__24935),
            .I(N__24919));
    LocalMux I__3435 (
            .O(N__24932),
            .I(N__24915));
    InMux I__3434 (
            .O(N__24929),
            .I(N__24912));
    CascadeMux I__3433 (
            .O(N__24928),
            .I(N__24909));
    CascadeMux I__3432 (
            .O(N__24927),
            .I(N__24905));
    InMux I__3431 (
            .O(N__24926),
            .I(N__24900));
    LocalMux I__3430 (
            .O(N__24919),
            .I(N__24897));
    InMux I__3429 (
            .O(N__24918),
            .I(N__24894));
    Span4Mux_v I__3428 (
            .O(N__24915),
            .I(N__24891));
    LocalMux I__3427 (
            .O(N__24912),
            .I(N__24888));
    InMux I__3426 (
            .O(N__24909),
            .I(N__24885));
    InMux I__3425 (
            .O(N__24908),
            .I(N__24878));
    InMux I__3424 (
            .O(N__24905),
            .I(N__24878));
    InMux I__3423 (
            .O(N__24904),
            .I(N__24878));
    InMux I__3422 (
            .O(N__24903),
            .I(N__24875));
    LocalMux I__3421 (
            .O(N__24900),
            .I(N__24868));
    Span4Mux_v I__3420 (
            .O(N__24897),
            .I(N__24868));
    LocalMux I__3419 (
            .O(N__24894),
            .I(N__24868));
    Odrv4 I__3418 (
            .O(N__24891),
            .I(DTRIG_N_958));
    Odrv4 I__3417 (
            .O(N__24888),
            .I(DTRIG_N_958));
    LocalMux I__3416 (
            .O(N__24885),
            .I(DTRIG_N_958));
    LocalMux I__3415 (
            .O(N__24878),
            .I(DTRIG_N_958));
    LocalMux I__3414 (
            .O(N__24875),
            .I(DTRIG_N_958));
    Odrv4 I__3413 (
            .O(N__24868),
            .I(DTRIG_N_958));
    InMux I__3412 (
            .O(N__24855),
            .I(N__24847));
    InMux I__3411 (
            .O(N__24854),
            .I(N__24843));
    InMux I__3410 (
            .O(N__24853),
            .I(N__24834));
    InMux I__3409 (
            .O(N__24852),
            .I(N__24834));
    InMux I__3408 (
            .O(N__24851),
            .I(N__24829));
    InMux I__3407 (
            .O(N__24850),
            .I(N__24829));
    LocalMux I__3406 (
            .O(N__24847),
            .I(N__24825));
    InMux I__3405 (
            .O(N__24846),
            .I(N__24822));
    LocalMux I__3404 (
            .O(N__24843),
            .I(N__24819));
    InMux I__3403 (
            .O(N__24842),
            .I(N__24816));
    InMux I__3402 (
            .O(N__24841),
            .I(N__24809));
    InMux I__3401 (
            .O(N__24840),
            .I(N__24809));
    InMux I__3400 (
            .O(N__24839),
            .I(N__24809));
    LocalMux I__3399 (
            .O(N__24834),
            .I(N__24804));
    LocalMux I__3398 (
            .O(N__24829),
            .I(N__24804));
    InMux I__3397 (
            .O(N__24828),
            .I(N__24801));
    Odrv4 I__3396 (
            .O(N__24825),
            .I(adc_state_1));
    LocalMux I__3395 (
            .O(N__24822),
            .I(adc_state_1));
    Odrv4 I__3394 (
            .O(N__24819),
            .I(adc_state_1));
    LocalMux I__3393 (
            .O(N__24816),
            .I(adc_state_1));
    LocalMux I__3392 (
            .O(N__24809),
            .I(adc_state_1));
    Odrv4 I__3391 (
            .O(N__24804),
            .I(adc_state_1));
    LocalMux I__3390 (
            .O(N__24801),
            .I(adc_state_1));
    IoInMux I__3389 (
            .O(N__24786),
            .I(N__24783));
    LocalMux I__3388 (
            .O(N__24783),
            .I(N__24780));
    IoSpan4Mux I__3387 (
            .O(N__24780),
            .I(N__24777));
    Span4Mux_s3_v I__3386 (
            .O(N__24777),
            .I(N__24773));
    CascadeMux I__3385 (
            .O(N__24776),
            .I(N__24770));
    Span4Mux_v I__3384 (
            .O(N__24773),
            .I(N__24767));
    InMux I__3383 (
            .O(N__24770),
            .I(N__24764));
    Odrv4 I__3382 (
            .O(N__24767),
            .I(IAC_SCLK));
    LocalMux I__3381 (
            .O(N__24764),
            .I(IAC_SCLK));
    InMux I__3380 (
            .O(N__24759),
            .I(N__24756));
    LocalMux I__3379 (
            .O(N__24756),
            .I(N__24753));
    Span4Mux_h I__3378 (
            .O(N__24753),
            .I(N__24750));
    Span4Mux_v I__3377 (
            .O(N__24750),
            .I(N__24746));
    InMux I__3376 (
            .O(N__24749),
            .I(N__24743));
    Span4Mux_v I__3375 (
            .O(N__24746),
            .I(N__24739));
    LocalMux I__3374 (
            .O(N__24743),
            .I(N__24736));
    InMux I__3373 (
            .O(N__24742),
            .I(N__24733));
    Sp12to4 I__3372 (
            .O(N__24739),
            .I(N__24730));
    Span4Mux_h I__3371 (
            .O(N__24736),
            .I(N__24727));
    LocalMux I__3370 (
            .O(N__24733),
            .I(buf_adcdata_iac_17));
    Odrv12 I__3369 (
            .O(N__24730),
            .I(buf_adcdata_iac_17));
    Odrv4 I__3368 (
            .O(N__24727),
            .I(buf_adcdata_iac_17));
    InMux I__3367 (
            .O(N__24720),
            .I(N__24717));
    LocalMux I__3366 (
            .O(N__24717),
            .I(N__24714));
    Span4Mux_v I__3365 (
            .O(N__24714),
            .I(N__24710));
    InMux I__3364 (
            .O(N__24713),
            .I(N__24707));
    Odrv4 I__3363 (
            .O(N__24710),
            .I(cmd_rdadctmp_4_adj_1488));
    LocalMux I__3362 (
            .O(N__24707),
            .I(cmd_rdadctmp_4_adj_1488));
    CascadeMux I__3361 (
            .O(N__24702),
            .I(N__24699));
    InMux I__3360 (
            .O(N__24699),
            .I(N__24693));
    InMux I__3359 (
            .O(N__24698),
            .I(N__24693));
    LocalMux I__3358 (
            .O(N__24693),
            .I(cmd_rdadctmp_5_adj_1487));
    CascadeMux I__3357 (
            .O(N__24690),
            .I(N__24687));
    InMux I__3356 (
            .O(N__24687),
            .I(N__24684));
    LocalMux I__3355 (
            .O(N__24684),
            .I(N__24681));
    Span4Mux_h I__3354 (
            .O(N__24681),
            .I(N__24677));
    InMux I__3353 (
            .O(N__24680),
            .I(N__24674));
    Odrv4 I__3352 (
            .O(N__24677),
            .I(cmd_rdadctmp_6_adj_1486));
    LocalMux I__3351 (
            .O(N__24674),
            .I(cmd_rdadctmp_6_adj_1486));
    CascadeMux I__3350 (
            .O(N__24669),
            .I(N__24666));
    InMux I__3349 (
            .O(N__24666),
            .I(N__24663));
    LocalMux I__3348 (
            .O(N__24663),
            .I(N__24660));
    Span4Mux_v I__3347 (
            .O(N__24660),
            .I(N__24655));
    InMux I__3346 (
            .O(N__24659),
            .I(N__24650));
    InMux I__3345 (
            .O(N__24658),
            .I(N__24650));
    Odrv4 I__3344 (
            .O(N__24655),
            .I(cmd_rdadctmp_22));
    LocalMux I__3343 (
            .O(N__24650),
            .I(cmd_rdadctmp_22));
    SRMux I__3342 (
            .O(N__24645),
            .I(N__24642));
    LocalMux I__3341 (
            .O(N__24642),
            .I(N__24638));
    CascadeMux I__3340 (
            .O(N__24641),
            .I(N__24635));
    Span4Mux_h I__3339 (
            .O(N__24638),
            .I(N__24632));
    InMux I__3338 (
            .O(N__24635),
            .I(N__24629));
    Odrv4 I__3337 (
            .O(N__24632),
            .I(n15092));
    LocalMux I__3336 (
            .O(N__24629),
            .I(n15092));
    CascadeMux I__3335 (
            .O(N__24624),
            .I(N__24620));
    CascadeMux I__3334 (
            .O(N__24623),
            .I(N__24617));
    InMux I__3333 (
            .O(N__24620),
            .I(N__24612));
    InMux I__3332 (
            .O(N__24617),
            .I(N__24607));
    InMux I__3331 (
            .O(N__24616),
            .I(N__24607));
    CascadeMux I__3330 (
            .O(N__24615),
            .I(N__24603));
    LocalMux I__3329 (
            .O(N__24612),
            .I(N__24598));
    LocalMux I__3328 (
            .O(N__24607),
            .I(N__24598));
    InMux I__3327 (
            .O(N__24606),
            .I(N__24595));
    InMux I__3326 (
            .O(N__24603),
            .I(N__24592));
    Span4Mux_v I__3325 (
            .O(N__24598),
            .I(N__24587));
    LocalMux I__3324 (
            .O(N__24595),
            .I(N__24587));
    LocalMux I__3323 (
            .O(N__24592),
            .I(N__24582));
    Sp12to4 I__3322 (
            .O(N__24587),
            .I(N__24582));
    Span12Mux_h I__3321 (
            .O(N__24582),
            .I(N__24579));
    Odrv12 I__3320 (
            .O(N__24579),
            .I(IAC_DRDY));
    CascadeMux I__3319 (
            .O(N__24576),
            .I(N__24573));
    InMux I__3318 (
            .O(N__24573),
            .I(N__24570));
    LocalMux I__3317 (
            .O(N__24570),
            .I(\CLK_DDS.tmp_buf_3 ));
    CascadeMux I__3316 (
            .O(N__24567),
            .I(N__24564));
    InMux I__3315 (
            .O(N__24564),
            .I(N__24561));
    LocalMux I__3314 (
            .O(N__24561),
            .I(\CLK_DDS.tmp_buf_4 ));
    CascadeMux I__3313 (
            .O(N__24558),
            .I(N__24555));
    InMux I__3312 (
            .O(N__24555),
            .I(N__24552));
    LocalMux I__3311 (
            .O(N__24552),
            .I(\CLK_DDS.tmp_buf_5 ));
    CascadeMux I__3310 (
            .O(N__24549),
            .I(N__24546));
    InMux I__3309 (
            .O(N__24546),
            .I(N__24543));
    LocalMux I__3308 (
            .O(N__24543),
            .I(\CLK_DDS.tmp_buf_6 ));
    CascadeMux I__3307 (
            .O(N__24540),
            .I(N__24537));
    InMux I__3306 (
            .O(N__24537),
            .I(N__24534));
    LocalMux I__3305 (
            .O(N__24534),
            .I(N__24531));
    Odrv12 I__3304 (
            .O(N__24531),
            .I(\CLK_DDS.tmp_buf_7 ));
    InMux I__3303 (
            .O(N__24528),
            .I(N__24525));
    LocalMux I__3302 (
            .O(N__24525),
            .I(N__24522));
    Span12Mux_s8_h I__3301 (
            .O(N__24522),
            .I(N__24517));
    InMux I__3300 (
            .O(N__24521),
            .I(N__24514));
    InMux I__3299 (
            .O(N__24520),
            .I(N__24511));
    Span12Mux_h I__3298 (
            .O(N__24517),
            .I(N__24508));
    LocalMux I__3297 (
            .O(N__24514),
            .I(N__24505));
    LocalMux I__3296 (
            .O(N__24511),
            .I(buf_adcdata_vac_17));
    Odrv12 I__3295 (
            .O(N__24508),
            .I(buf_adcdata_vac_17));
    Odrv12 I__3294 (
            .O(N__24505),
            .I(buf_adcdata_vac_17));
    CascadeMux I__3293 (
            .O(N__24498),
            .I(N__24494));
    InMux I__3292 (
            .O(N__24497),
            .I(N__24487));
    InMux I__3291 (
            .O(N__24494),
            .I(N__24487));
    InMux I__3290 (
            .O(N__24493),
            .I(N__24484));
    InMux I__3289 (
            .O(N__24492),
            .I(N__24481));
    LocalMux I__3288 (
            .O(N__24487),
            .I(\SIG_DDS.bit_cnt_1 ));
    LocalMux I__3287 (
            .O(N__24484),
            .I(\SIG_DDS.bit_cnt_1 ));
    LocalMux I__3286 (
            .O(N__24481),
            .I(\SIG_DDS.bit_cnt_1 ));
    InMux I__3285 (
            .O(N__24474),
            .I(N__24467));
    InMux I__3284 (
            .O(N__24473),
            .I(N__24467));
    CascadeMux I__3283 (
            .O(N__24472),
            .I(N__24464));
    LocalMux I__3282 (
            .O(N__24467),
            .I(N__24461));
    InMux I__3281 (
            .O(N__24464),
            .I(N__24458));
    Odrv4 I__3280 (
            .O(N__24461),
            .I(\SIG_DDS.bit_cnt_2 ));
    LocalMux I__3279 (
            .O(N__24458),
            .I(\SIG_DDS.bit_cnt_2 ));
    CascadeMux I__3278 (
            .O(N__24453),
            .I(N__24450));
    InMux I__3277 (
            .O(N__24450),
            .I(N__24447));
    LocalMux I__3276 (
            .O(N__24447),
            .I(N__24444));
    Odrv4 I__3275 (
            .O(N__24444),
            .I(\SIG_DDS.n10 ));
    InMux I__3274 (
            .O(N__24441),
            .I(N__24430));
    InMux I__3273 (
            .O(N__24440),
            .I(N__24430));
    InMux I__3272 (
            .O(N__24439),
            .I(N__24430));
    InMux I__3271 (
            .O(N__24438),
            .I(N__24427));
    InMux I__3270 (
            .O(N__24437),
            .I(N__24424));
    LocalMux I__3269 (
            .O(N__24430),
            .I(bit_cnt_0));
    LocalMux I__3268 (
            .O(N__24427),
            .I(bit_cnt_0));
    LocalMux I__3267 (
            .O(N__24424),
            .I(bit_cnt_0));
    CascadeMux I__3266 (
            .O(N__24417),
            .I(N__24413));
    CascadeMux I__3265 (
            .O(N__24416),
            .I(N__24409));
    InMux I__3264 (
            .O(N__24413),
            .I(N__24406));
    InMux I__3263 (
            .O(N__24412),
            .I(N__24401));
    InMux I__3262 (
            .O(N__24409),
            .I(N__24401));
    LocalMux I__3261 (
            .O(N__24406),
            .I(cmd_rdadctmp_28_adj_1464));
    LocalMux I__3260 (
            .O(N__24401),
            .I(cmd_rdadctmp_28_adj_1464));
    InMux I__3259 (
            .O(N__24396),
            .I(N__24393));
    LocalMux I__3258 (
            .O(N__24393),
            .I(N__24389));
    InMux I__3257 (
            .O(N__24392),
            .I(N__24386));
    Odrv12 I__3256 (
            .O(N__24389),
            .I(tmp_buf_15_adj_1497));
    LocalMux I__3255 (
            .O(N__24386),
            .I(tmp_buf_15_adj_1497));
    CascadeMux I__3254 (
            .O(N__24381),
            .I(N__24378));
    InMux I__3253 (
            .O(N__24378),
            .I(N__24375));
    LocalMux I__3252 (
            .O(N__24375),
            .I(\CLK_DDS.tmp_buf_0 ));
    InMux I__3251 (
            .O(N__24372),
            .I(N__24369));
    LocalMux I__3250 (
            .O(N__24369),
            .I(\CLK_DDS.tmp_buf_1 ));
    CascadeMux I__3249 (
            .O(N__24366),
            .I(N__24363));
    InMux I__3248 (
            .O(N__24363),
            .I(N__24360));
    LocalMux I__3247 (
            .O(N__24360),
            .I(\CLK_DDS.tmp_buf_2 ));
    InMux I__3246 (
            .O(N__24357),
            .I(N__24354));
    LocalMux I__3245 (
            .O(N__24354),
            .I(N__24350));
    InMux I__3244 (
            .O(N__24353),
            .I(N__24347));
    Span4Mux_h I__3243 (
            .O(N__24350),
            .I(N__24343));
    LocalMux I__3242 (
            .O(N__24347),
            .I(N__24340));
    InMux I__3241 (
            .O(N__24346),
            .I(N__24337));
    Odrv4 I__3240 (
            .O(N__24343),
            .I(cmd_rdadctmp_13));
    Odrv4 I__3239 (
            .O(N__24340),
            .I(cmd_rdadctmp_13));
    LocalMux I__3238 (
            .O(N__24337),
            .I(cmd_rdadctmp_13));
    InMux I__3237 (
            .O(N__24330),
            .I(N__24327));
    LocalMux I__3236 (
            .O(N__24327),
            .I(N__24323));
    CascadeMux I__3235 (
            .O(N__24326),
            .I(N__24320));
    Span4Mux_h I__3234 (
            .O(N__24323),
            .I(N__24317));
    InMux I__3233 (
            .O(N__24320),
            .I(N__24314));
    Sp12to4 I__3232 (
            .O(N__24317),
            .I(N__24308));
    LocalMux I__3231 (
            .O(N__24314),
            .I(N__24308));
    InMux I__3230 (
            .O(N__24313),
            .I(N__24305));
    Odrv12 I__3229 (
            .O(N__24308),
            .I(cmd_rdadctmp_10));
    LocalMux I__3228 (
            .O(N__24305),
            .I(cmd_rdadctmp_10));
    InMux I__3227 (
            .O(N__24300),
            .I(N__24297));
    LocalMux I__3226 (
            .O(N__24297),
            .I(N__24294));
    Span4Mux_v I__3225 (
            .O(N__24294),
            .I(N__24291));
    Span4Mux_h I__3224 (
            .O(N__24291),
            .I(N__24287));
    CascadeMux I__3223 (
            .O(N__24290),
            .I(N__24284));
    Span4Mux_h I__3222 (
            .O(N__24287),
            .I(N__24280));
    InMux I__3221 (
            .O(N__24284),
            .I(N__24277));
    InMux I__3220 (
            .O(N__24283),
            .I(N__24274));
    Span4Mux_h I__3219 (
            .O(N__24280),
            .I(N__24271));
    LocalMux I__3218 (
            .O(N__24277),
            .I(buf_adcdata_iac_2));
    LocalMux I__3217 (
            .O(N__24274),
            .I(buf_adcdata_iac_2));
    Odrv4 I__3216 (
            .O(N__24271),
            .I(buf_adcdata_iac_2));
    InMux I__3215 (
            .O(N__24264),
            .I(N__24261));
    LocalMux I__3214 (
            .O(N__24261),
            .I(N__24258));
    Span4Mux_h I__3213 (
            .O(N__24258),
            .I(N__24254));
    InMux I__3212 (
            .O(N__24257),
            .I(N__24250));
    Span4Mux_v I__3211 (
            .O(N__24254),
            .I(N__24247));
    InMux I__3210 (
            .O(N__24253),
            .I(N__24244));
    LocalMux I__3209 (
            .O(N__24250),
            .I(buf_adcdata_vac_5));
    Odrv4 I__3208 (
            .O(N__24247),
            .I(buf_adcdata_vac_5));
    LocalMux I__3207 (
            .O(N__24244),
            .I(buf_adcdata_vac_5));
    InMux I__3206 (
            .O(N__24237),
            .I(N__24234));
    LocalMux I__3205 (
            .O(N__24234),
            .I(N__24231));
    Span4Mux_h I__3204 (
            .O(N__24231),
            .I(N__24228));
    Span4Mux_h I__3203 (
            .O(N__24228),
            .I(N__24223));
    InMux I__3202 (
            .O(N__24227),
            .I(N__24218));
    InMux I__3201 (
            .O(N__24226),
            .I(N__24218));
    Odrv4 I__3200 (
            .O(N__24223),
            .I(buf_adcdata_iac_5));
    LocalMux I__3199 (
            .O(N__24218),
            .I(buf_adcdata_iac_5));
    CascadeMux I__3198 (
            .O(N__24213),
            .I(n19_adj_1603_cascade_));
    CascadeMux I__3197 (
            .O(N__24210),
            .I(n22377_cascade_));
    InMux I__3196 (
            .O(N__24207),
            .I(N__24204));
    LocalMux I__3195 (
            .O(N__24204),
            .I(n21237));
    InMux I__3194 (
            .O(N__24201),
            .I(\ADC_VDC.n19869 ));
    InMux I__3193 (
            .O(N__24198),
            .I(N__24195));
    LocalMux I__3192 (
            .O(N__24195),
            .I(N__24192));
    Span4Mux_v I__3191 (
            .O(N__24192),
            .I(N__24188));
    InMux I__3190 (
            .O(N__24191),
            .I(N__24185));
    Odrv4 I__3189 (
            .O(N__24188),
            .I(cmd_rdadcbuf_29));
    LocalMux I__3188 (
            .O(N__24185),
            .I(cmd_rdadcbuf_29));
    InMux I__3187 (
            .O(N__24180),
            .I(\ADC_VDC.n19870 ));
    InMux I__3186 (
            .O(N__24177),
            .I(\ADC_VDC.n19871 ));
    InMux I__3185 (
            .O(N__24174),
            .I(\ADC_VDC.n19872 ));
    InMux I__3184 (
            .O(N__24171),
            .I(bfn_8_10_0_));
    InMux I__3183 (
            .O(N__24168),
            .I(\ADC_VDC.n19874 ));
    InMux I__3182 (
            .O(N__24165),
            .I(\ADC_VDC.n19875 ));
    InMux I__3181 (
            .O(N__24162),
            .I(N__24159));
    LocalMux I__3180 (
            .O(N__24159),
            .I(N__24156));
    Sp12to4 I__3179 (
            .O(N__24156),
            .I(N__24152));
    CascadeMux I__3178 (
            .O(N__24155),
            .I(N__24149));
    Span12Mux_v I__3177 (
            .O(N__24152),
            .I(N__24146));
    InMux I__3176 (
            .O(N__24149),
            .I(N__24143));
    Odrv12 I__3175 (
            .O(N__24146),
            .I(buf_adcdata_vdc_18));
    LocalMux I__3174 (
            .O(N__24143),
            .I(buf_adcdata_vdc_18));
    InMux I__3173 (
            .O(N__24138),
            .I(N__24135));
    LocalMux I__3172 (
            .O(N__24135),
            .I(N__24132));
    Sp12to4 I__3171 (
            .O(N__24132),
            .I(N__24127));
    InMux I__3170 (
            .O(N__24131),
            .I(N__24124));
    CascadeMux I__3169 (
            .O(N__24130),
            .I(N__24121));
    Span12Mux_v I__3168 (
            .O(N__24127),
            .I(N__24118));
    LocalMux I__3167 (
            .O(N__24124),
            .I(N__24115));
    InMux I__3166 (
            .O(N__24121),
            .I(N__24112));
    Span12Mux_h I__3165 (
            .O(N__24118),
            .I(N__24109));
    Span4Mux_h I__3164 (
            .O(N__24115),
            .I(N__24106));
    LocalMux I__3163 (
            .O(N__24112),
            .I(buf_adcdata_vac_18));
    Odrv12 I__3162 (
            .O(N__24109),
            .I(buf_adcdata_vac_18));
    Odrv4 I__3161 (
            .O(N__24106),
            .I(buf_adcdata_vac_18));
    InMux I__3160 (
            .O(N__24099),
            .I(N__24096));
    LocalMux I__3159 (
            .O(N__24096),
            .I(n19_adj_1692));
    InMux I__3158 (
            .O(N__24093),
            .I(\ADC_VDC.n19860 ));
    InMux I__3157 (
            .O(N__24090),
            .I(\ADC_VDC.n19861 ));
    InMux I__3156 (
            .O(N__24087),
            .I(\ADC_VDC.n19862 ));
    InMux I__3155 (
            .O(N__24084),
            .I(\ADC_VDC.n19863 ));
    InMux I__3154 (
            .O(N__24081),
            .I(\ADC_VDC.n19864 ));
    InMux I__3153 (
            .O(N__24078),
            .I(bfn_8_9_0_));
    InMux I__3152 (
            .O(N__24075),
            .I(\ADC_VDC.n19866 ));
    InMux I__3151 (
            .O(N__24072),
            .I(\ADC_VDC.n19867 ));
    InMux I__3150 (
            .O(N__24069),
            .I(\ADC_VDC.n19868 ));
    InMux I__3149 (
            .O(N__24066),
            .I(\ADC_VDC.n19852 ));
    InMux I__3148 (
            .O(N__24063),
            .I(\ADC_VDC.n19853 ));
    InMux I__3147 (
            .O(N__24060),
            .I(\ADC_VDC.n19854 ));
    InMux I__3146 (
            .O(N__24057),
            .I(N__24054));
    LocalMux I__3145 (
            .O(N__24054),
            .I(N__24051));
    Span4Mux_h I__3144 (
            .O(N__24051),
            .I(N__24047));
    InMux I__3143 (
            .O(N__24050),
            .I(N__24044));
    Odrv4 I__3142 (
            .O(N__24047),
            .I(cmd_rdadcbuf_14));
    LocalMux I__3141 (
            .O(N__24044),
            .I(cmd_rdadcbuf_14));
    InMux I__3140 (
            .O(N__24039),
            .I(\ADC_VDC.n19855 ));
    InMux I__3139 (
            .O(N__24036),
            .I(\ADC_VDC.n19856 ));
    CascadeMux I__3138 (
            .O(N__24033),
            .I(N__24030));
    InMux I__3137 (
            .O(N__24030),
            .I(N__24025));
    InMux I__3136 (
            .O(N__24029),
            .I(N__24020));
    InMux I__3135 (
            .O(N__24028),
            .I(N__24020));
    LocalMux I__3134 (
            .O(N__24025),
            .I(N__24017));
    LocalMux I__3133 (
            .O(N__24020),
            .I(cmd_rdadctmp_16_adj_1507));
    Odrv12 I__3132 (
            .O(N__24017),
            .I(cmd_rdadctmp_16_adj_1507));
    InMux I__3131 (
            .O(N__24012),
            .I(bfn_8_8_0_));
    CascadeMux I__3130 (
            .O(N__24009),
            .I(N__24006));
    InMux I__3129 (
            .O(N__24006),
            .I(N__24001));
    InMux I__3128 (
            .O(N__24005),
            .I(N__23996));
    InMux I__3127 (
            .O(N__24004),
            .I(N__23996));
    LocalMux I__3126 (
            .O(N__24001),
            .I(N__23993));
    LocalMux I__3125 (
            .O(N__23996),
            .I(cmd_rdadctmp_17_adj_1506));
    Odrv12 I__3124 (
            .O(N__23993),
            .I(cmd_rdadctmp_17_adj_1506));
    InMux I__3123 (
            .O(N__23988),
            .I(\ADC_VDC.n19858 ));
    CascadeMux I__3122 (
            .O(N__23985),
            .I(N__23982));
    InMux I__3121 (
            .O(N__23982),
            .I(N__23978));
    CascadeMux I__3120 (
            .O(N__23981),
            .I(N__23975));
    LocalMux I__3119 (
            .O(N__23978),
            .I(N__23971));
    InMux I__3118 (
            .O(N__23975),
            .I(N__23968));
    InMux I__3117 (
            .O(N__23974),
            .I(N__23965));
    Span4Mux_v I__3116 (
            .O(N__23971),
            .I(N__23962));
    LocalMux I__3115 (
            .O(N__23968),
            .I(cmd_rdadctmp_18_adj_1505));
    LocalMux I__3114 (
            .O(N__23965),
            .I(cmd_rdadctmp_18_adj_1505));
    Odrv4 I__3113 (
            .O(N__23962),
            .I(cmd_rdadctmp_18_adj_1505));
    InMux I__3112 (
            .O(N__23955),
            .I(\ADC_VDC.n19859 ));
    InMux I__3111 (
            .O(N__23952),
            .I(N__23949));
    LocalMux I__3110 (
            .O(N__23949),
            .I(\ADC_VDC.cmd_rdadcbuf_2 ));
    InMux I__3109 (
            .O(N__23946),
            .I(\ADC_VDC.n19843 ));
    InMux I__3108 (
            .O(N__23943),
            .I(N__23940));
    LocalMux I__3107 (
            .O(N__23940),
            .I(\ADC_VDC.cmd_rdadcbuf_3 ));
    InMux I__3106 (
            .O(N__23937),
            .I(\ADC_VDC.n19844 ));
    CascadeMux I__3105 (
            .O(N__23934),
            .I(N__23931));
    InMux I__3104 (
            .O(N__23931),
            .I(N__23928));
    LocalMux I__3103 (
            .O(N__23928),
            .I(N__23925));
    Odrv4 I__3102 (
            .O(N__23925),
            .I(\ADC_VDC.cmd_rdadcbuf_4 ));
    InMux I__3101 (
            .O(N__23922),
            .I(\ADC_VDC.n19845 ));
    InMux I__3100 (
            .O(N__23919),
            .I(N__23916));
    LocalMux I__3099 (
            .O(N__23916),
            .I(\ADC_VDC.cmd_rdadcbuf_5 ));
    InMux I__3098 (
            .O(N__23913),
            .I(\ADC_VDC.n19846 ));
    CascadeMux I__3097 (
            .O(N__23910),
            .I(N__23906));
    CascadeMux I__3096 (
            .O(N__23909),
            .I(N__23903));
    InMux I__3095 (
            .O(N__23906),
            .I(N__23899));
    InMux I__3094 (
            .O(N__23903),
            .I(N__23896));
    InMux I__3093 (
            .O(N__23902),
            .I(N__23893));
    LocalMux I__3092 (
            .O(N__23899),
            .I(N__23890));
    LocalMux I__3091 (
            .O(N__23896),
            .I(cmd_rdadctmp_6_adj_1517));
    LocalMux I__3090 (
            .O(N__23893),
            .I(cmd_rdadctmp_6_adj_1517));
    Odrv4 I__3089 (
            .O(N__23890),
            .I(cmd_rdadctmp_6_adj_1517));
    InMux I__3088 (
            .O(N__23883),
            .I(N__23880));
    LocalMux I__3087 (
            .O(N__23880),
            .I(\ADC_VDC.cmd_rdadcbuf_6 ));
    InMux I__3086 (
            .O(N__23877),
            .I(\ADC_VDC.n19847 ));
    CascadeMux I__3085 (
            .O(N__23874),
            .I(N__23871));
    InMux I__3084 (
            .O(N__23871),
            .I(N__23868));
    LocalMux I__3083 (
            .O(N__23868),
            .I(\ADC_VDC.cmd_rdadcbuf_7 ));
    InMux I__3082 (
            .O(N__23865),
            .I(\ADC_VDC.n19848 ));
    InMux I__3081 (
            .O(N__23862),
            .I(N__23859));
    LocalMux I__3080 (
            .O(N__23859),
            .I(\ADC_VDC.cmd_rdadcbuf_8 ));
    InMux I__3079 (
            .O(N__23856),
            .I(bfn_8_7_0_));
    InMux I__3078 (
            .O(N__23853),
            .I(N__23850));
    LocalMux I__3077 (
            .O(N__23850),
            .I(\ADC_VDC.cmd_rdadcbuf_9 ));
    InMux I__3076 (
            .O(N__23847),
            .I(\ADC_VDC.n19850 ));
    InMux I__3075 (
            .O(N__23844),
            .I(N__23841));
    LocalMux I__3074 (
            .O(N__23841),
            .I(\ADC_VDC.cmd_rdadcbuf_10 ));
    InMux I__3073 (
            .O(N__23838),
            .I(\ADC_VDC.n19851 ));
    CascadeMux I__3072 (
            .O(N__23835),
            .I(N__23832));
    InMux I__3071 (
            .O(N__23832),
            .I(N__23827));
    InMux I__3070 (
            .O(N__23831),
            .I(N__23822));
    InMux I__3069 (
            .O(N__23830),
            .I(N__23822));
    LocalMux I__3068 (
            .O(N__23827),
            .I(N__23819));
    LocalMux I__3067 (
            .O(N__23822),
            .I(cmd_rdadctmp_0_adj_1523));
    Odrv4 I__3066 (
            .O(N__23819),
            .I(cmd_rdadctmp_0_adj_1523));
    InMux I__3065 (
            .O(N__23814),
            .I(N__23811));
    LocalMux I__3064 (
            .O(N__23811),
            .I(\ADC_VDC.cmd_rdadcbuf_0 ));
    InMux I__3063 (
            .O(N__23808),
            .I(N__23805));
    LocalMux I__3062 (
            .O(N__23805),
            .I(\ADC_VDC.cmd_rdadcbuf_1 ));
    InMux I__3061 (
            .O(N__23802),
            .I(\ADC_VDC.n19842 ));
    InMux I__3060 (
            .O(N__23799),
            .I(N__23796));
    LocalMux I__3059 (
            .O(N__23796),
            .I(n21082));
    CascadeMux I__3058 (
            .O(N__23793),
            .I(n21082_cascade_));
    InMux I__3057 (
            .O(N__23790),
            .I(N__23784));
    InMux I__3056 (
            .O(N__23789),
            .I(N__23784));
    LocalMux I__3055 (
            .O(N__23784),
            .I(cmd_rdadctmp_3));
    CascadeMux I__3054 (
            .O(N__23781),
            .I(n12771_cascade_));
    CascadeMux I__3053 (
            .O(N__23778),
            .I(N__23775));
    InMux I__3052 (
            .O(N__23775),
            .I(N__23769));
    InMux I__3051 (
            .O(N__23774),
            .I(N__23769));
    LocalMux I__3050 (
            .O(N__23769),
            .I(cmd_rdadctmp_4));
    InMux I__3049 (
            .O(N__23766),
            .I(N__23760));
    InMux I__3048 (
            .O(N__23765),
            .I(N__23760));
    LocalMux I__3047 (
            .O(N__23760),
            .I(cmd_rdadctmp_5));
    InMux I__3046 (
            .O(N__23757),
            .I(N__23754));
    LocalMux I__3045 (
            .O(N__23754),
            .I(\ADC_IAC.n17 ));
    IoInMux I__3044 (
            .O(N__23751),
            .I(N__23748));
    LocalMux I__3043 (
            .O(N__23748),
            .I(N__23745));
    Span4Mux_s2_v I__3042 (
            .O(N__23745),
            .I(N__23742));
    Span4Mux_v I__3041 (
            .O(N__23742),
            .I(N__23739));
    Span4Mux_h I__3040 (
            .O(N__23739),
            .I(N__23736));
    Odrv4 I__3039 (
            .O(N__23736),
            .I(DDS_MCLK1));
    InMux I__3038 (
            .O(N__23733),
            .I(N__23730));
    LocalMux I__3037 (
            .O(N__23730),
            .I(N__23727));
    Span4Mux_v I__3036 (
            .O(N__23727),
            .I(N__23724));
    Span4Mux_v I__3035 (
            .O(N__23724),
            .I(N__23720));
    CascadeMux I__3034 (
            .O(N__23723),
            .I(N__23717));
    Span4Mux_h I__3033 (
            .O(N__23720),
            .I(N__23714));
    InMux I__3032 (
            .O(N__23717),
            .I(N__23711));
    Odrv4 I__3031 (
            .O(N__23714),
            .I(buf_readRTD_7));
    LocalMux I__3030 (
            .O(N__23711),
            .I(buf_readRTD_7));
    InMux I__3029 (
            .O(N__23706),
            .I(N__23703));
    LocalMux I__3028 (
            .O(N__23703),
            .I(N__23700));
    Odrv12 I__3027 (
            .O(N__23700),
            .I(n16_adj_1690));
    CascadeMux I__3026 (
            .O(N__23697),
            .I(N__23694));
    InMux I__3025 (
            .O(N__23694),
            .I(N__23691));
    LocalMux I__3024 (
            .O(N__23691),
            .I(N__23688));
    Span4Mux_v I__3023 (
            .O(N__23688),
            .I(N__23685));
    Odrv4 I__3022 (
            .O(N__23685),
            .I(n17_adj_1691));
    CEMux I__3021 (
            .O(N__23682),
            .I(N__23679));
    LocalMux I__3020 (
            .O(N__23679),
            .I(N__23676));
    Odrv4 I__3019 (
            .O(N__23676),
            .I(\ADC_IAC.n12 ));
    InMux I__3018 (
            .O(N__23673),
            .I(N__23670));
    LocalMux I__3017 (
            .O(N__23670),
            .I(\ADC_IAC.n21457 ));
    CascadeMux I__3016 (
            .O(N__23667),
            .I(N__23664));
    InMux I__3015 (
            .O(N__23664),
            .I(N__23661));
    LocalMux I__3014 (
            .O(N__23661),
            .I(N__23658));
    Span4Mux_v I__3013 (
            .O(N__23658),
            .I(N__23654));
    InMux I__3012 (
            .O(N__23657),
            .I(N__23651));
    Odrv4 I__3011 (
            .O(N__23654),
            .I(cmd_rdadctmp_7));
    LocalMux I__3010 (
            .O(N__23651),
            .I(cmd_rdadctmp_7));
    CascadeMux I__3009 (
            .O(N__23646),
            .I(N__23643));
    InMux I__3008 (
            .O(N__23643),
            .I(N__23637));
    InMux I__3007 (
            .O(N__23642),
            .I(N__23637));
    LocalMux I__3006 (
            .O(N__23637),
            .I(cmd_rdadctmp_6));
    CascadeMux I__3005 (
            .O(N__23634),
            .I(N__23631));
    InMux I__3004 (
            .O(N__23631),
            .I(N__23628));
    LocalMux I__3003 (
            .O(N__23628),
            .I(\CLK_DDS.tmp_buf_10 ));
    CascadeMux I__3002 (
            .O(N__23625),
            .I(N__23622));
    InMux I__3001 (
            .O(N__23622),
            .I(N__23619));
    LocalMux I__3000 (
            .O(N__23619),
            .I(\CLK_DDS.tmp_buf_11 ));
    InMux I__2999 (
            .O(N__23616),
            .I(N__23613));
    LocalMux I__2998 (
            .O(N__23613),
            .I(N__23610));
    Odrv4 I__2997 (
            .O(N__23610),
            .I(\CLK_DDS.tmp_buf_12 ));
    CascadeMux I__2996 (
            .O(N__23607),
            .I(N__23604));
    InMux I__2995 (
            .O(N__23604),
            .I(N__23601));
    LocalMux I__2994 (
            .O(N__23601),
            .I(N__23598));
    Odrv4 I__2993 (
            .O(N__23598),
            .I(\CLK_DDS.tmp_buf_13 ));
    CascadeMux I__2992 (
            .O(N__23595),
            .I(N__23592));
    InMux I__2991 (
            .O(N__23592),
            .I(N__23589));
    LocalMux I__2990 (
            .O(N__23589),
            .I(\CLK_DDS.tmp_buf_14 ));
    CascadeMux I__2989 (
            .O(N__23586),
            .I(N__23583));
    InMux I__2988 (
            .O(N__23583),
            .I(N__23580));
    LocalMux I__2987 (
            .O(N__23580),
            .I(\CLK_DDS.tmp_buf_9 ));
    CascadeMux I__2986 (
            .O(N__23577),
            .I(N__23574));
    InMux I__2985 (
            .O(N__23574),
            .I(N__23571));
    LocalMux I__2984 (
            .O(N__23571),
            .I(\CLK_DDS.tmp_buf_8 ));
    InMux I__2983 (
            .O(N__23568),
            .I(N__23565));
    LocalMux I__2982 (
            .O(N__23565),
            .I(N__23562));
    Span12Mux_v I__2981 (
            .O(N__23562),
            .I(N__23557));
    InMux I__2980 (
            .O(N__23561),
            .I(N__23554));
    InMux I__2979 (
            .O(N__23560),
            .I(N__23551));
    Span12Mux_h I__2978 (
            .O(N__23557),
            .I(N__23548));
    LocalMux I__2977 (
            .O(N__23554),
            .I(N__23545));
    LocalMux I__2976 (
            .O(N__23551),
            .I(buf_adcdata_vac_9));
    Odrv12 I__2975 (
            .O(N__23548),
            .I(buf_adcdata_vac_9));
    Odrv4 I__2974 (
            .O(N__23545),
            .I(buf_adcdata_vac_9));
    CascadeMux I__2973 (
            .O(N__23538),
            .I(N__23535));
    InMux I__2972 (
            .O(N__23535),
            .I(N__23531));
    CascadeMux I__2971 (
            .O(N__23534),
            .I(N__23528));
    LocalMux I__2970 (
            .O(N__23531),
            .I(N__23524));
    InMux I__2969 (
            .O(N__23528),
            .I(N__23519));
    InMux I__2968 (
            .O(N__23527),
            .I(N__23519));
    Odrv4 I__2967 (
            .O(N__23524),
            .I(cmd_rdadctmp_11));
    LocalMux I__2966 (
            .O(N__23519),
            .I(cmd_rdadctmp_11));
    CascadeMux I__2965 (
            .O(N__23514),
            .I(N__23510));
    InMux I__2964 (
            .O(N__23513),
            .I(N__23504));
    InMux I__2963 (
            .O(N__23510),
            .I(N__23504));
    InMux I__2962 (
            .O(N__23509),
            .I(N__23501));
    LocalMux I__2961 (
            .O(N__23504),
            .I(cmd_rdadctmp_12));
    LocalMux I__2960 (
            .O(N__23501),
            .I(cmd_rdadctmp_12));
    CascadeMux I__2959 (
            .O(N__23496),
            .I(N__23493));
    InMux I__2958 (
            .O(N__23493),
            .I(N__23490));
    LocalMux I__2957 (
            .O(N__23490),
            .I(N__23486));
    CascadeMux I__2956 (
            .O(N__23489),
            .I(N__23483));
    Span4Mux_h I__2955 (
            .O(N__23486),
            .I(N__23479));
    InMux I__2954 (
            .O(N__23483),
            .I(N__23476));
    InMux I__2953 (
            .O(N__23482),
            .I(N__23473));
    Odrv4 I__2952 (
            .O(N__23479),
            .I(cmd_rdadctmp_8));
    LocalMux I__2951 (
            .O(N__23476),
            .I(cmd_rdadctmp_8));
    LocalMux I__2950 (
            .O(N__23473),
            .I(cmd_rdadctmp_8));
    CascadeMux I__2949 (
            .O(N__23466),
            .I(N__23462));
    InMux I__2948 (
            .O(N__23465),
            .I(N__23458));
    InMux I__2947 (
            .O(N__23462),
            .I(N__23453));
    InMux I__2946 (
            .O(N__23461),
            .I(N__23453));
    LocalMux I__2945 (
            .O(N__23458),
            .I(cmd_rdadctmp_17_adj_1475));
    LocalMux I__2944 (
            .O(N__23453),
            .I(cmd_rdadctmp_17_adj_1475));
    CascadeMux I__2943 (
            .O(N__23448),
            .I(N__23444));
    InMux I__2942 (
            .O(N__23447),
            .I(N__23438));
    InMux I__2941 (
            .O(N__23444),
            .I(N__23438));
    CascadeMux I__2940 (
            .O(N__23443),
            .I(N__23435));
    LocalMux I__2939 (
            .O(N__23438),
            .I(N__23432));
    InMux I__2938 (
            .O(N__23435),
            .I(N__23429));
    Odrv4 I__2937 (
            .O(N__23432),
            .I(cmd_rdadctmp_29_adj_1463));
    LocalMux I__2936 (
            .O(N__23429),
            .I(cmd_rdadctmp_29_adj_1463));
    CascadeMux I__2935 (
            .O(N__23424),
            .I(N__23420));
    CascadeMux I__2934 (
            .O(N__23423),
            .I(N__23417));
    InMux I__2933 (
            .O(N__23420),
            .I(N__23413));
    InMux I__2932 (
            .O(N__23417),
            .I(N__23408));
    InMux I__2931 (
            .O(N__23416),
            .I(N__23408));
    LocalMux I__2930 (
            .O(N__23413),
            .I(cmd_rdadctmp_9_adj_1483));
    LocalMux I__2929 (
            .O(N__23408),
            .I(cmd_rdadctmp_9_adj_1483));
    InMux I__2928 (
            .O(N__23403),
            .I(N__23400));
    LocalMux I__2927 (
            .O(N__23400),
            .I(N__23397));
    Span4Mux_v I__2926 (
            .O(N__23397),
            .I(N__23394));
    Span4Mux_h I__2925 (
            .O(N__23394),
            .I(N__23391));
    Odrv4 I__2924 (
            .O(N__23391),
            .I(buf_data_iac_6));
    InMux I__2923 (
            .O(N__23388),
            .I(N__23385));
    LocalMux I__2922 (
            .O(N__23385),
            .I(N__23382));
    Odrv4 I__2921 (
            .O(N__23382),
            .I(n22_adj_1601));
    InMux I__2920 (
            .O(N__23379),
            .I(N__23376));
    LocalMux I__2919 (
            .O(N__23376),
            .I(N__23373));
    Span4Mux_v I__2918 (
            .O(N__23373),
            .I(N__23370));
    Span4Mux_v I__2917 (
            .O(N__23370),
            .I(N__23367));
    Sp12to4 I__2916 (
            .O(N__23367),
            .I(N__23364));
    Span12Mux_h I__2915 (
            .O(N__23364),
            .I(N__23361));
    Odrv12 I__2914 (
            .O(N__23361),
            .I(buf_data_iac_2));
    InMux I__2913 (
            .O(N__23358),
            .I(N__23355));
    LocalMux I__2912 (
            .O(N__23355),
            .I(n22_adj_1613));
    InMux I__2911 (
            .O(N__23352),
            .I(N__23349));
    LocalMux I__2910 (
            .O(N__23349),
            .I(N__23345));
    InMux I__2909 (
            .O(N__23348),
            .I(N__23342));
    Span4Mux_h I__2908 (
            .O(N__23345),
            .I(N__23337));
    LocalMux I__2907 (
            .O(N__23342),
            .I(N__23337));
    Odrv4 I__2906 (
            .O(N__23337),
            .I(buf_readRTD_10));
    CascadeMux I__2905 (
            .O(N__23334),
            .I(N__23331));
    InMux I__2904 (
            .O(N__23331),
            .I(N__23327));
    CascadeMux I__2903 (
            .O(N__23330),
            .I(N__23324));
    LocalMux I__2902 (
            .O(N__23327),
            .I(N__23320));
    InMux I__2901 (
            .O(N__23324),
            .I(N__23315));
    InMux I__2900 (
            .O(N__23323),
            .I(N__23315));
    Span4Mux_h I__2899 (
            .O(N__23320),
            .I(N__23308));
    LocalMux I__2898 (
            .O(N__23315),
            .I(N__23308));
    InMux I__2897 (
            .O(N__23314),
            .I(N__23303));
    InMux I__2896 (
            .O(N__23313),
            .I(N__23303));
    Odrv4 I__2895 (
            .O(N__23308),
            .I(buf_cfgRTD_2));
    LocalMux I__2894 (
            .O(N__23303),
            .I(buf_cfgRTD_2));
    CascadeMux I__2893 (
            .O(N__23298),
            .I(N__23294));
    CascadeMux I__2892 (
            .O(N__23297),
            .I(N__23291));
    InMux I__2891 (
            .O(N__23294),
            .I(N__23288));
    InMux I__2890 (
            .O(N__23291),
            .I(N__23285));
    LocalMux I__2889 (
            .O(N__23288),
            .I(N__23281));
    LocalMux I__2888 (
            .O(N__23285),
            .I(N__23278));
    InMux I__2887 (
            .O(N__23284),
            .I(N__23275));
    Odrv12 I__2886 (
            .O(N__23281),
            .I(cmd_rdadctmp_11_adj_1481));
    Odrv4 I__2885 (
            .O(N__23278),
            .I(cmd_rdadctmp_11_adj_1481));
    LocalMux I__2884 (
            .O(N__23275),
            .I(cmd_rdadctmp_11_adj_1481));
    InMux I__2883 (
            .O(N__23268),
            .I(N__23265));
    LocalMux I__2882 (
            .O(N__23265),
            .I(N__23262));
    Span4Mux_v I__2881 (
            .O(N__23262),
            .I(N__23259));
    Sp12to4 I__2880 (
            .O(N__23259),
            .I(N__23254));
    InMux I__2879 (
            .O(N__23258),
            .I(N__23251));
    InMux I__2878 (
            .O(N__23257),
            .I(N__23248));
    Span12Mux_h I__2877 (
            .O(N__23254),
            .I(N__23245));
    LocalMux I__2876 (
            .O(N__23251),
            .I(N__23242));
    LocalMux I__2875 (
            .O(N__23248),
            .I(buf_adcdata_vac_3));
    Odrv12 I__2874 (
            .O(N__23245),
            .I(buf_adcdata_vac_3));
    Odrv4 I__2873 (
            .O(N__23242),
            .I(buf_adcdata_vac_3));
    CascadeMux I__2872 (
            .O(N__23235),
            .I(N__23232));
    InMux I__2871 (
            .O(N__23232),
            .I(N__23229));
    LocalMux I__2870 (
            .O(N__23229),
            .I(N__23224));
    CascadeMux I__2869 (
            .O(N__23228),
            .I(N__23221));
    CascadeMux I__2868 (
            .O(N__23227),
            .I(N__23218));
    Span4Mux_v I__2867 (
            .O(N__23224),
            .I(N__23215));
    InMux I__2866 (
            .O(N__23221),
            .I(N__23212));
    InMux I__2865 (
            .O(N__23218),
            .I(N__23209));
    Odrv4 I__2864 (
            .O(N__23215),
            .I(cmd_rdadctmp_13_adj_1479));
    LocalMux I__2863 (
            .O(N__23212),
            .I(cmd_rdadctmp_13_adj_1479));
    LocalMux I__2862 (
            .O(N__23209),
            .I(cmd_rdadctmp_13_adj_1479));
    InMux I__2861 (
            .O(N__23202),
            .I(N__23197));
    InMux I__2860 (
            .O(N__23201),
            .I(N__23194));
    InMux I__2859 (
            .O(N__23200),
            .I(N__23191));
    LocalMux I__2858 (
            .O(N__23197),
            .I(cmd_rdadctmp_30_adj_1462));
    LocalMux I__2857 (
            .O(N__23194),
            .I(cmd_rdadctmp_30_adj_1462));
    LocalMux I__2856 (
            .O(N__23191),
            .I(cmd_rdadctmp_30_adj_1462));
    CascadeMux I__2855 (
            .O(N__23184),
            .I(N__23181));
    InMux I__2854 (
            .O(N__23181),
            .I(N__23178));
    LocalMux I__2853 (
            .O(N__23178),
            .I(n20_adj_1693));
    InMux I__2852 (
            .O(N__23175),
            .I(N__23172));
    LocalMux I__2851 (
            .O(N__23172),
            .I(n22407));
    InMux I__2850 (
            .O(N__23169),
            .I(N__23166));
    LocalMux I__2849 (
            .O(N__23166),
            .I(N__23163));
    Span12Mux_s9_h I__2848 (
            .O(N__23163),
            .I(N__23160));
    Span12Mux_h I__2847 (
            .O(N__23160),
            .I(N__23155));
    InMux I__2846 (
            .O(N__23159),
            .I(N__23150));
    InMux I__2845 (
            .O(N__23158),
            .I(N__23150));
    Odrv12 I__2844 (
            .O(N__23155),
            .I(buf_adcdata_vac_2));
    LocalMux I__2843 (
            .O(N__23150),
            .I(buf_adcdata_vac_2));
    CascadeMux I__2842 (
            .O(N__23145),
            .I(n19_adj_1612_cascade_));
    InMux I__2841 (
            .O(N__23142),
            .I(N__23139));
    LocalMux I__2840 (
            .O(N__23139),
            .I(N__23134));
    InMux I__2839 (
            .O(N__23138),
            .I(N__23131));
    InMux I__2838 (
            .O(N__23137),
            .I(N__23128));
    Span4Mux_h I__2837 (
            .O(N__23134),
            .I(N__23125));
    LocalMux I__2836 (
            .O(N__23131),
            .I(N__23122));
    LocalMux I__2835 (
            .O(N__23128),
            .I(N__23117));
    Span4Mux_v I__2834 (
            .O(N__23125),
            .I(N__23117));
    Span4Mux_h I__2833 (
            .O(N__23122),
            .I(N__23114));
    Odrv4 I__2832 (
            .O(N__23117),
            .I(buf_adcdata_vac_6));
    Odrv4 I__2831 (
            .O(N__23114),
            .I(buf_adcdata_vac_6));
    InMux I__2830 (
            .O(N__23109),
            .I(N__23106));
    LocalMux I__2829 (
            .O(N__23106),
            .I(N__23103));
    Span4Mux_h I__2828 (
            .O(N__23103),
            .I(N__23100));
    Span4Mux_v I__2827 (
            .O(N__23100),
            .I(N__23096));
    CascadeMux I__2826 (
            .O(N__23099),
            .I(N__23093));
    Sp12to4 I__2825 (
            .O(N__23096),
            .I(N__23089));
    InMux I__2824 (
            .O(N__23093),
            .I(N__23086));
    InMux I__2823 (
            .O(N__23092),
            .I(N__23083));
    Span12Mux_h I__2822 (
            .O(N__23089),
            .I(N__23080));
    LocalMux I__2821 (
            .O(N__23086),
            .I(buf_adcdata_vac_22));
    LocalMux I__2820 (
            .O(N__23083),
            .I(buf_adcdata_vac_22));
    Odrv12 I__2819 (
            .O(N__23080),
            .I(buf_adcdata_vac_22));
    InMux I__2818 (
            .O(N__23073),
            .I(N__23070));
    LocalMux I__2817 (
            .O(N__23070),
            .I(N__23067));
    Odrv4 I__2816 (
            .O(N__23067),
            .I(n22629));
    CascadeMux I__2815 (
            .O(N__23064),
            .I(N__23061));
    InMux I__2814 (
            .O(N__23061),
            .I(N__23057));
    CascadeMux I__2813 (
            .O(N__23060),
            .I(N__23054));
    LocalMux I__2812 (
            .O(N__23057),
            .I(N__23050));
    InMux I__2811 (
            .O(N__23054),
            .I(N__23047));
    InMux I__2810 (
            .O(N__23053),
            .I(N__23044));
    Odrv4 I__2809 (
            .O(N__23050),
            .I(cmd_rdadctmp_14_adj_1478));
    LocalMux I__2808 (
            .O(N__23047),
            .I(cmd_rdadctmp_14_adj_1478));
    LocalMux I__2807 (
            .O(N__23044),
            .I(cmd_rdadctmp_14_adj_1478));
    CascadeMux I__2806 (
            .O(N__23037),
            .I(N__23034));
    InMux I__2805 (
            .O(N__23034),
            .I(N__23031));
    LocalMux I__2804 (
            .O(N__23031),
            .I(N__23027));
    CascadeMux I__2803 (
            .O(N__23030),
            .I(N__23024));
    Span4Mux_v I__2802 (
            .O(N__23027),
            .I(N__23020));
    InMux I__2801 (
            .O(N__23024),
            .I(N__23015));
    InMux I__2800 (
            .O(N__23023),
            .I(N__23015));
    Odrv4 I__2799 (
            .O(N__23020),
            .I(cmd_rdadctmp_15_adj_1477));
    LocalMux I__2798 (
            .O(N__23015),
            .I(cmd_rdadctmp_15_adj_1477));
    CascadeMux I__2797 (
            .O(N__23010),
            .I(N__23002));
    CascadeMux I__2796 (
            .O(N__23009),
            .I(N__22999));
    InMux I__2795 (
            .O(N__23008),
            .I(N__22995));
    InMux I__2794 (
            .O(N__23007),
            .I(N__22992));
    InMux I__2793 (
            .O(N__23006),
            .I(N__22989));
    InMux I__2792 (
            .O(N__23005),
            .I(N__22980));
    InMux I__2791 (
            .O(N__23002),
            .I(N__22980));
    InMux I__2790 (
            .O(N__22999),
            .I(N__22980));
    InMux I__2789 (
            .O(N__22998),
            .I(N__22980));
    LocalMux I__2788 (
            .O(N__22995),
            .I(\RTD.n13090 ));
    LocalMux I__2787 (
            .O(N__22992),
            .I(\RTD.n13090 ));
    LocalMux I__2786 (
            .O(N__22989),
            .I(\RTD.n13090 ));
    LocalMux I__2785 (
            .O(N__22980),
            .I(\RTD.n13090 ));
    CascadeMux I__2784 (
            .O(N__22971),
            .I(N__22964));
    CascadeMux I__2783 (
            .O(N__22970),
            .I(N__22961));
    CascadeMux I__2782 (
            .O(N__22969),
            .I(N__22957));
    CascadeMux I__2781 (
            .O(N__22968),
            .I(N__22954));
    CascadeMux I__2780 (
            .O(N__22967),
            .I(N__22951));
    InMux I__2779 (
            .O(N__22964),
            .I(N__22945));
    InMux I__2778 (
            .O(N__22961),
            .I(N__22942));
    InMux I__2777 (
            .O(N__22960),
            .I(N__22939));
    InMux I__2776 (
            .O(N__22957),
            .I(N__22936));
    InMux I__2775 (
            .O(N__22954),
            .I(N__22925));
    InMux I__2774 (
            .O(N__22951),
            .I(N__22925));
    InMux I__2773 (
            .O(N__22950),
            .I(N__22925));
    InMux I__2772 (
            .O(N__22949),
            .I(N__22925));
    InMux I__2771 (
            .O(N__22948),
            .I(N__22925));
    LocalMux I__2770 (
            .O(N__22945),
            .I(N__22916));
    LocalMux I__2769 (
            .O(N__22942),
            .I(N__22916));
    LocalMux I__2768 (
            .O(N__22939),
            .I(N__22916));
    LocalMux I__2767 (
            .O(N__22936),
            .I(N__22916));
    LocalMux I__2766 (
            .O(N__22925),
            .I(N__22913));
    Span4Mux_h I__2765 (
            .O(N__22916),
            .I(N__22910));
    Span4Mux_h I__2764 (
            .O(N__22913),
            .I(N__22907));
    Odrv4 I__2763 (
            .O(N__22910),
            .I(\RTD.n21061 ));
    Odrv4 I__2762 (
            .O(N__22907),
            .I(\RTD.n21061 ));
    InMux I__2761 (
            .O(N__22902),
            .I(N__22898));
    InMux I__2760 (
            .O(N__22901),
            .I(N__22895));
    LocalMux I__2759 (
            .O(N__22898),
            .I(N__22892));
    LocalMux I__2758 (
            .O(N__22895),
            .I(\RTD.cfg_buf_0 ));
    Odrv4 I__2757 (
            .O(N__22892),
            .I(\RTD.cfg_buf_0 ));
    InMux I__2756 (
            .O(N__22887),
            .I(N__22883));
    InMux I__2755 (
            .O(N__22886),
            .I(N__22880));
    LocalMux I__2754 (
            .O(N__22883),
            .I(buf_readRTD_9));
    LocalMux I__2753 (
            .O(N__22880),
            .I(buf_readRTD_9));
    InMux I__2752 (
            .O(N__22875),
            .I(N__22871));
    CascadeMux I__2751 (
            .O(N__22874),
            .I(N__22868));
    LocalMux I__2750 (
            .O(N__22871),
            .I(N__22865));
    InMux I__2749 (
            .O(N__22868),
            .I(N__22862));
    Odrv12 I__2748 (
            .O(N__22865),
            .I(buf_adcdata_vdc_3));
    LocalMux I__2747 (
            .O(N__22862),
            .I(buf_adcdata_vdc_3));
    InMux I__2746 (
            .O(N__22857),
            .I(N__22854));
    LocalMux I__2745 (
            .O(N__22854),
            .I(N__22850));
    InMux I__2744 (
            .O(N__22853),
            .I(N__22847));
    Span12Mux_v I__2743 (
            .O(N__22850),
            .I(N__22843));
    LocalMux I__2742 (
            .O(N__22847),
            .I(N__22840));
    InMux I__2741 (
            .O(N__22846),
            .I(N__22837));
    Span12Mux_h I__2740 (
            .O(N__22843),
            .I(N__22834));
    Span4Mux_h I__2739 (
            .O(N__22840),
            .I(N__22831));
    LocalMux I__2738 (
            .O(N__22837),
            .I(buf_adcdata_iac_3));
    Odrv12 I__2737 (
            .O(N__22834),
            .I(buf_adcdata_iac_3));
    Odrv4 I__2736 (
            .O(N__22831),
            .I(buf_adcdata_iac_3));
    CascadeMux I__2735 (
            .O(N__22824),
            .I(n19_adj_1609_cascade_));
    CascadeMux I__2734 (
            .O(N__22821),
            .I(N__22818));
    InMux I__2733 (
            .O(N__22818),
            .I(N__22815));
    LocalMux I__2732 (
            .O(N__22815),
            .I(N__22811));
    InMux I__2731 (
            .O(N__22814),
            .I(N__22808));
    Odrv12 I__2730 (
            .O(N__22811),
            .I(buf_readRTD_14));
    LocalMux I__2729 (
            .O(N__22808),
            .I(buf_readRTD_14));
    CascadeMux I__2728 (
            .O(N__22803),
            .I(N__22800));
    InMux I__2727 (
            .O(N__22800),
            .I(N__22796));
    CascadeMux I__2726 (
            .O(N__22799),
            .I(N__22793));
    LocalMux I__2725 (
            .O(N__22796),
            .I(N__22789));
    InMux I__2724 (
            .O(N__22793),
            .I(N__22786));
    InMux I__2723 (
            .O(N__22792),
            .I(N__22783));
    Span4Mux_h I__2722 (
            .O(N__22789),
            .I(N__22780));
    LocalMux I__2721 (
            .O(N__22786),
            .I(cmd_rdadctmp_10_adj_1482));
    LocalMux I__2720 (
            .O(N__22783),
            .I(cmd_rdadctmp_10_adj_1482));
    Odrv4 I__2719 (
            .O(N__22780),
            .I(cmd_rdadctmp_10_adj_1482));
    IoInMux I__2718 (
            .O(N__22773),
            .I(N__22770));
    LocalMux I__2717 (
            .O(N__22770),
            .I(N__22767));
    Span12Mux_s5_v I__2716 (
            .O(N__22767),
            .I(N__22763));
    InMux I__2715 (
            .O(N__22766),
            .I(N__22760));
    Odrv12 I__2714 (
            .O(N__22763),
            .I(DDS_MOSI1));
    LocalMux I__2713 (
            .O(N__22760),
            .I(DDS_MOSI1));
    InMux I__2712 (
            .O(N__22755),
            .I(N__22749));
    InMux I__2711 (
            .O(N__22754),
            .I(N__22749));
    LocalMux I__2710 (
            .O(N__22749),
            .I(\RTD.cfg_buf_5 ));
    InMux I__2709 (
            .O(N__22746),
            .I(N__22743));
    LocalMux I__2708 (
            .O(N__22743),
            .I(\RTD.n11_adj_1444 ));
    InMux I__2707 (
            .O(N__22740),
            .I(N__22734));
    InMux I__2706 (
            .O(N__22739),
            .I(N__22734));
    LocalMux I__2705 (
            .O(N__22734),
            .I(\RTD.cfg_buf_3 ));
    InMux I__2704 (
            .O(N__22731),
            .I(N__22725));
    InMux I__2703 (
            .O(N__22730),
            .I(N__22725));
    LocalMux I__2702 (
            .O(N__22725),
            .I(\RTD.cfg_buf_4 ));
    InMux I__2701 (
            .O(N__22722),
            .I(N__22716));
    InMux I__2700 (
            .O(N__22721),
            .I(N__22716));
    LocalMux I__2699 (
            .O(N__22716),
            .I(\RTD.cfg_buf_2 ));
    InMux I__2698 (
            .O(N__22713),
            .I(N__22710));
    LocalMux I__2697 (
            .O(N__22710),
            .I(\RTD.n10 ));
    InMux I__2696 (
            .O(N__22707),
            .I(N__22703));
    InMux I__2695 (
            .O(N__22706),
            .I(N__22700));
    LocalMux I__2694 (
            .O(N__22703),
            .I(\RTD.n11 ));
    LocalMux I__2693 (
            .O(N__22700),
            .I(\RTD.n11 ));
    CascadeMux I__2692 (
            .O(N__22695),
            .I(N__22688));
    InMux I__2691 (
            .O(N__22694),
            .I(N__22680));
    InMux I__2690 (
            .O(N__22693),
            .I(N__22674));
    CascadeMux I__2689 (
            .O(N__22692),
            .I(N__22671));
    InMux I__2688 (
            .O(N__22691),
            .I(N__22663));
    InMux I__2687 (
            .O(N__22688),
            .I(N__22663));
    InMux I__2686 (
            .O(N__22687),
            .I(N__22663));
    InMux I__2685 (
            .O(N__22686),
            .I(N__22660));
    InMux I__2684 (
            .O(N__22685),
            .I(N__22653));
    InMux I__2683 (
            .O(N__22684),
            .I(N__22653));
    InMux I__2682 (
            .O(N__22683),
            .I(N__22653));
    LocalMux I__2681 (
            .O(N__22680),
            .I(N__22649));
    InMux I__2680 (
            .O(N__22679),
            .I(N__22646));
    CascadeMux I__2679 (
            .O(N__22678),
            .I(N__22641));
    CascadeMux I__2678 (
            .O(N__22677),
            .I(N__22636));
    LocalMux I__2677 (
            .O(N__22674),
            .I(N__22632));
    InMux I__2676 (
            .O(N__22671),
            .I(N__22627));
    InMux I__2675 (
            .O(N__22670),
            .I(N__22627));
    LocalMux I__2674 (
            .O(N__22663),
            .I(N__22620));
    LocalMux I__2673 (
            .O(N__22660),
            .I(N__22620));
    LocalMux I__2672 (
            .O(N__22653),
            .I(N__22620));
    InMux I__2671 (
            .O(N__22652),
            .I(N__22617));
    Span4Mux_v I__2670 (
            .O(N__22649),
            .I(N__22614));
    LocalMux I__2669 (
            .O(N__22646),
            .I(N__22611));
    CascadeMux I__2668 (
            .O(N__22645),
            .I(N__22606));
    InMux I__2667 (
            .O(N__22644),
            .I(N__22600));
    InMux I__2666 (
            .O(N__22641),
            .I(N__22597));
    InMux I__2665 (
            .O(N__22640),
            .I(N__22594));
    InMux I__2664 (
            .O(N__22639),
            .I(N__22587));
    InMux I__2663 (
            .O(N__22636),
            .I(N__22587));
    InMux I__2662 (
            .O(N__22635),
            .I(N__22587));
    Span4Mux_v I__2661 (
            .O(N__22632),
            .I(N__22580));
    LocalMux I__2660 (
            .O(N__22627),
            .I(N__22580));
    Span4Mux_v I__2659 (
            .O(N__22620),
            .I(N__22580));
    LocalMux I__2658 (
            .O(N__22617),
            .I(N__22573));
    Span4Mux_h I__2657 (
            .O(N__22614),
            .I(N__22573));
    Span4Mux_h I__2656 (
            .O(N__22611),
            .I(N__22573));
    InMux I__2655 (
            .O(N__22610),
            .I(N__22560));
    InMux I__2654 (
            .O(N__22609),
            .I(N__22560));
    InMux I__2653 (
            .O(N__22606),
            .I(N__22560));
    InMux I__2652 (
            .O(N__22605),
            .I(N__22560));
    InMux I__2651 (
            .O(N__22604),
            .I(N__22560));
    InMux I__2650 (
            .O(N__22603),
            .I(N__22560));
    LocalMux I__2649 (
            .O(N__22600),
            .I(\RTD.adc_state_3 ));
    LocalMux I__2648 (
            .O(N__22597),
            .I(\RTD.adc_state_3 ));
    LocalMux I__2647 (
            .O(N__22594),
            .I(\RTD.adc_state_3 ));
    LocalMux I__2646 (
            .O(N__22587),
            .I(\RTD.adc_state_3 ));
    Odrv4 I__2645 (
            .O(N__22580),
            .I(\RTD.adc_state_3 ));
    Odrv4 I__2644 (
            .O(N__22573),
            .I(\RTD.adc_state_3 ));
    LocalMux I__2643 (
            .O(N__22560),
            .I(\RTD.adc_state_3 ));
    CascadeMux I__2642 (
            .O(N__22545),
            .I(N__22541));
    InMux I__2641 (
            .O(N__22544),
            .I(N__22538));
    InMux I__2640 (
            .O(N__22541),
            .I(N__22535));
    LocalMux I__2639 (
            .O(N__22538),
            .I(N__22532));
    LocalMux I__2638 (
            .O(N__22535),
            .I(\RTD.n21036 ));
    Odrv12 I__2637 (
            .O(N__22532),
            .I(\RTD.n21036 ));
    InMux I__2636 (
            .O(N__22527),
            .I(N__22523));
    InMux I__2635 (
            .O(N__22526),
            .I(N__22520));
    LocalMux I__2634 (
            .O(N__22523),
            .I(N__22517));
    LocalMux I__2633 (
            .O(N__22520),
            .I(N__22513));
    Span4Mux_v I__2632 (
            .O(N__22517),
            .I(N__22509));
    InMux I__2631 (
            .O(N__22516),
            .I(N__22506));
    Span4Mux_h I__2630 (
            .O(N__22513),
            .I(N__22503));
    InMux I__2629 (
            .O(N__22512),
            .I(N__22500));
    Odrv4 I__2628 (
            .O(N__22509),
            .I(\RTD.n21199 ));
    LocalMux I__2627 (
            .O(N__22506),
            .I(\RTD.n21199 ));
    Odrv4 I__2626 (
            .O(N__22503),
            .I(\RTD.n21199 ));
    LocalMux I__2625 (
            .O(N__22500),
            .I(\RTD.n21199 ));
    CascadeMux I__2624 (
            .O(N__22491),
            .I(\RTD.n13090_cascade_ ));
    InMux I__2623 (
            .O(N__22488),
            .I(N__22484));
    InMux I__2622 (
            .O(N__22487),
            .I(N__22481));
    LocalMux I__2621 (
            .O(N__22484),
            .I(\RTD.cfg_buf_1 ));
    LocalMux I__2620 (
            .O(N__22481),
            .I(\RTD.cfg_buf_1 ));
    InMux I__2619 (
            .O(N__22476),
            .I(N__22473));
    LocalMux I__2618 (
            .O(N__22473),
            .I(\RTD.n12 ));
    InMux I__2617 (
            .O(N__22470),
            .I(N__22464));
    InMux I__2616 (
            .O(N__22469),
            .I(N__22464));
    LocalMux I__2615 (
            .O(N__22464),
            .I(\RTD.cfg_buf_7 ));
    InMux I__2614 (
            .O(N__22461),
            .I(N__22458));
    LocalMux I__2613 (
            .O(N__22458),
            .I(\RTD.cfg_tmp_1 ));
    CascadeMux I__2612 (
            .O(N__22455),
            .I(N__22452));
    InMux I__2611 (
            .O(N__22452),
            .I(N__22449));
    LocalMux I__2610 (
            .O(N__22449),
            .I(\RTD.cfg_tmp_2 ));
    InMux I__2609 (
            .O(N__22446),
            .I(N__22443));
    LocalMux I__2608 (
            .O(N__22443),
            .I(\RTD.cfg_tmp_3 ));
    InMux I__2607 (
            .O(N__22440),
            .I(N__22437));
    LocalMux I__2606 (
            .O(N__22437),
            .I(\RTD.cfg_tmp_4 ));
    InMux I__2605 (
            .O(N__22434),
            .I(N__22431));
    LocalMux I__2604 (
            .O(N__22431),
            .I(\RTD.cfg_tmp_5 ));
    InMux I__2603 (
            .O(N__22428),
            .I(N__22425));
    LocalMux I__2602 (
            .O(N__22425),
            .I(\RTD.cfg_tmp_6 ));
    CascadeMux I__2601 (
            .O(N__22422),
            .I(N__22418));
    CascadeMux I__2600 (
            .O(N__22421),
            .I(N__22415));
    InMux I__2599 (
            .O(N__22418),
            .I(N__22406));
    InMux I__2598 (
            .O(N__22415),
            .I(N__22383));
    InMux I__2597 (
            .O(N__22414),
            .I(N__22383));
    InMux I__2596 (
            .O(N__22413),
            .I(N__22383));
    InMux I__2595 (
            .O(N__22412),
            .I(N__22383));
    InMux I__2594 (
            .O(N__22411),
            .I(N__22383));
    InMux I__2593 (
            .O(N__22410),
            .I(N__22383));
    InMux I__2592 (
            .O(N__22409),
            .I(N__22383));
    LocalMux I__2591 (
            .O(N__22406),
            .I(N__22380));
    InMux I__2590 (
            .O(N__22405),
            .I(N__22370));
    InMux I__2589 (
            .O(N__22404),
            .I(N__22370));
    InMux I__2588 (
            .O(N__22403),
            .I(N__22361));
    InMux I__2587 (
            .O(N__22402),
            .I(N__22361));
    InMux I__2586 (
            .O(N__22401),
            .I(N__22361));
    InMux I__2585 (
            .O(N__22400),
            .I(N__22361));
    InMux I__2584 (
            .O(N__22399),
            .I(N__22356));
    InMux I__2583 (
            .O(N__22398),
            .I(N__22356));
    LocalMux I__2582 (
            .O(N__22383),
            .I(N__22353));
    Span4Mux_v I__2581 (
            .O(N__22380),
            .I(N__22347));
    InMux I__2580 (
            .O(N__22379),
            .I(N__22344));
    CascadeMux I__2579 (
            .O(N__22378),
            .I(N__22333));
    CascadeMux I__2578 (
            .O(N__22377),
            .I(N__22328));
    InMux I__2577 (
            .O(N__22376),
            .I(N__22324));
    InMux I__2576 (
            .O(N__22375),
            .I(N__22321));
    LocalMux I__2575 (
            .O(N__22370),
            .I(N__22314));
    LocalMux I__2574 (
            .O(N__22361),
            .I(N__22314));
    LocalMux I__2573 (
            .O(N__22356),
            .I(N__22314));
    Span4Mux_v I__2572 (
            .O(N__22353),
            .I(N__22311));
    InMux I__2571 (
            .O(N__22352),
            .I(N__22308));
    InMux I__2570 (
            .O(N__22351),
            .I(N__22305));
    InMux I__2569 (
            .O(N__22350),
            .I(N__22302));
    Span4Mux_h I__2568 (
            .O(N__22347),
            .I(N__22297));
    LocalMux I__2567 (
            .O(N__22344),
            .I(N__22297));
    InMux I__2566 (
            .O(N__22343),
            .I(N__22284));
    InMux I__2565 (
            .O(N__22342),
            .I(N__22284));
    InMux I__2564 (
            .O(N__22341),
            .I(N__22284));
    InMux I__2563 (
            .O(N__22340),
            .I(N__22284));
    InMux I__2562 (
            .O(N__22339),
            .I(N__22284));
    InMux I__2561 (
            .O(N__22338),
            .I(N__22284));
    InMux I__2560 (
            .O(N__22337),
            .I(N__22269));
    InMux I__2559 (
            .O(N__22336),
            .I(N__22269));
    InMux I__2558 (
            .O(N__22333),
            .I(N__22269));
    InMux I__2557 (
            .O(N__22332),
            .I(N__22269));
    InMux I__2556 (
            .O(N__22331),
            .I(N__22269));
    InMux I__2555 (
            .O(N__22328),
            .I(N__22269));
    InMux I__2554 (
            .O(N__22327),
            .I(N__22269));
    LocalMux I__2553 (
            .O(N__22324),
            .I(N__22262));
    LocalMux I__2552 (
            .O(N__22321),
            .I(N__22262));
    Span4Mux_v I__2551 (
            .O(N__22314),
            .I(N__22262));
    Sp12to4 I__2550 (
            .O(N__22311),
            .I(N__22257));
    LocalMux I__2549 (
            .O(N__22308),
            .I(N__22257));
    LocalMux I__2548 (
            .O(N__22305),
            .I(\RTD.adc_state_0 ));
    LocalMux I__2547 (
            .O(N__22302),
            .I(\RTD.adc_state_0 ));
    Odrv4 I__2546 (
            .O(N__22297),
            .I(\RTD.adc_state_0 ));
    LocalMux I__2545 (
            .O(N__22284),
            .I(\RTD.adc_state_0 ));
    LocalMux I__2544 (
            .O(N__22269),
            .I(\RTD.adc_state_0 ));
    Odrv4 I__2543 (
            .O(N__22262),
            .I(\RTD.adc_state_0 ));
    Odrv12 I__2542 (
            .O(N__22257),
            .I(\RTD.adc_state_0 ));
    InMux I__2541 (
            .O(N__22242),
            .I(N__22239));
    LocalMux I__2540 (
            .O(N__22239),
            .I(N__22236));
    Span4Mux_v I__2539 (
            .O(N__22236),
            .I(N__22232));
    InMux I__2538 (
            .O(N__22235),
            .I(N__22229));
    Odrv4 I__2537 (
            .O(N__22232),
            .I(\RTD.cfg_tmp_7 ));
    LocalMux I__2536 (
            .O(N__22229),
            .I(\RTD.cfg_tmp_7 ));
    InMux I__2535 (
            .O(N__22224),
            .I(N__22198));
    InMux I__2534 (
            .O(N__22223),
            .I(N__22198));
    InMux I__2533 (
            .O(N__22222),
            .I(N__22198));
    InMux I__2532 (
            .O(N__22221),
            .I(N__22198));
    InMux I__2531 (
            .O(N__22220),
            .I(N__22198));
    InMux I__2530 (
            .O(N__22219),
            .I(N__22198));
    InMux I__2529 (
            .O(N__22218),
            .I(N__22198));
    InMux I__2528 (
            .O(N__22217),
            .I(N__22198));
    InMux I__2527 (
            .O(N__22216),
            .I(N__22189));
    CascadeMux I__2526 (
            .O(N__22215),
            .I(N__22183));
    LocalMux I__2525 (
            .O(N__22198),
            .I(N__22170));
    InMux I__2524 (
            .O(N__22197),
            .I(N__22157));
    InMux I__2523 (
            .O(N__22196),
            .I(N__22157));
    InMux I__2522 (
            .O(N__22195),
            .I(N__22157));
    InMux I__2521 (
            .O(N__22194),
            .I(N__22157));
    InMux I__2520 (
            .O(N__22193),
            .I(N__22157));
    CascadeMux I__2519 (
            .O(N__22192),
            .I(N__22149));
    LocalMux I__2518 (
            .O(N__22189),
            .I(N__22146));
    InMux I__2517 (
            .O(N__22188),
            .I(N__22141));
    InMux I__2516 (
            .O(N__22187),
            .I(N__22141));
    InMux I__2515 (
            .O(N__22186),
            .I(N__22138));
    InMux I__2514 (
            .O(N__22183),
            .I(N__22135));
    InMux I__2513 (
            .O(N__22182),
            .I(N__22130));
    InMux I__2512 (
            .O(N__22181),
            .I(N__22130));
    InMux I__2511 (
            .O(N__22180),
            .I(N__22125));
    InMux I__2510 (
            .O(N__22179),
            .I(N__22125));
    InMux I__2509 (
            .O(N__22178),
            .I(N__22116));
    InMux I__2508 (
            .O(N__22177),
            .I(N__22116));
    InMux I__2507 (
            .O(N__22176),
            .I(N__22116));
    InMux I__2506 (
            .O(N__22175),
            .I(N__22116));
    CascadeMux I__2505 (
            .O(N__22174),
            .I(N__22112));
    CascadeMux I__2504 (
            .O(N__22173),
            .I(N__22108));
    Span4Mux_v I__2503 (
            .O(N__22170),
            .I(N__22105));
    InMux I__2502 (
            .O(N__22169),
            .I(N__22102));
    CascadeMux I__2501 (
            .O(N__22168),
            .I(N__22099));
    LocalMux I__2500 (
            .O(N__22157),
            .I(N__22091));
    InMux I__2499 (
            .O(N__22156),
            .I(N__22080));
    InMux I__2498 (
            .O(N__22155),
            .I(N__22080));
    InMux I__2497 (
            .O(N__22154),
            .I(N__22080));
    InMux I__2496 (
            .O(N__22153),
            .I(N__22080));
    InMux I__2495 (
            .O(N__22152),
            .I(N__22080));
    InMux I__2494 (
            .O(N__22149),
            .I(N__22077));
    Span4Mux_v I__2493 (
            .O(N__22146),
            .I(N__22074));
    LocalMux I__2492 (
            .O(N__22141),
            .I(N__22069));
    LocalMux I__2491 (
            .O(N__22138),
            .I(N__22069));
    LocalMux I__2490 (
            .O(N__22135),
            .I(N__22063));
    LocalMux I__2489 (
            .O(N__22130),
            .I(N__22058));
    LocalMux I__2488 (
            .O(N__22125),
            .I(N__22058));
    LocalMux I__2487 (
            .O(N__22116),
            .I(N__22055));
    InMux I__2486 (
            .O(N__22115),
            .I(N__22052));
    InMux I__2485 (
            .O(N__22112),
            .I(N__22047));
    InMux I__2484 (
            .O(N__22111),
            .I(N__22047));
    InMux I__2483 (
            .O(N__22108),
            .I(N__22044));
    Span4Mux_h I__2482 (
            .O(N__22105),
            .I(N__22039));
    LocalMux I__2481 (
            .O(N__22102),
            .I(N__22039));
    InMux I__2480 (
            .O(N__22099),
            .I(N__22034));
    InMux I__2479 (
            .O(N__22098),
            .I(N__22034));
    InMux I__2478 (
            .O(N__22097),
            .I(N__22025));
    InMux I__2477 (
            .O(N__22096),
            .I(N__22025));
    InMux I__2476 (
            .O(N__22095),
            .I(N__22025));
    InMux I__2475 (
            .O(N__22094),
            .I(N__22025));
    Span4Mux_v I__2474 (
            .O(N__22091),
            .I(N__22014));
    LocalMux I__2473 (
            .O(N__22080),
            .I(N__22014));
    LocalMux I__2472 (
            .O(N__22077),
            .I(N__22014));
    Span4Mux_h I__2471 (
            .O(N__22074),
            .I(N__22014));
    Span4Mux_v I__2470 (
            .O(N__22069),
            .I(N__22014));
    InMux I__2469 (
            .O(N__22068),
            .I(N__22007));
    InMux I__2468 (
            .O(N__22067),
            .I(N__22007));
    InMux I__2467 (
            .O(N__22066),
            .I(N__22007));
    Span4Mux_v I__2466 (
            .O(N__22063),
            .I(N__22000));
    Span4Mux_v I__2465 (
            .O(N__22058),
            .I(N__22000));
    Span4Mux_h I__2464 (
            .O(N__22055),
            .I(N__22000));
    LocalMux I__2463 (
            .O(N__22052),
            .I(adc_state_2));
    LocalMux I__2462 (
            .O(N__22047),
            .I(adc_state_2));
    LocalMux I__2461 (
            .O(N__22044),
            .I(adc_state_2));
    Odrv4 I__2460 (
            .O(N__22039),
            .I(adc_state_2));
    LocalMux I__2459 (
            .O(N__22034),
            .I(adc_state_2));
    LocalMux I__2458 (
            .O(N__22025),
            .I(adc_state_2));
    Odrv4 I__2457 (
            .O(N__22014),
            .I(adc_state_2));
    LocalMux I__2456 (
            .O(N__22007),
            .I(adc_state_2));
    Odrv4 I__2455 (
            .O(N__22000),
            .I(adc_state_2));
    InMux I__2454 (
            .O(N__21981),
            .I(N__21978));
    LocalMux I__2453 (
            .O(N__21978),
            .I(\RTD.cfg_tmp_0 ));
    CEMux I__2452 (
            .O(N__21975),
            .I(N__21972));
    LocalMux I__2451 (
            .O(N__21972),
            .I(\RTD.n13137 ));
    SRMux I__2450 (
            .O(N__21969),
            .I(N__21966));
    LocalMux I__2449 (
            .O(N__21966),
            .I(\RTD.n15115 ));
    CascadeMux I__2448 (
            .O(N__21963),
            .I(N__21959));
    InMux I__2447 (
            .O(N__21962),
            .I(N__21956));
    InMux I__2446 (
            .O(N__21959),
            .I(N__21953));
    LocalMux I__2445 (
            .O(N__21956),
            .I(\ADC_IAC.bit_cnt_6 ));
    LocalMux I__2444 (
            .O(N__21953),
            .I(\ADC_IAC.bit_cnt_6 ));
    InMux I__2443 (
            .O(N__21948),
            .I(\ADC_IAC.n19833 ));
    InMux I__2442 (
            .O(N__21945),
            .I(\ADC_IAC.n19834 ));
    InMux I__2441 (
            .O(N__21942),
            .I(N__21938));
    InMux I__2440 (
            .O(N__21941),
            .I(N__21935));
    LocalMux I__2439 (
            .O(N__21938),
            .I(\ADC_IAC.bit_cnt_7 ));
    LocalMux I__2438 (
            .O(N__21935),
            .I(\ADC_IAC.bit_cnt_7 ));
    CEMux I__2437 (
            .O(N__21930),
            .I(N__21927));
    LocalMux I__2436 (
            .O(N__21927),
            .I(N__21924));
    Span4Mux_v I__2435 (
            .O(N__21924),
            .I(N__21921));
    Odrv4 I__2434 (
            .O(N__21921),
            .I(\ADC_IAC.n12698 ));
    CascadeMux I__2433 (
            .O(N__21918),
            .I(\ADC_IAC.n12698_cascade_ ));
    SRMux I__2432 (
            .O(N__21915),
            .I(N__21912));
    LocalMux I__2431 (
            .O(N__21912),
            .I(N__21909));
    Span4Mux_h I__2430 (
            .O(N__21909),
            .I(N__21906));
    Odrv4 I__2429 (
            .O(N__21906),
            .I(\ADC_IAC.n15014 ));
    IoInMux I__2428 (
            .O(N__21903),
            .I(N__21900));
    LocalMux I__2427 (
            .O(N__21900),
            .I(N__21897));
    IoSpan4Mux I__2426 (
            .O(N__21897),
            .I(N__21894));
    IoSpan4Mux I__2425 (
            .O(N__21894),
            .I(N__21891));
    Span4Mux_s3_v I__2424 (
            .O(N__21891),
            .I(N__21888));
    Span4Mux_v I__2423 (
            .O(N__21888),
            .I(N__21885));
    Odrv4 I__2422 (
            .O(N__21885),
            .I(AC_ADC_SYNC));
    CascadeMux I__2421 (
            .O(N__21882),
            .I(n14_adj_1662_cascade_));
    IoInMux I__2420 (
            .O(N__21879),
            .I(N__21876));
    LocalMux I__2419 (
            .O(N__21876),
            .I(N__21873));
    Span4Mux_s3_v I__2418 (
            .O(N__21873),
            .I(N__21870));
    Span4Mux_v I__2417 (
            .O(N__21870),
            .I(N__21866));
    InMux I__2416 (
            .O(N__21869),
            .I(N__21863));
    Odrv4 I__2415 (
            .O(N__21866),
            .I(IAC_CS));
    LocalMux I__2414 (
            .O(N__21863),
            .I(IAC_CS));
    IoInMux I__2413 (
            .O(N__21858),
            .I(N__21855));
    LocalMux I__2412 (
            .O(N__21855),
            .I(N__21852));
    Span4Mux_s3_v I__2411 (
            .O(N__21852),
            .I(N__21849));
    Span4Mux_v I__2410 (
            .O(N__21849),
            .I(N__21846));
    Span4Mux_h I__2409 (
            .O(N__21846),
            .I(N__21843));
    Odrv4 I__2408 (
            .O(N__21843),
            .I(DDS_CS1));
    CascadeMux I__2407 (
            .O(N__21840),
            .I(\ADC_IAC.n21458_cascade_ ));
    InMux I__2406 (
            .O(N__21837),
            .I(N__21834));
    LocalMux I__2405 (
            .O(N__21834),
            .I(\ADC_IAC.n16 ));
    InMux I__2404 (
            .O(N__21831),
            .I(N__21827));
    InMux I__2403 (
            .O(N__21830),
            .I(N__21824));
    LocalMux I__2402 (
            .O(N__21827),
            .I(\ADC_IAC.bit_cnt_0 ));
    LocalMux I__2401 (
            .O(N__21824),
            .I(\ADC_IAC.bit_cnt_0 ));
    InMux I__2400 (
            .O(N__21819),
            .I(bfn_6_18_0_));
    InMux I__2399 (
            .O(N__21816),
            .I(N__21812));
    InMux I__2398 (
            .O(N__21815),
            .I(N__21809));
    LocalMux I__2397 (
            .O(N__21812),
            .I(\ADC_IAC.bit_cnt_1 ));
    LocalMux I__2396 (
            .O(N__21809),
            .I(\ADC_IAC.bit_cnt_1 ));
    InMux I__2395 (
            .O(N__21804),
            .I(\ADC_IAC.n19828 ));
    InMux I__2394 (
            .O(N__21801),
            .I(N__21797));
    InMux I__2393 (
            .O(N__21800),
            .I(N__21794));
    LocalMux I__2392 (
            .O(N__21797),
            .I(\ADC_IAC.bit_cnt_2 ));
    LocalMux I__2391 (
            .O(N__21794),
            .I(\ADC_IAC.bit_cnt_2 ));
    InMux I__2390 (
            .O(N__21789),
            .I(\ADC_IAC.n19829 ));
    InMux I__2389 (
            .O(N__21786),
            .I(N__21782));
    InMux I__2388 (
            .O(N__21785),
            .I(N__21779));
    LocalMux I__2387 (
            .O(N__21782),
            .I(\ADC_IAC.bit_cnt_3 ));
    LocalMux I__2386 (
            .O(N__21779),
            .I(\ADC_IAC.bit_cnt_3 ));
    InMux I__2385 (
            .O(N__21774),
            .I(\ADC_IAC.n19830 ));
    InMux I__2384 (
            .O(N__21771),
            .I(N__21767));
    InMux I__2383 (
            .O(N__21770),
            .I(N__21764));
    LocalMux I__2382 (
            .O(N__21767),
            .I(\ADC_IAC.bit_cnt_4 ));
    LocalMux I__2381 (
            .O(N__21764),
            .I(\ADC_IAC.bit_cnt_4 ));
    InMux I__2380 (
            .O(N__21759),
            .I(\ADC_IAC.n19831 ));
    CascadeMux I__2379 (
            .O(N__21756),
            .I(N__21752));
    InMux I__2378 (
            .O(N__21755),
            .I(N__21749));
    InMux I__2377 (
            .O(N__21752),
            .I(N__21746));
    LocalMux I__2376 (
            .O(N__21749),
            .I(\ADC_IAC.bit_cnt_5 ));
    LocalMux I__2375 (
            .O(N__21746),
            .I(\ADC_IAC.bit_cnt_5 ));
    InMux I__2374 (
            .O(N__21741),
            .I(\ADC_IAC.n19832 ));
    CEMux I__2373 (
            .O(N__21738),
            .I(N__21735));
    LocalMux I__2372 (
            .O(N__21735),
            .I(N__21732));
    Odrv4 I__2371 (
            .O(N__21732),
            .I(\ADC_VAC.n12 ));
    InMux I__2370 (
            .O(N__21729),
            .I(N__21726));
    LocalMux I__2369 (
            .O(N__21726),
            .I(n21050));
    CascadeMux I__2368 (
            .O(N__21723),
            .I(N__21719));
    CascadeMux I__2367 (
            .O(N__21722),
            .I(N__21716));
    InMux I__2366 (
            .O(N__21719),
            .I(N__21710));
    InMux I__2365 (
            .O(N__21716),
            .I(N__21707));
    InMux I__2364 (
            .O(N__21715),
            .I(N__21704));
    InMux I__2363 (
            .O(N__21714),
            .I(N__21701));
    CascadeMux I__2362 (
            .O(N__21713),
            .I(N__21698));
    LocalMux I__2361 (
            .O(N__21710),
            .I(N__21695));
    LocalMux I__2360 (
            .O(N__21707),
            .I(N__21692));
    LocalMux I__2359 (
            .O(N__21704),
            .I(N__21689));
    LocalMux I__2358 (
            .O(N__21701),
            .I(N__21686));
    InMux I__2357 (
            .O(N__21698),
            .I(N__21683));
    Span4Mux_v I__2356 (
            .O(N__21695),
            .I(N__21678));
    Span4Mux_v I__2355 (
            .O(N__21692),
            .I(N__21678));
    Span4Mux_v I__2354 (
            .O(N__21689),
            .I(N__21671));
    Span4Mux_v I__2353 (
            .O(N__21686),
            .I(N__21671));
    LocalMux I__2352 (
            .O(N__21683),
            .I(N__21671));
    Sp12to4 I__2351 (
            .O(N__21678),
            .I(N__21666));
    Sp12to4 I__2350 (
            .O(N__21671),
            .I(N__21666));
    Odrv12 I__2349 (
            .O(N__21666),
            .I(VAC_DRDY));
    CascadeMux I__2348 (
            .O(N__21663),
            .I(n21050_cascade_));
    IoInMux I__2347 (
            .O(N__21660),
            .I(N__21657));
    LocalMux I__2346 (
            .O(N__21657),
            .I(N__21654));
    Span4Mux_s3_h I__2345 (
            .O(N__21654),
            .I(N__21651));
    Span4Mux_h I__2344 (
            .O(N__21651),
            .I(N__21647));
    InMux I__2343 (
            .O(N__21650),
            .I(N__21644));
    Span4Mux_v I__2342 (
            .O(N__21647),
            .I(N__21641));
    LocalMux I__2341 (
            .O(N__21644),
            .I(N__21638));
    Odrv4 I__2340 (
            .O(N__21641),
            .I(VAC_CS));
    Odrv4 I__2339 (
            .O(N__21638),
            .I(VAC_CS));
    InMux I__2338 (
            .O(N__21633),
            .I(N__21630));
    LocalMux I__2337 (
            .O(N__21630),
            .I(n14_adj_1657));
    CascadeMux I__2336 (
            .O(N__21627),
            .I(N__21622));
    CascadeMux I__2335 (
            .O(N__21626),
            .I(N__21613));
    CascadeMux I__2334 (
            .O(N__21625),
            .I(N__21609));
    InMux I__2333 (
            .O(N__21622),
            .I(N__21604));
    InMux I__2332 (
            .O(N__21621),
            .I(N__21601));
    InMux I__2331 (
            .O(N__21620),
            .I(N__21598));
    InMux I__2330 (
            .O(N__21619),
            .I(N__21595));
    InMux I__2329 (
            .O(N__21618),
            .I(N__21592));
    InMux I__2328 (
            .O(N__21617),
            .I(N__21587));
    InMux I__2327 (
            .O(N__21616),
            .I(N__21587));
    InMux I__2326 (
            .O(N__21613),
            .I(N__21576));
    InMux I__2325 (
            .O(N__21612),
            .I(N__21576));
    InMux I__2324 (
            .O(N__21609),
            .I(N__21576));
    InMux I__2323 (
            .O(N__21608),
            .I(N__21576));
    InMux I__2322 (
            .O(N__21607),
            .I(N__21576));
    LocalMux I__2321 (
            .O(N__21604),
            .I(N__21569));
    LocalMux I__2320 (
            .O(N__21601),
            .I(N__21569));
    LocalMux I__2319 (
            .O(N__21598),
            .I(N__21569));
    LocalMux I__2318 (
            .O(N__21595),
            .I(DTRIG_N_958_adj_1493));
    LocalMux I__2317 (
            .O(N__21592),
            .I(DTRIG_N_958_adj_1493));
    LocalMux I__2316 (
            .O(N__21587),
            .I(DTRIG_N_958_adj_1493));
    LocalMux I__2315 (
            .O(N__21576),
            .I(DTRIG_N_958_adj_1493));
    Odrv4 I__2314 (
            .O(N__21569),
            .I(DTRIG_N_958_adj_1493));
    InMux I__2313 (
            .O(N__21558),
            .I(N__21547));
    InMux I__2312 (
            .O(N__21557),
            .I(N__21547));
    InMux I__2311 (
            .O(N__21556),
            .I(N__21544));
    InMux I__2310 (
            .O(N__21555),
            .I(N__21536));
    InMux I__2309 (
            .O(N__21554),
            .I(N__21533));
    InMux I__2308 (
            .O(N__21553),
            .I(N__21528));
    InMux I__2307 (
            .O(N__21552),
            .I(N__21528));
    LocalMux I__2306 (
            .O(N__21547),
            .I(N__21523));
    LocalMux I__2305 (
            .O(N__21544),
            .I(N__21523));
    InMux I__2304 (
            .O(N__21543),
            .I(N__21512));
    InMux I__2303 (
            .O(N__21542),
            .I(N__21512));
    InMux I__2302 (
            .O(N__21541),
            .I(N__21512));
    InMux I__2301 (
            .O(N__21540),
            .I(N__21512));
    InMux I__2300 (
            .O(N__21539),
            .I(N__21512));
    LocalMux I__2299 (
            .O(N__21536),
            .I(adc_state_1_adj_1459));
    LocalMux I__2298 (
            .O(N__21533),
            .I(adc_state_1_adj_1459));
    LocalMux I__2297 (
            .O(N__21528),
            .I(adc_state_1_adj_1459));
    Odrv4 I__2296 (
            .O(N__21523),
            .I(adc_state_1_adj_1459));
    LocalMux I__2295 (
            .O(N__21512),
            .I(adc_state_1_adj_1459));
    CascadeMux I__2294 (
            .O(N__21501),
            .I(N__21498));
    InMux I__2293 (
            .O(N__21498),
            .I(N__21493));
    CascadeMux I__2292 (
            .O(N__21497),
            .I(N__21490));
    CascadeMux I__2291 (
            .O(N__21496),
            .I(N__21487));
    LocalMux I__2290 (
            .O(N__21493),
            .I(N__21484));
    InMux I__2289 (
            .O(N__21490),
            .I(N__21479));
    InMux I__2288 (
            .O(N__21487),
            .I(N__21479));
    Odrv12 I__2287 (
            .O(N__21484),
            .I(cmd_rdadctmp_14));
    LocalMux I__2286 (
            .O(N__21479),
            .I(cmd_rdadctmp_14));
    InMux I__2285 (
            .O(N__21474),
            .I(N__21471));
    LocalMux I__2284 (
            .O(N__21471),
            .I(\ADC_VAC.n17 ));
    IoInMux I__2283 (
            .O(N__21468),
            .I(N__21465));
    LocalMux I__2282 (
            .O(N__21465),
            .I(N__21462));
    IoSpan4Mux I__2281 (
            .O(N__21462),
            .I(N__21459));
    Span4Mux_s2_h I__2280 (
            .O(N__21459),
            .I(N__21455));
    CascadeMux I__2279 (
            .O(N__21458),
            .I(N__21452));
    Span4Mux_h I__2278 (
            .O(N__21455),
            .I(N__21449));
    InMux I__2277 (
            .O(N__21452),
            .I(N__21446));
    Odrv4 I__2276 (
            .O(N__21449),
            .I(VAC_SCLK));
    LocalMux I__2275 (
            .O(N__21446),
            .I(VAC_SCLK));
    CascadeMux I__2274 (
            .O(N__21441),
            .I(N__21437));
    InMux I__2273 (
            .O(N__21440),
            .I(N__21429));
    InMux I__2272 (
            .O(N__21437),
            .I(N__21429));
    InMux I__2271 (
            .O(N__21436),
            .I(N__21429));
    LocalMux I__2270 (
            .O(N__21429),
            .I(cmd_rdadctmp_26_adj_1466));
    CascadeMux I__2269 (
            .O(N__21426),
            .I(N__21423));
    InMux I__2268 (
            .O(N__21423),
            .I(N__21420));
    LocalMux I__2267 (
            .O(N__21420),
            .I(N__21417));
    Span4Mux_v I__2266 (
            .O(N__21417),
            .I(N__21413));
    InMux I__2265 (
            .O(N__21416),
            .I(N__21410));
    Odrv4 I__2264 (
            .O(N__21413),
            .I(cmd_rdadctmp_3_adj_1489));
    LocalMux I__2263 (
            .O(N__21410),
            .I(cmd_rdadctmp_3_adj_1489));
    InMux I__2262 (
            .O(N__21405),
            .I(N__21402));
    LocalMux I__2261 (
            .O(N__21402),
            .I(N__21399));
    Span4Mux_h I__2260 (
            .O(N__21399),
            .I(N__21395));
    InMux I__2259 (
            .O(N__21398),
            .I(N__21391));
    Span4Mux_v I__2258 (
            .O(N__21395),
            .I(N__21388));
    InMux I__2257 (
            .O(N__21394),
            .I(N__21385));
    LocalMux I__2256 (
            .O(N__21391),
            .I(buf_adcdata_iac_7));
    Odrv4 I__2255 (
            .O(N__21388),
            .I(buf_adcdata_iac_7));
    LocalMux I__2254 (
            .O(N__21385),
            .I(buf_adcdata_iac_7));
    CascadeMux I__2253 (
            .O(N__21378),
            .I(N__21374));
    CascadeMux I__2252 (
            .O(N__21377),
            .I(N__21371));
    InMux I__2251 (
            .O(N__21374),
            .I(N__21368));
    InMux I__2250 (
            .O(N__21371),
            .I(N__21364));
    LocalMux I__2249 (
            .O(N__21368),
            .I(N__21361));
    InMux I__2248 (
            .O(N__21367),
            .I(N__21358));
    LocalMux I__2247 (
            .O(N__21364),
            .I(cmd_rdadctmp_8_adj_1484));
    Odrv4 I__2246 (
            .O(N__21361),
            .I(cmd_rdadctmp_8_adj_1484));
    LocalMux I__2245 (
            .O(N__21358),
            .I(cmd_rdadctmp_8_adj_1484));
    InMux I__2244 (
            .O(N__21351),
            .I(N__21348));
    LocalMux I__2243 (
            .O(N__21348),
            .I(N__21345));
    Span4Mux_h I__2242 (
            .O(N__21345),
            .I(N__21342));
    Sp12to4 I__2241 (
            .O(N__21342),
            .I(N__21339));
    Odrv12 I__2240 (
            .O(N__21339),
            .I(buf_data_iac_7));
    InMux I__2239 (
            .O(N__21336),
            .I(N__21333));
    LocalMux I__2238 (
            .O(N__21333),
            .I(n22_adj_1598));
    InMux I__2237 (
            .O(N__21330),
            .I(N__21323));
    InMux I__2236 (
            .O(N__21329),
            .I(N__21323));
    InMux I__2235 (
            .O(N__21328),
            .I(N__21320));
    LocalMux I__2234 (
            .O(N__21323),
            .I(cmd_rdadctmp_12_adj_1480));
    LocalMux I__2233 (
            .O(N__21320),
            .I(cmd_rdadctmp_12_adj_1480));
    InMux I__2232 (
            .O(N__21315),
            .I(N__21311));
    CascadeMux I__2231 (
            .O(N__21314),
            .I(N__21308));
    LocalMux I__2230 (
            .O(N__21311),
            .I(N__21304));
    InMux I__2229 (
            .O(N__21308),
            .I(N__21301));
    InMux I__2228 (
            .O(N__21307),
            .I(N__21298));
    Span12Mux_s9_h I__2227 (
            .O(N__21304),
            .I(N__21295));
    LocalMux I__2226 (
            .O(N__21301),
            .I(buf_adcdata_iac_4));
    LocalMux I__2225 (
            .O(N__21298),
            .I(buf_adcdata_iac_4));
    Odrv12 I__2224 (
            .O(N__21295),
            .I(buf_adcdata_iac_4));
    InMux I__2223 (
            .O(N__21288),
            .I(N__21284));
    CascadeMux I__2222 (
            .O(N__21287),
            .I(N__21281));
    LocalMux I__2221 (
            .O(N__21284),
            .I(N__21278));
    InMux I__2220 (
            .O(N__21281),
            .I(N__21274));
    Span4Mux_h I__2219 (
            .O(N__21278),
            .I(N__21271));
    InMux I__2218 (
            .O(N__21277),
            .I(N__21268));
    LocalMux I__2217 (
            .O(N__21274),
            .I(buf_adcdata_vac_4));
    Odrv4 I__2216 (
            .O(N__21271),
            .I(buf_adcdata_vac_4));
    LocalMux I__2215 (
            .O(N__21268),
            .I(buf_adcdata_vac_4));
    CascadeMux I__2214 (
            .O(N__21261),
            .I(n19_adj_1606_cascade_));
    InMux I__2213 (
            .O(N__21258),
            .I(N__21255));
    LocalMux I__2212 (
            .O(N__21255),
            .I(N__21252));
    Span4Mux_h I__2211 (
            .O(N__21252),
            .I(N__21249));
    Span4Mux_v I__2210 (
            .O(N__21249),
            .I(N__21246));
    Odrv4 I__2209 (
            .O(N__21246),
            .I(buf_data_iac_4));
    CascadeMux I__2208 (
            .O(N__21243),
            .I(n22_adj_1607_cascade_));
    CascadeMux I__2207 (
            .O(N__21240),
            .I(N__21237));
    InMux I__2206 (
            .O(N__21237),
            .I(N__21233));
    InMux I__2205 (
            .O(N__21236),
            .I(N__21230));
    LocalMux I__2204 (
            .O(N__21233),
            .I(cmd_rdadctmp_31_adj_1461));
    LocalMux I__2203 (
            .O(N__21230),
            .I(cmd_rdadctmp_31_adj_1461));
    CascadeMux I__2202 (
            .O(N__21225),
            .I(N__21222));
    InMux I__2201 (
            .O(N__21222),
            .I(N__21219));
    LocalMux I__2200 (
            .O(N__21219),
            .I(N__21215));
    InMux I__2199 (
            .O(N__21218),
            .I(N__21212));
    Span4Mux_v I__2198 (
            .O(N__21215),
            .I(N__21206));
    LocalMux I__2197 (
            .O(N__21212),
            .I(N__21206));
    InMux I__2196 (
            .O(N__21211),
            .I(N__21203));
    Odrv4 I__2195 (
            .O(N__21206),
            .I(read_buf_0));
    LocalMux I__2194 (
            .O(N__21203),
            .I(read_buf_0));
    InMux I__2193 (
            .O(N__21198),
            .I(N__21193));
    CascadeMux I__2192 (
            .O(N__21197),
            .I(N__21190));
    CascadeMux I__2191 (
            .O(N__21196),
            .I(N__21187));
    LocalMux I__2190 (
            .O(N__21193),
            .I(N__21184));
    InMux I__2189 (
            .O(N__21190),
            .I(N__21179));
    InMux I__2188 (
            .O(N__21187),
            .I(N__21179));
    Odrv12 I__2187 (
            .O(N__21184),
            .I(read_buf_2));
    LocalMux I__2186 (
            .O(N__21179),
            .I(read_buf_2));
    CascadeMux I__2185 (
            .O(N__21174),
            .I(N__21170));
    CascadeMux I__2184 (
            .O(N__21173),
            .I(N__21166));
    InMux I__2183 (
            .O(N__21170),
            .I(N__21156));
    InMux I__2182 (
            .O(N__21169),
            .I(N__21156));
    InMux I__2181 (
            .O(N__21166),
            .I(N__21142));
    InMux I__2180 (
            .O(N__21165),
            .I(N__21142));
    InMux I__2179 (
            .O(N__21164),
            .I(N__21142));
    InMux I__2178 (
            .O(N__21163),
            .I(N__21137));
    InMux I__2177 (
            .O(N__21162),
            .I(N__21137));
    InMux I__2176 (
            .O(N__21161),
            .I(N__21134));
    LocalMux I__2175 (
            .O(N__21156),
            .I(N__21131));
    InMux I__2174 (
            .O(N__21155),
            .I(N__21126));
    InMux I__2173 (
            .O(N__21154),
            .I(N__21126));
    InMux I__2172 (
            .O(N__21153),
            .I(N__21115));
    InMux I__2171 (
            .O(N__21152),
            .I(N__21115));
    InMux I__2170 (
            .O(N__21151),
            .I(N__21115));
    InMux I__2169 (
            .O(N__21150),
            .I(N__21115));
    InMux I__2168 (
            .O(N__21149),
            .I(N__21115));
    LocalMux I__2167 (
            .O(N__21142),
            .I(n11856));
    LocalMux I__2166 (
            .O(N__21137),
            .I(n11856));
    LocalMux I__2165 (
            .O(N__21134),
            .I(n11856));
    Odrv4 I__2164 (
            .O(N__21131),
            .I(n11856));
    LocalMux I__2163 (
            .O(N__21126),
            .I(n11856));
    LocalMux I__2162 (
            .O(N__21115),
            .I(n11856));
    CascadeMux I__2161 (
            .O(N__21102),
            .I(N__21097));
    InMux I__2160 (
            .O(N__21101),
            .I(N__21092));
    InMux I__2159 (
            .O(N__21100),
            .I(N__21092));
    InMux I__2158 (
            .O(N__21097),
            .I(N__21089));
    LocalMux I__2157 (
            .O(N__21092),
            .I(read_buf_1));
    LocalMux I__2156 (
            .O(N__21089),
            .I(read_buf_1));
    InMux I__2155 (
            .O(N__21084),
            .I(N__21079));
    InMux I__2154 (
            .O(N__21083),
            .I(N__21074));
    InMux I__2153 (
            .O(N__21082),
            .I(N__21074));
    LocalMux I__2152 (
            .O(N__21079),
            .I(read_buf_12));
    LocalMux I__2151 (
            .O(N__21074),
            .I(read_buf_12));
    InMux I__2150 (
            .O(N__21069),
            .I(N__21064));
    CascadeMux I__2149 (
            .O(N__21068),
            .I(N__21061));
    CascadeMux I__2148 (
            .O(N__21067),
            .I(N__21058));
    LocalMux I__2147 (
            .O(N__21064),
            .I(N__21055));
    InMux I__2146 (
            .O(N__21061),
            .I(N__21050));
    InMux I__2145 (
            .O(N__21058),
            .I(N__21050));
    Odrv4 I__2144 (
            .O(N__21055),
            .I(read_buf_13));
    LocalMux I__2143 (
            .O(N__21050),
            .I(read_buf_13));
    InMux I__2142 (
            .O(N__21045),
            .I(N__21035));
    CascadeMux I__2141 (
            .O(N__21044),
            .I(N__21032));
    InMux I__2140 (
            .O(N__21043),
            .I(N__21018));
    InMux I__2139 (
            .O(N__21042),
            .I(N__21018));
    InMux I__2138 (
            .O(N__21041),
            .I(N__21018));
    InMux I__2137 (
            .O(N__21040),
            .I(N__21011));
    InMux I__2136 (
            .O(N__21039),
            .I(N__21011));
    InMux I__2135 (
            .O(N__21038),
            .I(N__21011));
    LocalMux I__2134 (
            .O(N__21035),
            .I(N__21008));
    InMux I__2133 (
            .O(N__21032),
            .I(N__21005));
    InMux I__2132 (
            .O(N__21031),
            .I(N__20996));
    InMux I__2131 (
            .O(N__21030),
            .I(N__20996));
    InMux I__2130 (
            .O(N__21029),
            .I(N__20996));
    InMux I__2129 (
            .O(N__21028),
            .I(N__20996));
    InMux I__2128 (
            .O(N__21027),
            .I(N__20989));
    InMux I__2127 (
            .O(N__21026),
            .I(N__20989));
    InMux I__2126 (
            .O(N__21025),
            .I(N__20989));
    LocalMux I__2125 (
            .O(N__21018),
            .I(n13212));
    LocalMux I__2124 (
            .O(N__21011),
            .I(n13212));
    Odrv4 I__2123 (
            .O(N__21008),
            .I(n13212));
    LocalMux I__2122 (
            .O(N__21005),
            .I(n13212));
    LocalMux I__2121 (
            .O(N__20996),
            .I(n13212));
    LocalMux I__2120 (
            .O(N__20989),
            .I(n13212));
    CascadeMux I__2119 (
            .O(N__20976),
            .I(N__20971));
    CascadeMux I__2118 (
            .O(N__20975),
            .I(N__20965));
    CascadeMux I__2117 (
            .O(N__20974),
            .I(N__20962));
    InMux I__2116 (
            .O(N__20971),
            .I(N__20952));
    InMux I__2115 (
            .O(N__20970),
            .I(N__20952));
    InMux I__2114 (
            .O(N__20969),
            .I(N__20952));
    InMux I__2113 (
            .O(N__20968),
            .I(N__20946));
    InMux I__2112 (
            .O(N__20965),
            .I(N__20935));
    InMux I__2111 (
            .O(N__20962),
            .I(N__20935));
    InMux I__2110 (
            .O(N__20961),
            .I(N__20935));
    InMux I__2109 (
            .O(N__20960),
            .I(N__20935));
    InMux I__2108 (
            .O(N__20959),
            .I(N__20935));
    LocalMux I__2107 (
            .O(N__20952),
            .I(N__20932));
    InMux I__2106 (
            .O(N__20951),
            .I(N__20925));
    InMux I__2105 (
            .O(N__20950),
            .I(N__20925));
    InMux I__2104 (
            .O(N__20949),
            .I(N__20925));
    LocalMux I__2103 (
            .O(N__20946),
            .I(N__20918));
    LocalMux I__2102 (
            .O(N__20935),
            .I(N__20915));
    Span4Mux_v I__2101 (
            .O(N__20932),
            .I(N__20910));
    LocalMux I__2100 (
            .O(N__20925),
            .I(N__20910));
    InMux I__2099 (
            .O(N__20924),
            .I(N__20903));
    InMux I__2098 (
            .O(N__20923),
            .I(N__20903));
    InMux I__2097 (
            .O(N__20922),
            .I(N__20903));
    InMux I__2096 (
            .O(N__20921),
            .I(N__20900));
    Span4Mux_v I__2095 (
            .O(N__20918),
            .I(N__20895));
    Span4Mux_v I__2094 (
            .O(N__20915),
            .I(N__20895));
    Span4Mux_h I__2093 (
            .O(N__20910),
            .I(N__20892));
    LocalMux I__2092 (
            .O(N__20903),
            .I(N__20887));
    LocalMux I__2091 (
            .O(N__20900),
            .I(N__20887));
    Odrv4 I__2090 (
            .O(N__20895),
            .I(n1_adj_1592));
    Odrv4 I__2089 (
            .O(N__20892),
            .I(n1_adj_1592));
    Odrv4 I__2088 (
            .O(N__20887),
            .I(n1_adj_1592));
    CascadeMux I__2087 (
            .O(N__20880),
            .I(N__20877));
    InMux I__2086 (
            .O(N__20877),
            .I(N__20873));
    InMux I__2085 (
            .O(N__20876),
            .I(N__20869));
    LocalMux I__2084 (
            .O(N__20873),
            .I(N__20866));
    InMux I__2083 (
            .O(N__20872),
            .I(N__20863));
    LocalMux I__2082 (
            .O(N__20869),
            .I(read_buf_6));
    Odrv4 I__2081 (
            .O(N__20866),
            .I(read_buf_6));
    LocalMux I__2080 (
            .O(N__20863),
            .I(read_buf_6));
    InMux I__2079 (
            .O(N__20856),
            .I(N__20851));
    InMux I__2078 (
            .O(N__20855),
            .I(N__20846));
    InMux I__2077 (
            .O(N__20854),
            .I(N__20846));
    LocalMux I__2076 (
            .O(N__20851),
            .I(read_buf_7));
    LocalMux I__2075 (
            .O(N__20846),
            .I(read_buf_7));
    InMux I__2074 (
            .O(N__20841),
            .I(N__20838));
    LocalMux I__2073 (
            .O(N__20838),
            .I(N__20835));
    Span4Mux_h I__2072 (
            .O(N__20835),
            .I(N__20831));
    InMux I__2071 (
            .O(N__20834),
            .I(N__20827));
    Span4Mux_v I__2070 (
            .O(N__20831),
            .I(N__20824));
    InMux I__2069 (
            .O(N__20830),
            .I(N__20821));
    LocalMux I__2068 (
            .O(N__20827),
            .I(buf_adcdata_iac_6));
    Odrv4 I__2067 (
            .O(N__20824),
            .I(buf_adcdata_iac_6));
    LocalMux I__2066 (
            .O(N__20821),
            .I(buf_adcdata_iac_6));
    SRMux I__2065 (
            .O(N__20814),
            .I(N__20811));
    LocalMux I__2064 (
            .O(N__20811),
            .I(N__20807));
    SRMux I__2063 (
            .O(N__20810),
            .I(N__20804));
    Span4Mux_v I__2062 (
            .O(N__20807),
            .I(N__20801));
    LocalMux I__2061 (
            .O(N__20804),
            .I(N__20798));
    Span4Mux_h I__2060 (
            .O(N__20801),
            .I(N__20795));
    Span4Mux_h I__2059 (
            .O(N__20798),
            .I(N__20790));
    Span4Mux_h I__2058 (
            .O(N__20795),
            .I(N__20790));
    Odrv4 I__2057 (
            .O(N__20790),
            .I(\RTD.n20370 ));
    InMux I__2056 (
            .O(N__20787),
            .I(N__20783));
    InMux I__2055 (
            .O(N__20786),
            .I(N__20780));
    LocalMux I__2054 (
            .O(N__20783),
            .I(\RTD.cfg_buf_6 ));
    LocalMux I__2053 (
            .O(N__20780),
            .I(\RTD.cfg_buf_6 ));
    CascadeMux I__2052 (
            .O(N__20775),
            .I(N__20771));
    CascadeMux I__2051 (
            .O(N__20774),
            .I(N__20768));
    InMux I__2050 (
            .O(N__20771),
            .I(N__20764));
    InMux I__2049 (
            .O(N__20768),
            .I(N__20759));
    InMux I__2048 (
            .O(N__20767),
            .I(N__20759));
    LocalMux I__2047 (
            .O(N__20764),
            .I(read_buf_9));
    LocalMux I__2046 (
            .O(N__20759),
            .I(read_buf_9));
    CascadeMux I__2045 (
            .O(N__20754),
            .I(N__20745));
    InMux I__2044 (
            .O(N__20753),
            .I(N__20735));
    InMux I__2043 (
            .O(N__20752),
            .I(N__20735));
    InMux I__2042 (
            .O(N__20751),
            .I(N__20735));
    InMux I__2041 (
            .O(N__20750),
            .I(N__20730));
    InMux I__2040 (
            .O(N__20749),
            .I(N__20730));
    InMux I__2039 (
            .O(N__20748),
            .I(N__20718));
    InMux I__2038 (
            .O(N__20745),
            .I(N__20718));
    InMux I__2037 (
            .O(N__20744),
            .I(N__20718));
    InMux I__2036 (
            .O(N__20743),
            .I(N__20713));
    InMux I__2035 (
            .O(N__20742),
            .I(N__20713));
    LocalMux I__2034 (
            .O(N__20735),
            .I(N__20706));
    LocalMux I__2033 (
            .O(N__20730),
            .I(N__20706));
    InMux I__2032 (
            .O(N__20729),
            .I(N__20697));
    InMux I__2031 (
            .O(N__20728),
            .I(N__20697));
    InMux I__2030 (
            .O(N__20727),
            .I(N__20697));
    InMux I__2029 (
            .O(N__20726),
            .I(N__20697));
    InMux I__2028 (
            .O(N__20725),
            .I(N__20694));
    LocalMux I__2027 (
            .O(N__20718),
            .I(N__20691));
    LocalMux I__2026 (
            .O(N__20713),
            .I(N__20688));
    InMux I__2025 (
            .O(N__20712),
            .I(N__20680));
    InMux I__2024 (
            .O(N__20711),
            .I(N__20680));
    Span4Mux_v I__2023 (
            .O(N__20706),
            .I(N__20674));
    LocalMux I__2022 (
            .O(N__20697),
            .I(N__20674));
    LocalMux I__2021 (
            .O(N__20694),
            .I(N__20666));
    Span4Mux_v I__2020 (
            .O(N__20691),
            .I(N__20666));
    Span4Mux_h I__2019 (
            .O(N__20688),
            .I(N__20663));
    InMux I__2018 (
            .O(N__20687),
            .I(N__20656));
    InMux I__2017 (
            .O(N__20686),
            .I(N__20656));
    InMux I__2016 (
            .O(N__20685),
            .I(N__20656));
    LocalMux I__2015 (
            .O(N__20680),
            .I(N__20653));
    InMux I__2014 (
            .O(N__20679),
            .I(N__20650));
    Span4Mux_h I__2013 (
            .O(N__20674),
            .I(N__20647));
    InMux I__2012 (
            .O(N__20673),
            .I(N__20640));
    InMux I__2011 (
            .O(N__20672),
            .I(N__20640));
    InMux I__2010 (
            .O(N__20671),
            .I(N__20640));
    Odrv4 I__2009 (
            .O(N__20666),
            .I(\RTD.adc_state_1 ));
    Odrv4 I__2008 (
            .O(N__20663),
            .I(\RTD.adc_state_1 ));
    LocalMux I__2007 (
            .O(N__20656),
            .I(\RTD.adc_state_1 ));
    Odrv4 I__2006 (
            .O(N__20653),
            .I(\RTD.adc_state_1 ));
    LocalMux I__2005 (
            .O(N__20650),
            .I(\RTD.adc_state_1 ));
    Odrv4 I__2004 (
            .O(N__20647),
            .I(\RTD.adc_state_1 ));
    LocalMux I__2003 (
            .O(N__20640),
            .I(\RTD.adc_state_1 ));
    CEMux I__2002 (
            .O(N__20625),
            .I(N__20622));
    LocalMux I__2001 (
            .O(N__20622),
            .I(N__20619));
    Span4Mux_v I__2000 (
            .O(N__20619),
            .I(N__20616));
    Span4Mux_h I__1999 (
            .O(N__20616),
            .I(N__20613));
    Odrv4 I__1998 (
            .O(N__20613),
            .I(\RTD.n11829 ));
    CascadeMux I__1997 (
            .O(N__20610),
            .I(N__20605));
    CascadeMux I__1996 (
            .O(N__20609),
            .I(N__20602));
    CascadeMux I__1995 (
            .O(N__20608),
            .I(N__20599));
    InMux I__1994 (
            .O(N__20605),
            .I(N__20592));
    InMux I__1993 (
            .O(N__20602),
            .I(N__20592));
    InMux I__1992 (
            .O(N__20599),
            .I(N__20592));
    LocalMux I__1991 (
            .O(N__20592),
            .I(read_buf_8));
    InMux I__1990 (
            .O(N__20589),
            .I(N__20586));
    LocalMux I__1989 (
            .O(N__20586),
            .I(N__20583));
    Span4Mux_v I__1988 (
            .O(N__20583),
            .I(N__20576));
    InMux I__1987 (
            .O(N__20582),
            .I(N__20571));
    InMux I__1986 (
            .O(N__20581),
            .I(N__20571));
    InMux I__1985 (
            .O(N__20580),
            .I(N__20566));
    InMux I__1984 (
            .O(N__20579),
            .I(N__20566));
    Odrv4 I__1983 (
            .O(N__20576),
            .I(\RTD.bit_cnt_3 ));
    LocalMux I__1982 (
            .O(N__20571),
            .I(\RTD.bit_cnt_3 ));
    LocalMux I__1981 (
            .O(N__20566),
            .I(\RTD.bit_cnt_3 ));
    InMux I__1980 (
            .O(N__20559),
            .I(N__20556));
    LocalMux I__1979 (
            .O(N__20556),
            .I(N__20551));
    InMux I__1978 (
            .O(N__20555),
            .I(N__20548));
    InMux I__1977 (
            .O(N__20554),
            .I(N__20545));
    Odrv4 I__1976 (
            .O(N__20551),
            .I(\RTD.n18043 ));
    LocalMux I__1975 (
            .O(N__20548),
            .I(\RTD.n18043 ));
    LocalMux I__1974 (
            .O(N__20545),
            .I(\RTD.n18043 ));
    InMux I__1973 (
            .O(N__20538),
            .I(N__20535));
    LocalMux I__1972 (
            .O(N__20535),
            .I(N__20531));
    InMux I__1971 (
            .O(N__20534),
            .I(N__20528));
    Span4Mux_h I__1970 (
            .O(N__20531),
            .I(N__20525));
    LocalMux I__1969 (
            .O(N__20528),
            .I(N__20522));
    Odrv4 I__1968 (
            .O(N__20525),
            .I(\RTD.n19026 ));
    Odrv12 I__1967 (
            .O(N__20522),
            .I(\RTD.n19026 ));
    CascadeMux I__1966 (
            .O(N__20517),
            .I(N__20513));
    InMux I__1965 (
            .O(N__20516),
            .I(N__20510));
    InMux I__1964 (
            .O(N__20513),
            .I(N__20507));
    LocalMux I__1963 (
            .O(N__20510),
            .I(adress_6));
    LocalMux I__1962 (
            .O(N__20507),
            .I(adress_6));
    CascadeMux I__1961 (
            .O(N__20502),
            .I(\RTD.n9_cascade_ ));
    CascadeMux I__1960 (
            .O(N__20499),
            .I(\RTD.adress_7_N_1086_7_cascade_ ));
    InMux I__1959 (
            .O(N__20496),
            .I(N__20491));
    InMux I__1958 (
            .O(N__20495),
            .I(N__20488));
    InMux I__1957 (
            .O(N__20494),
            .I(N__20485));
    LocalMux I__1956 (
            .O(N__20491),
            .I(N__20482));
    LocalMux I__1955 (
            .O(N__20488),
            .I(N__20479));
    LocalMux I__1954 (
            .O(N__20485),
            .I(N__20476));
    Span4Mux_h I__1953 (
            .O(N__20482),
            .I(N__20469));
    Span4Mux_h I__1952 (
            .O(N__20479),
            .I(N__20469));
    Span4Mux_v I__1951 (
            .O(N__20476),
            .I(N__20469));
    Sp12to4 I__1950 (
            .O(N__20469),
            .I(N__20466));
    Span12Mux_v I__1949 (
            .O(N__20466),
            .I(N__20463));
    Odrv12 I__1948 (
            .O(N__20463),
            .I(RTD_DRDY));
    CascadeMux I__1947 (
            .O(N__20460),
            .I(\RTD.n11_cascade_ ));
    CascadeMux I__1946 (
            .O(N__20457),
            .I(\RTD.n19_cascade_ ));
    CascadeMux I__1945 (
            .O(N__20454),
            .I(N__20451));
    InMux I__1944 (
            .O(N__20451),
            .I(N__20447));
    CascadeMux I__1943 (
            .O(N__20450),
            .I(N__20444));
    LocalMux I__1942 (
            .O(N__20447),
            .I(N__20441));
    InMux I__1941 (
            .O(N__20444),
            .I(N__20438));
    Span4Mux_v I__1940 (
            .O(N__20441),
            .I(N__20435));
    LocalMux I__1939 (
            .O(N__20438),
            .I(\RTD.adress_7 ));
    Odrv4 I__1938 (
            .O(N__20435),
            .I(\RTD.adress_7 ));
    InMux I__1937 (
            .O(N__20430),
            .I(N__20424));
    InMux I__1936 (
            .O(N__20429),
            .I(N__20419));
    InMux I__1935 (
            .O(N__20428),
            .I(N__20419));
    InMux I__1934 (
            .O(N__20427),
            .I(N__20416));
    LocalMux I__1933 (
            .O(N__20424),
            .I(\RTD.adress_7_N_1086_7 ));
    LocalMux I__1932 (
            .O(N__20419),
            .I(\RTD.adress_7_N_1086_7 ));
    LocalMux I__1931 (
            .O(N__20416),
            .I(\RTD.adress_7_N_1086_7 ));
    CascadeMux I__1930 (
            .O(N__20409),
            .I(N__20406));
    InMux I__1929 (
            .O(N__20406),
            .I(N__20403));
    LocalMux I__1928 (
            .O(N__20403),
            .I(N__20400));
    Odrv4 I__1927 (
            .O(N__20400),
            .I(adress_0));
    CEMux I__1926 (
            .O(N__20397),
            .I(N__20394));
    LocalMux I__1925 (
            .O(N__20394),
            .I(N__20385));
    InMux I__1924 (
            .O(N__20393),
            .I(N__20372));
    InMux I__1923 (
            .O(N__20392),
            .I(N__20372));
    InMux I__1922 (
            .O(N__20391),
            .I(N__20372));
    InMux I__1921 (
            .O(N__20390),
            .I(N__20372));
    InMux I__1920 (
            .O(N__20389),
            .I(N__20372));
    InMux I__1919 (
            .O(N__20388),
            .I(N__20372));
    Odrv4 I__1918 (
            .O(N__20385),
            .I(n13054));
    LocalMux I__1917 (
            .O(N__20372),
            .I(n13054));
    CascadeMux I__1916 (
            .O(N__20367),
            .I(\ADC_VAC.n21157_cascade_ ));
    InMux I__1915 (
            .O(N__20364),
            .I(N__20361));
    LocalMux I__1914 (
            .O(N__20361),
            .I(\ADC_VAC.n21468 ));
    CEMux I__1913 (
            .O(N__20358),
            .I(N__20355));
    LocalMux I__1912 (
            .O(N__20355),
            .I(N__20352));
    Span4Mux_v I__1911 (
            .O(N__20352),
            .I(N__20349));
    Odrv4 I__1910 (
            .O(N__20349),
            .I(\ADC_VAC.n21158 ));
    CascadeMux I__1909 (
            .O(N__20346),
            .I(N__20342));
    InMux I__1908 (
            .O(N__20345),
            .I(N__20339));
    InMux I__1907 (
            .O(N__20342),
            .I(N__20336));
    LocalMux I__1906 (
            .O(N__20339),
            .I(N__20333));
    LocalMux I__1905 (
            .O(N__20336),
            .I(N__20330));
    Span4Mux_h I__1904 (
            .O(N__20333),
            .I(N__20327));
    Odrv4 I__1903 (
            .O(N__20330),
            .I(\RTD.n16766 ));
    Odrv4 I__1902 (
            .O(N__20327),
            .I(\RTD.n16766 ));
    IoInMux I__1901 (
            .O(N__20322),
            .I(N__20319));
    LocalMux I__1900 (
            .O(N__20319),
            .I(N__20316));
    IoSpan4Mux I__1899 (
            .O(N__20316),
            .I(N__20313));
    IoSpan4Mux I__1898 (
            .O(N__20313),
            .I(N__20310));
    Span4Mux_s3_h I__1897 (
            .O(N__20310),
            .I(N__20307));
    Span4Mux_v I__1896 (
            .O(N__20307),
            .I(N__20304));
    Span4Mux_h I__1895 (
            .O(N__20304),
            .I(N__20301));
    Odrv4 I__1894 (
            .O(N__20301),
            .I(RTD_CS));
    InMux I__1893 (
            .O(N__20298),
            .I(N__20295));
    LocalMux I__1892 (
            .O(N__20295),
            .I(N__20292));
    Span4Mux_h I__1891 (
            .O(N__20292),
            .I(N__20289));
    Odrv4 I__1890 (
            .O(N__20289),
            .I(\RTD.n14 ));
    CascadeMux I__1889 (
            .O(N__20286),
            .I(\RTD.n21181_cascade_ ));
    CascadeMux I__1888 (
            .O(N__20283),
            .I(\RTD.n13137_cascade_ ));
    InMux I__1887 (
            .O(N__20280),
            .I(N__20276));
    InMux I__1886 (
            .O(N__20279),
            .I(N__20273));
    LocalMux I__1885 (
            .O(N__20276),
            .I(N__20268));
    LocalMux I__1884 (
            .O(N__20273),
            .I(N__20268));
    Span4Mux_v I__1883 (
            .O(N__20268),
            .I(N__20265));
    Odrv4 I__1882 (
            .O(N__20265),
            .I(\RTD.n7889 ));
    InMux I__1881 (
            .O(N__20262),
            .I(\ADC_VAC.n19838 ));
    InMux I__1880 (
            .O(N__20259),
            .I(\ADC_VAC.n19839 ));
    InMux I__1879 (
            .O(N__20256),
            .I(\ADC_VAC.n19840 ));
    InMux I__1878 (
            .O(N__20253),
            .I(\ADC_VAC.n19841 ));
    InMux I__1877 (
            .O(N__20250),
            .I(N__20246));
    InMux I__1876 (
            .O(N__20249),
            .I(N__20243));
    LocalMux I__1875 (
            .O(N__20246),
            .I(\ADC_VAC.bit_cnt_4 ));
    LocalMux I__1874 (
            .O(N__20243),
            .I(\ADC_VAC.bit_cnt_4 ));
    InMux I__1873 (
            .O(N__20238),
            .I(N__20234));
    InMux I__1872 (
            .O(N__20237),
            .I(N__20231));
    LocalMux I__1871 (
            .O(N__20234),
            .I(\ADC_VAC.bit_cnt_3 ));
    LocalMux I__1870 (
            .O(N__20231),
            .I(\ADC_VAC.bit_cnt_3 ));
    CascadeMux I__1869 (
            .O(N__20226),
            .I(N__20222));
    InMux I__1868 (
            .O(N__20225),
            .I(N__20219));
    InMux I__1867 (
            .O(N__20222),
            .I(N__20216));
    LocalMux I__1866 (
            .O(N__20219),
            .I(\ADC_VAC.bit_cnt_1 ));
    LocalMux I__1865 (
            .O(N__20216),
            .I(\ADC_VAC.bit_cnt_1 ));
    InMux I__1864 (
            .O(N__20211),
            .I(N__20207));
    InMux I__1863 (
            .O(N__20210),
            .I(N__20204));
    LocalMux I__1862 (
            .O(N__20207),
            .I(\ADC_VAC.bit_cnt_2 ));
    LocalMux I__1861 (
            .O(N__20204),
            .I(\ADC_VAC.bit_cnt_2 ));
    InMux I__1860 (
            .O(N__20199),
            .I(N__20195));
    InMux I__1859 (
            .O(N__20198),
            .I(N__20192));
    LocalMux I__1858 (
            .O(N__20195),
            .I(N__20189));
    LocalMux I__1857 (
            .O(N__20192),
            .I(\ADC_VAC.bit_cnt_6 ));
    Odrv4 I__1856 (
            .O(N__20189),
            .I(\ADC_VAC.bit_cnt_6 ));
    InMux I__1855 (
            .O(N__20184),
            .I(N__20180));
    InMux I__1854 (
            .O(N__20183),
            .I(N__20177));
    LocalMux I__1853 (
            .O(N__20180),
            .I(\ADC_VAC.bit_cnt_0 ));
    LocalMux I__1852 (
            .O(N__20177),
            .I(\ADC_VAC.bit_cnt_0 ));
    CascadeMux I__1851 (
            .O(N__20172),
            .I(\ADC_VAC.n21224_cascade_ ));
    InMux I__1850 (
            .O(N__20169),
            .I(N__20165));
    InMux I__1849 (
            .O(N__20168),
            .I(N__20162));
    LocalMux I__1848 (
            .O(N__20165),
            .I(\ADC_VAC.bit_cnt_7 ));
    LocalMux I__1847 (
            .O(N__20162),
            .I(\ADC_VAC.bit_cnt_7 ));
    InMux I__1846 (
            .O(N__20157),
            .I(N__20153));
    InMux I__1845 (
            .O(N__20156),
            .I(N__20150));
    LocalMux I__1844 (
            .O(N__20153),
            .I(\ADC_VAC.bit_cnt_5 ));
    LocalMux I__1843 (
            .O(N__20150),
            .I(\ADC_VAC.bit_cnt_5 ));
    CascadeMux I__1842 (
            .O(N__20145),
            .I(\ADC_VAC.n21234_cascade_ ));
    CEMux I__1841 (
            .O(N__20142),
            .I(N__20139));
    LocalMux I__1840 (
            .O(N__20139),
            .I(N__20135));
    InMux I__1839 (
            .O(N__20138),
            .I(N__20132));
    Sp12to4 I__1838 (
            .O(N__20135),
            .I(N__20127));
    LocalMux I__1837 (
            .O(N__20132),
            .I(N__20127));
    Odrv12 I__1836 (
            .O(N__20127),
            .I(\ADC_VAC.n12803 ));
    SRMux I__1835 (
            .O(N__20124),
            .I(N__20121));
    LocalMux I__1834 (
            .O(N__20121),
            .I(N__20118));
    Span4Mux_h I__1833 (
            .O(N__20118),
            .I(N__20115));
    Odrv4 I__1832 (
            .O(N__20115),
            .I(\ADC_VAC.n15052 ));
    InMux I__1831 (
            .O(N__20112),
            .I(N__20106));
    InMux I__1830 (
            .O(N__20111),
            .I(N__20106));
    LocalMux I__1829 (
            .O(N__20106),
            .I(cmd_rdadctmp_7_adj_1485));
    CascadeMux I__1828 (
            .O(N__20103),
            .I(N__20100));
    InMux I__1827 (
            .O(N__20100),
            .I(N__20097));
    LocalMux I__1826 (
            .O(N__20097),
            .I(N__20094));
    Span4Mux_v I__1825 (
            .O(N__20094),
            .I(N__20091));
    Sp12to4 I__1824 (
            .O(N__20091),
            .I(N__20088));
    Odrv12 I__1823 (
            .O(N__20088),
            .I(VAC_MISO));
    InMux I__1822 (
            .O(N__20085),
            .I(N__20079));
    InMux I__1821 (
            .O(N__20084),
            .I(N__20079));
    LocalMux I__1820 (
            .O(N__20079),
            .I(cmd_rdadctmp_0_adj_1492));
    CascadeMux I__1819 (
            .O(N__20076),
            .I(N__20073));
    InMux I__1818 (
            .O(N__20073),
            .I(N__20067));
    InMux I__1817 (
            .O(N__20072),
            .I(N__20067));
    LocalMux I__1816 (
            .O(N__20067),
            .I(cmd_rdadctmp_1_adj_1491));
    InMux I__1815 (
            .O(N__20064),
            .I(N__20058));
    InMux I__1814 (
            .O(N__20063),
            .I(N__20058));
    LocalMux I__1813 (
            .O(N__20058),
            .I(cmd_rdadctmp_2_adj_1490));
    InMux I__1812 (
            .O(N__20055),
            .I(bfn_5_14_0_));
    InMux I__1811 (
            .O(N__20052),
            .I(\ADC_VAC.n19835 ));
    InMux I__1810 (
            .O(N__20049),
            .I(\ADC_VAC.n19836 ));
    InMux I__1809 (
            .O(N__20046),
            .I(\ADC_VAC.n19837 ));
    CascadeMux I__1808 (
            .O(N__20043),
            .I(n19_adj_1597_cascade_));
    InMux I__1807 (
            .O(N__20040),
            .I(N__20037));
    LocalMux I__1806 (
            .O(N__20037),
            .I(N__20034));
    Span4Mux_v I__1805 (
            .O(N__20034),
            .I(N__20029));
    InMux I__1804 (
            .O(N__20033),
            .I(N__20024));
    InMux I__1803 (
            .O(N__20032),
            .I(N__20024));
    Odrv4 I__1802 (
            .O(N__20029),
            .I(buf_adcdata_vac_7));
    LocalMux I__1801 (
            .O(N__20024),
            .I(buf_adcdata_vac_7));
    CascadeMux I__1800 (
            .O(N__20019),
            .I(N__20014));
    CascadeMux I__1799 (
            .O(N__20018),
            .I(N__20011));
    InMux I__1798 (
            .O(N__20017),
            .I(N__20004));
    InMux I__1797 (
            .O(N__20014),
            .I(N__20004));
    InMux I__1796 (
            .O(N__20011),
            .I(N__20004));
    LocalMux I__1795 (
            .O(N__20004),
            .I(read_buf_4));
    CascadeMux I__1794 (
            .O(N__20001),
            .I(N__19996));
    CascadeMux I__1793 (
            .O(N__20000),
            .I(N__19993));
    InMux I__1792 (
            .O(N__19999),
            .I(N__19988));
    InMux I__1791 (
            .O(N__19996),
            .I(N__19988));
    InMux I__1790 (
            .O(N__19993),
            .I(N__19985));
    LocalMux I__1789 (
            .O(N__19988),
            .I(N__19982));
    LocalMux I__1788 (
            .O(N__19985),
            .I(read_buf_11));
    Odrv4 I__1787 (
            .O(N__19982),
            .I(read_buf_11));
    InMux I__1786 (
            .O(N__19977),
            .I(N__19974));
    LocalMux I__1785 (
            .O(N__19974),
            .I(N__19969));
    InMux I__1784 (
            .O(N__19973),
            .I(N__19964));
    InMux I__1783 (
            .O(N__19972),
            .I(N__19964));
    Odrv12 I__1782 (
            .O(N__19969),
            .I(read_buf_5));
    LocalMux I__1781 (
            .O(N__19964),
            .I(read_buf_5));
    CascadeMux I__1780 (
            .O(N__19959),
            .I(N__19955));
    CascadeMux I__1779 (
            .O(N__19958),
            .I(N__19951));
    InMux I__1778 (
            .O(N__19955),
            .I(N__19948));
    InMux I__1777 (
            .O(N__19954),
            .I(N__19943));
    InMux I__1776 (
            .O(N__19951),
            .I(N__19943));
    LocalMux I__1775 (
            .O(N__19948),
            .I(read_buf_3));
    LocalMux I__1774 (
            .O(N__19943),
            .I(read_buf_3));
    CascadeMux I__1773 (
            .O(N__19938),
            .I(n19_adj_1600_cascade_));
    InMux I__1772 (
            .O(N__19935),
            .I(N__19932));
    LocalMux I__1771 (
            .O(N__19932),
            .I(N__19927));
    InMux I__1770 (
            .O(N__19931),
            .I(N__19922));
    InMux I__1769 (
            .O(N__19930),
            .I(N__19922));
    Odrv12 I__1768 (
            .O(N__19927),
            .I(read_buf_10));
    LocalMux I__1767 (
            .O(N__19922),
            .I(read_buf_10));
    CascadeMux I__1766 (
            .O(N__19917),
            .I(n13212_cascade_));
    CascadeMux I__1765 (
            .O(N__19914),
            .I(N__19911));
    InMux I__1764 (
            .O(N__19911),
            .I(N__19905));
    InMux I__1763 (
            .O(N__19910),
            .I(N__19905));
    LocalMux I__1762 (
            .O(N__19905),
            .I(read_buf_15));
    CascadeMux I__1761 (
            .O(N__19902),
            .I(n11856_cascade_));
    CascadeMux I__1760 (
            .O(N__19899),
            .I(N__19894));
    InMux I__1759 (
            .O(N__19898),
            .I(N__19889));
    InMux I__1758 (
            .O(N__19897),
            .I(N__19889));
    InMux I__1757 (
            .O(N__19894),
            .I(N__19886));
    LocalMux I__1756 (
            .O(N__19889),
            .I(read_buf_14));
    LocalMux I__1755 (
            .O(N__19886),
            .I(read_buf_14));
    InMux I__1754 (
            .O(N__19881),
            .I(N__19878));
    LocalMux I__1753 (
            .O(N__19878),
            .I(N__19875));
    Odrv4 I__1752 (
            .O(N__19875),
            .I(\RTD.n12_adj_1445 ));
    CascadeMux I__1751 (
            .O(N__19872),
            .I(N__19869));
    InMux I__1750 (
            .O(N__19869),
            .I(N__19863));
    InMux I__1749 (
            .O(N__19868),
            .I(N__19858));
    InMux I__1748 (
            .O(N__19867),
            .I(N__19858));
    InMux I__1747 (
            .O(N__19866),
            .I(N__19855));
    LocalMux I__1746 (
            .O(N__19863),
            .I(N__19852));
    LocalMux I__1745 (
            .O(N__19858),
            .I(N__19847));
    LocalMux I__1744 (
            .O(N__19855),
            .I(N__19847));
    Span4Mux_h I__1743 (
            .O(N__19852),
            .I(N__19844));
    Odrv4 I__1742 (
            .O(N__19847),
            .I(\RTD.mode ));
    Odrv4 I__1741 (
            .O(N__19844),
            .I(\RTD.mode ));
    InMux I__1740 (
            .O(N__19839),
            .I(N__19833));
    InMux I__1739 (
            .O(N__19838),
            .I(N__19833));
    LocalMux I__1738 (
            .O(N__19833),
            .I(adress_5));
    CascadeMux I__1737 (
            .O(N__19830),
            .I(N__19827));
    InMux I__1736 (
            .O(N__19827),
            .I(N__19824));
    LocalMux I__1735 (
            .O(N__19824),
            .I(N__19821));
    Span4Mux_v I__1734 (
            .O(N__19821),
            .I(N__19818));
    Span4Mux_v I__1733 (
            .O(N__19818),
            .I(N__19815));
    Span4Mux_v I__1732 (
            .O(N__19815),
            .I(N__19812));
    Sp12to4 I__1731 (
            .O(N__19812),
            .I(N__19809));
    Odrv12 I__1730 (
            .O(N__19809),
            .I(RTD_SDO));
    CEMux I__1729 (
            .O(N__19806),
            .I(N__19803));
    LocalMux I__1728 (
            .O(N__19803),
            .I(N__19800));
    Odrv12 I__1727 (
            .O(N__19800),
            .I(\RTD.n11915 ));
    CascadeMux I__1726 (
            .O(N__19797),
            .I(N__19792));
    CascadeMux I__1725 (
            .O(N__19796),
            .I(N__19789));
    InMux I__1724 (
            .O(N__19795),
            .I(N__19783));
    InMux I__1723 (
            .O(N__19792),
            .I(N__19772));
    InMux I__1722 (
            .O(N__19789),
            .I(N__19772));
    InMux I__1721 (
            .O(N__19788),
            .I(N__19772));
    InMux I__1720 (
            .O(N__19787),
            .I(N__19772));
    InMux I__1719 (
            .O(N__19786),
            .I(N__19772));
    LocalMux I__1718 (
            .O(N__19783),
            .I(n14692));
    LocalMux I__1717 (
            .O(N__19772),
            .I(n14692));
    SRMux I__1716 (
            .O(N__19767),
            .I(N__19764));
    LocalMux I__1715 (
            .O(N__19764),
            .I(N__19761));
    Odrv4 I__1714 (
            .O(N__19761),
            .I(\RTD.n15280 ));
    CEMux I__1713 (
            .O(N__19758),
            .I(N__19755));
    LocalMux I__1712 (
            .O(N__19755),
            .I(N__19752));
    Span12Mux_v I__1711 (
            .O(N__19752),
            .I(N__19749));
    Odrv12 I__1710 (
            .O(N__19749),
            .I(\RTD.n11860 ));
    CEMux I__1709 (
            .O(N__19746),
            .I(N__19743));
    LocalMux I__1708 (
            .O(N__19743),
            .I(N__19740));
    Odrv4 I__1707 (
            .O(N__19740),
            .I(\RTD.n8 ));
    CascadeMux I__1706 (
            .O(N__19737),
            .I(N__19734));
    InMux I__1705 (
            .O(N__19734),
            .I(N__19730));
    InMux I__1704 (
            .O(N__19733),
            .I(N__19727));
    LocalMux I__1703 (
            .O(N__19730),
            .I(adress_1));
    LocalMux I__1702 (
            .O(N__19727),
            .I(adress_1));
    CascadeMux I__1701 (
            .O(N__19722),
            .I(N__19719));
    InMux I__1700 (
            .O(N__19719),
            .I(N__19713));
    InMux I__1699 (
            .O(N__19718),
            .I(N__19713));
    LocalMux I__1698 (
            .O(N__19713),
            .I(N__19710));
    Odrv4 I__1697 (
            .O(N__19710),
            .I(adress_2));
    InMux I__1696 (
            .O(N__19707),
            .I(N__19701));
    InMux I__1695 (
            .O(N__19706),
            .I(N__19701));
    LocalMux I__1694 (
            .O(N__19701),
            .I(adress_3));
    CascadeMux I__1693 (
            .O(N__19698),
            .I(N__19695));
    InMux I__1692 (
            .O(N__19695),
            .I(N__19689));
    InMux I__1691 (
            .O(N__19694),
            .I(N__19689));
    LocalMux I__1690 (
            .O(N__19689),
            .I(adress_4));
    CascadeMux I__1689 (
            .O(N__19686),
            .I(N__19683));
    InMux I__1688 (
            .O(N__19683),
            .I(N__19680));
    LocalMux I__1687 (
            .O(N__19680),
            .I(\RTD.n19032 ));
    CascadeMux I__1686 (
            .O(N__19677),
            .I(\RTD.n4_cascade_ ));
    InMux I__1685 (
            .O(N__19674),
            .I(N__19671));
    LocalMux I__1684 (
            .O(N__19671),
            .I(\RTD.n21387 ));
    CascadeMux I__1683 (
            .O(N__19668),
            .I(\RTD.n21199_cascade_ ));
    InMux I__1682 (
            .O(N__19665),
            .I(N__19662));
    LocalMux I__1681 (
            .O(N__19662),
            .I(N__19658));
    InMux I__1680 (
            .O(N__19661),
            .I(N__19655));
    Odrv4 I__1679 (
            .O(N__19658),
            .I(\RTD.adc_state_3_N_1114_1 ));
    LocalMux I__1678 (
            .O(N__19655),
            .I(\RTD.adc_state_3_N_1114_1 ));
    CascadeMux I__1677 (
            .O(N__19650),
            .I(\RTD.n7_cascade_ ));
    CEMux I__1676 (
            .O(N__19647),
            .I(N__19644));
    LocalMux I__1675 (
            .O(N__19644),
            .I(N__19640));
    CEMux I__1674 (
            .O(N__19643),
            .I(N__19637));
    Span4Mux_v I__1673 (
            .O(N__19640),
            .I(N__19632));
    LocalMux I__1672 (
            .O(N__19637),
            .I(N__19632));
    Odrv4 I__1671 (
            .O(N__19632),
            .I(\RTD.n11868 ));
    CascadeMux I__1670 (
            .O(N__19629),
            .I(\RTD.n21492_cascade_ ));
    InMux I__1669 (
            .O(N__19626),
            .I(N__19623));
    LocalMux I__1668 (
            .O(N__19623),
            .I(N__19620));
    Odrv4 I__1667 (
            .O(N__19620),
            .I(\RTD.n7_adj_1435 ));
    CascadeMux I__1666 (
            .O(N__19617),
            .I(N__19614));
    InMux I__1665 (
            .O(N__19614),
            .I(N__19607));
    InMux I__1664 (
            .O(N__19613),
            .I(N__19607));
    InMux I__1663 (
            .O(N__19612),
            .I(N__19604));
    LocalMux I__1662 (
            .O(N__19607),
            .I(\RTD.bit_cnt_2 ));
    LocalMux I__1661 (
            .O(N__19604),
            .I(\RTD.bit_cnt_2 ));
    InMux I__1660 (
            .O(N__19599),
            .I(N__19589));
    InMux I__1659 (
            .O(N__19598),
            .I(N__19589));
    InMux I__1658 (
            .O(N__19597),
            .I(N__19589));
    InMux I__1657 (
            .O(N__19596),
            .I(N__19586));
    LocalMux I__1656 (
            .O(N__19589),
            .I(\RTD.bit_cnt_1 ));
    LocalMux I__1655 (
            .O(N__19586),
            .I(\RTD.bit_cnt_1 ));
    InMux I__1654 (
            .O(N__19581),
            .I(N__19568));
    InMux I__1653 (
            .O(N__19580),
            .I(N__19568));
    InMux I__1652 (
            .O(N__19579),
            .I(N__19568));
    InMux I__1651 (
            .O(N__19578),
            .I(N__19568));
    InMux I__1650 (
            .O(N__19577),
            .I(N__19565));
    LocalMux I__1649 (
            .O(N__19568),
            .I(\RTD.bit_cnt_0 ));
    LocalMux I__1648 (
            .O(N__19565),
            .I(\RTD.bit_cnt_0 ));
    IoInMux I__1647 (
            .O(N__19560),
            .I(N__19557));
    LocalMux I__1646 (
            .O(N__19557),
            .I(N__19554));
    Span4Mux_s2_h I__1645 (
            .O(N__19554),
            .I(N__19551));
    Sp12to4 I__1644 (
            .O(N__19551),
            .I(N__19548));
    Span12Mux_v I__1643 (
            .O(N__19548),
            .I(N__19545));
    Odrv12 I__1642 (
            .O(N__19545),
            .I(RTD_SDI));
    CascadeMux I__1641 (
            .O(N__19542),
            .I(\RTD.n21471_cascade_ ));
    IoInMux I__1640 (
            .O(N__19539),
            .I(N__19536));
    LocalMux I__1639 (
            .O(N__19536),
            .I(N__19533));
    IoSpan4Mux I__1638 (
            .O(N__19533),
            .I(N__19530));
    Span4Mux_s3_h I__1637 (
            .O(N__19530),
            .I(N__19527));
    Span4Mux_v I__1636 (
            .O(N__19527),
            .I(N__19524));
    Span4Mux_v I__1635 (
            .O(N__19524),
            .I(N__19521));
    Odrv4 I__1634 (
            .O(N__19521),
            .I(RTD_SCLK));
    SRMux I__1633 (
            .O(N__19518),
            .I(N__19515));
    LocalMux I__1632 (
            .O(N__19515),
            .I(\CLK_DDS.n16974 ));
    InMux I__1631 (
            .O(N__19512),
            .I(N__19501));
    InMux I__1630 (
            .O(N__19511),
            .I(N__19501));
    InMux I__1629 (
            .O(N__19510),
            .I(N__19501));
    InMux I__1628 (
            .O(N__19509),
            .I(N__19496));
    InMux I__1627 (
            .O(N__19508),
            .I(N__19496));
    LocalMux I__1626 (
            .O(N__19501),
            .I(bit_cnt_0_adj_1498));
    LocalMux I__1625 (
            .O(N__19496),
            .I(bit_cnt_0_adj_1498));
    InMux I__1624 (
            .O(N__19491),
            .I(N__19487));
    InMux I__1623 (
            .O(N__19490),
            .I(N__19484));
    LocalMux I__1622 (
            .O(N__19487),
            .I(bit_cnt_3));
    LocalMux I__1621 (
            .O(N__19484),
            .I(bit_cnt_3));
    InMux I__1620 (
            .O(N__19479),
            .I(N__19474));
    InMux I__1619 (
            .O(N__19478),
            .I(N__19471));
    InMux I__1618 (
            .O(N__19477),
            .I(N__19468));
    LocalMux I__1617 (
            .O(N__19474),
            .I(bit_cnt_2));
    LocalMux I__1616 (
            .O(N__19471),
            .I(bit_cnt_2));
    LocalMux I__1615 (
            .O(N__19468),
            .I(bit_cnt_2));
    CascadeMux I__1614 (
            .O(N__19461),
            .I(N__19458));
    InMux I__1613 (
            .O(N__19458),
            .I(N__19450));
    InMux I__1612 (
            .O(N__19457),
            .I(N__19450));
    InMux I__1611 (
            .O(N__19456),
            .I(N__19447));
    InMux I__1610 (
            .O(N__19455),
            .I(N__19444));
    LocalMux I__1609 (
            .O(N__19450),
            .I(bit_cnt_1));
    LocalMux I__1608 (
            .O(N__19447),
            .I(bit_cnt_1));
    LocalMux I__1607 (
            .O(N__19444),
            .I(bit_cnt_1));
    CascadeMux I__1606 (
            .O(N__19437),
            .I(n8_adj_1680_cascade_));
    InMux I__1605 (
            .O(N__19434),
            .I(N__19431));
    LocalMux I__1604 (
            .O(N__19431),
            .I(n21625));
    CascadeMux I__1603 (
            .O(N__19428),
            .I(\RTD.n18043_cascade_ ));
    InMux I__1602 (
            .O(N__19425),
            .I(N__19422));
    LocalMux I__1601 (
            .O(N__19422),
            .I(\RTD.n21494 ));
    InMux I__1600 (
            .O(N__19419),
            .I(N__19416));
    LocalMux I__1599 (
            .O(N__19416),
            .I(\RTD.n18092 ));
    IoInMux I__1598 (
            .O(N__19413),
            .I(N__19410));
    LocalMux I__1597 (
            .O(N__19410),
            .I(N__19407));
    IoSpan4Mux I__1596 (
            .O(N__19407),
            .I(N__19404));
    IoSpan4Mux I__1595 (
            .O(N__19404),
            .I(N__19401));
    Odrv4 I__1594 (
            .O(N__19401),
            .I(ICE_SYSCLK));
    IoInMux I__1593 (
            .O(N__19398),
            .I(N__19395));
    LocalMux I__1592 (
            .O(N__19395),
            .I(N__19392));
    IoSpan4Mux I__1591 (
            .O(N__19392),
            .I(N__19389));
    Span4Mux_s3_v I__1590 (
            .O(N__19389),
            .I(N__19386));
    Sp12to4 I__1589 (
            .O(N__19386),
            .I(N__19383));
    Span12Mux_h I__1588 (
            .O(N__19383),
            .I(N__19380));
    Odrv12 I__1587 (
            .O(N__19380),
            .I(ICE_GPMO_2));
    INV \INVADC_VDC.genclk.t0on_i8C  (
            .O(\INVADC_VDC.genclk.t0on_i8C_net ),
            .I(N__50798));
    INV \INVADC_VDC.genclk.t0on_i0C  (
            .O(\INVADC_VDC.genclk.t0on_i0C_net ),
            .I(N__50797));
    INV \INVADC_VDC.genclk.div_state_i0C  (
            .O(\INVADC_VDC.genclk.div_state_i0C_net ),
            .I(N__50796));
    INV \INVADC_VDC.genclk.t0off_i8C  (
            .O(\INVADC_VDC.genclk.t0off_i8C_net ),
            .I(N__50795));
    INV \INVADC_VDC.genclk.t0off_i0C  (
            .O(\INVADC_VDC.genclk.t0off_i0C_net ),
            .I(N__50794));
    INV \INVADC_VDC.genclk.div_state_i1C  (
            .O(\INVADC_VDC.genclk.div_state_i1C_net ),
            .I(N__50793));
    INV INVdds0_mclkcnt_i7_3772__i0C (
            .O(INVdds0_mclkcnt_i7_3772__i0C_net),
            .I(N__50803));
    INV INVdds0_mclk_294C (
            .O(INVdds0_mclk_294C_net),
            .I(N__50799));
    INV \INVcomm_spi.data_valid_85C  (
            .O(\INVcomm_spi.data_valid_85C_net ),
            .I(N__55969));
    INV \INVcomm_spi.MISO_48_12291_12292_setC  (
            .O(\INVcomm_spi.MISO_48_12291_12292_setC_net ),
            .I(N__55941));
    INV \INVcomm_spi.MISO_48_12291_12292_resetC  (
            .O(\INVcomm_spi.MISO_48_12291_12292_resetC_net ),
            .I(N__55939));
    INV \INVcomm_spi.imiso_83_12297_12298_setC  (
            .O(\INVcomm_spi.imiso_83_12297_12298_setC_net ),
            .I(N__58307));
    INV INVdata_cntvec_i0_i8C (
            .O(INVdata_cntvec_i0_i8C_net),
            .I(N__56006));
    INV INVdata_cntvec_i0_i0C (
            .O(INVdata_cntvec_i0_i0C_net),
            .I(N__55992));
    INV \INVcomm_spi.bit_cnt_3767__i3C  (
            .O(\INVcomm_spi.bit_cnt_3767__i3C_net ),
            .I(N__58391));
    INV \INVADC_VDC.genclk.t_clk_24C  (
            .O(\INVADC_VDC.genclk.t_clk_24C_net ),
            .I(N__50781));
    INV \INVcomm_spi.imiso_83_12297_12298_resetC  (
            .O(\INVcomm_spi.imiso_83_12297_12298_resetC_net ),
            .I(N__58357));
    INV INVacadc_skipcnt_i0_i9C (
            .O(INVacadc_skipcnt_i0_i9C_net),
            .I(N__56078));
    INV INVacadc_skipcnt_i0_i1C (
            .O(INVacadc_skipcnt_i0_i1C_net),
            .I(N__56065));
    INV INVacadc_skipcnt_i0_i0C (
            .O(INVacadc_skipcnt_i0_i0C_net),
            .I(N__56052));
    INV INVdata_count_i0_i8C (
            .O(INVdata_count_i0_i8C_net),
            .I(N__56045));
    INV INVdata_count_i0_i0C (
            .O(INVdata_count_i0_i0C_net),
            .I(N__56029));
    INV INVeis_state_i0C (
            .O(INVeis_state_i0C_net),
            .I(N__55990));
    INV INVeis_state_i1C (
            .O(INVeis_state_i1C_net),
            .I(N__56020));
    INV INVacadc_trig_300C (
            .O(INVacadc_trig_300C_net),
            .I(N__56003));
    INV INViac_raw_buf_vac_raw_buf_merged2WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged2WCLKN_net),
            .I(N__56043));
    INV INViac_raw_buf_vac_raw_buf_merged7WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged7WCLKN_net),
            .I(N__56103));
    INV INViac_raw_buf_vac_raw_buf_merged1WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged1WCLKN_net),
            .I(N__55961));
    INV INViac_raw_buf_vac_raw_buf_merged6WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged6WCLKN_net),
            .I(N__56101));
    INV INViac_raw_buf_vac_raw_buf_merged0WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged0WCLKN_net),
            .I(N__55949));
    INV INViac_raw_buf_vac_raw_buf_merged5WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged5WCLKN_net),
            .I(N__56098));
    INV INViac_raw_buf_vac_raw_buf_merged9WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged9WCLKN_net),
            .I(N__55998));
    INV INViac_raw_buf_vac_raw_buf_merged4WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged4WCLKN_net),
            .I(N__56091));
    INV INViac_raw_buf_vac_raw_buf_merged8WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged8WCLKN_net),
            .I(N__55973));
    INV INViac_raw_buf_vac_raw_buf_merged10WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged10WCLKN_net),
            .I(N__55985));
    INV INViac_raw_buf_vac_raw_buf_merged3WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged3WCLKN_net),
            .I(N__56072));
    INV INViac_raw_buf_vac_raw_buf_merged11WCLKN (
            .O(INViac_raw_buf_vac_raw_buf_merged11WCLKN_net),
            .I(N__56013));
    defparam IN_MUX_bfv_15_5_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_15_5_0_));
    defparam IN_MUX_bfv_15_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_6_0_ (
            .carryinitin(n19939),
            .carryinitout(bfn_15_6_0_));
    defparam IN_MUX_bfv_15_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_7_0_ (
            .carryinitin(n19947),
            .carryinitout(bfn_15_7_0_));
    defparam IN_MUX_bfv_15_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_15_8_0_ (
            .carryinitin(n19955),
            .carryinitout(bfn_15_8_0_));
    defparam IN_MUX_bfv_11_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_7_0_));
    defparam IN_MUX_bfv_11_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_8_0_ (
            .carryinitin(n19963),
            .carryinitout(bfn_11_8_0_));
    defparam IN_MUX_bfv_11_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_9_0_ (
            .carryinitin(n19971),
            .carryinitout(bfn_11_9_0_));
    defparam IN_MUX_bfv_18_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_16_0_));
    defparam IN_MUX_bfv_13_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_18_0_));
    defparam IN_MUX_bfv_13_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_19_0_ (
            .carryinitin(n19789_THRU_CRY_6_THRU_CO),
            .carryinitout(bfn_13_19_0_));
    defparam IN_MUX_bfv_13_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_20_0_ (
            .carryinitin(n19797),
            .carryinitout(bfn_13_20_0_));
    defparam IN_MUX_bfv_14_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_13_0_));
    defparam IN_MUX_bfv_14_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_14_0_ (
            .carryinitin(n19781),
            .carryinitout(bfn_14_14_0_));
    defparam IN_MUX_bfv_12_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_18_0_));
    defparam IN_MUX_bfv_12_19_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_19_0_ (
            .carryinitin(n19772),
            .carryinitout(bfn_12_19_0_));
    defparam IN_MUX_bfv_9_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_11_0_));
    defparam IN_MUX_bfv_9_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_12_0_ (
            .carryinitin(n19820),
            .carryinitout(bfn_9_12_0_));
    defparam IN_MUX_bfv_14_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_15_0_));
    defparam IN_MUX_bfv_14_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_16_0_ (
            .carryinitin(n19811),
            .carryinitout(bfn_14_16_0_));
    defparam IN_MUX_bfv_19_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_19_7_0_));
    defparam IN_MUX_bfv_19_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_19_8_0_ (
            .carryinitin(\ADC_VDC.genclk.n19895 ),
            .carryinitout(bfn_19_8_0_));
    defparam IN_MUX_bfv_22_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_22_7_0_));
    defparam IN_MUX_bfv_22_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_22_8_0_ (
            .carryinitin(\ADC_VDC.genclk.n19910 ),
            .carryinitout(bfn_22_8_0_));
    defparam IN_MUX_bfv_13_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_6_0_));
    defparam IN_MUX_bfv_10_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_6_0_));
    defparam IN_MUX_bfv_10_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_7_0_ (
            .carryinitin(\ADC_VDC.n19884 ),
            .carryinitout(bfn_10_7_0_));
    defparam IN_MUX_bfv_8_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_6_0_));
    defparam IN_MUX_bfv_8_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_7_0_ (
            .carryinitin(\ADC_VDC.n19849 ),
            .carryinitout(bfn_8_7_0_));
    defparam IN_MUX_bfv_8_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_8_0_ (
            .carryinitin(\ADC_VDC.n19857 ),
            .carryinitout(bfn_8_8_0_));
    defparam IN_MUX_bfv_8_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_9_0_ (
            .carryinitin(\ADC_VDC.n19865 ),
            .carryinitout(bfn_8_9_0_));
    defparam IN_MUX_bfv_8_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_10_0_ (
            .carryinitin(\ADC_VDC.n19873 ),
            .carryinitout(bfn_8_10_0_));
    defparam IN_MUX_bfv_5_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_14_0_));
    defparam IN_MUX_bfv_6_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_18_0_));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \CLK_DDS.bit_cnt_i3_LC_2_7_0 .C_ON=1'b0;
    defparam \CLK_DDS.bit_cnt_i3_LC_2_7_0 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.bit_cnt_i3_LC_2_7_0 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \CLK_DDS.bit_cnt_i3_LC_2_7_0  (
            .in0(N__19479),
            .in1(N__19512),
            .in2(N__19461),
            .in3(N__19491),
            .lcout(bit_cnt_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56028),
            .ce(N__29821),
            .sr(N__19518));
    defparam \CLK_DDS.bit_cnt_i2_LC_2_7_2 .C_ON=1'b0;
    defparam \CLK_DDS.bit_cnt_i2_LC_2_7_2 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.bit_cnt_i2_LC_2_7_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \CLK_DDS.bit_cnt_i2_LC_2_7_2  (
            .in0(N__19457),
            .in1(N__19478),
            .in2(_gnd_net_),
            .in3(N__19511),
            .lcout(bit_cnt_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56028),
            .ce(N__29821),
            .sr(N__19518));
    defparam \CLK_DDS.bit_cnt_i1_LC_2_7_4 .C_ON=1'b0;
    defparam \CLK_DDS.bit_cnt_i1_LC_2_7_4 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.bit_cnt_i1_LC_2_7_4 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \CLK_DDS.bit_cnt_i1_LC_2_7_4  (
            .in0(_gnd_net_),
            .in1(N__19456),
            .in2(_gnd_net_),
            .in3(N__19510),
            .lcout(bit_cnt_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56028),
            .ce(N__29821),
            .sr(N__19518));
    defparam \RTD.adc_state_3__I_0_66_Mux_0_i14_4_lut_LC_2_8_4 .C_ON=1'b0;
    defparam \RTD.adc_state_3__I_0_66_Mux_0_i14_4_lut_LC_2_8_4 .SEQ_MODE=4'b0000;
    defparam \RTD.adc_state_3__I_0_66_Mux_0_i14_4_lut_LC_2_8_4 .LUT_INIT=16'b1100101011000000;
    LogicCell40 \RTD.adc_state_3__I_0_66_Mux_0_i14_4_lut_LC_2_8_4  (
            .in0(N__22350),
            .in1(N__20279),
            .in2(N__22173),
            .in3(N__19425),
            .lcout(\RTD.n18092 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.dds_state_i2_LC_2_8_7 .C_ON=1'b0;
    defparam \CLK_DDS.dds_state_i2_LC_2_8_7 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.dds_state_i2_LC_2_8_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \CLK_DDS.dds_state_i2_LC_2_8_7  (
            .in0(_gnd_net_),
            .in1(N__30007),
            .in2(_gnd_net_),
            .in3(N__29819),
            .lcout(dds_state_2_adj_1494),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56044),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adc_state_i0_LC_2_9_0 .C_ON=1'b0;
    defparam \RTD.adc_state_i0_LC_2_9_0 .SEQ_MODE=4'b1000;
    defparam \RTD.adc_state_i0_LC_2_9_0 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \RTD.adc_state_i0_LC_2_9_0  (
            .in0(N__22693),
            .in1(N__19419),
            .in2(_gnd_net_),
            .in3(N__19626),
            .lcout(\RTD.adc_state_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40617),
            .ce(N__19647),
            .sr(_gnd_net_));
    defparam \RTD.adc_state_i3_LC_2_9_1 .C_ON=1'b0;
    defparam \RTD.adc_state_i3_LC_2_9_1 .SEQ_MODE=4'b1000;
    defparam \RTD.adc_state_i3_LC_2_9_1 .LUT_INIT=16'b0010001000100111;
    LogicCell40 \RTD.adc_state_i3_LC_2_9_1  (
            .in0(N__22640),
            .in1(N__22111),
            .in2(N__19686),
            .in3(N__20538),
            .lcout(\RTD.adc_state_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40617),
            .ce(N__19647),
            .sr(_gnd_net_));
    defparam \RTD.adc_state_i2_LC_2_9_2 .C_ON=1'b0;
    defparam \RTD.adc_state_i2_LC_2_9_2 .SEQ_MODE=4'b1000;
    defparam \RTD.adc_state_i2_LC_2_9_2 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \RTD.adc_state_i2_LC_2_9_2  (
            .in0(N__19674),
            .in1(N__20280),
            .in2(N__22174),
            .in3(N__22644),
            .lcout(adc_state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40617),
            .ce(N__19647),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_LC_2_9_7.C_ON=1'b0;
    defparam i1_2_lut_3_lut_LC_2_9_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_LC_2_9_7.LUT_INIT=16'b0000000000100010;
    LogicCell40 i1_2_lut_3_lut_LC_2_9_7 (
            .in0(N__52285),
            .in1(N__54857),
            .in2(_gnd_net_),
            .in3(N__54554),
            .lcout(n14_adj_1578),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.SCLK_51_LC_2_10_4 .C_ON=1'b0;
    defparam \RTD.SCLK_51_LC_2_10_4 .SEQ_MODE=4'b1000;
    defparam \RTD.SCLK_51_LC_2_10_4 .LUT_INIT=16'b0000101111010100;
    LogicCell40 \RTD.SCLK_51_LC_2_10_4  (
            .in0(N__22351),
            .in1(N__20725),
            .in2(N__22678),
            .in3(N__22115),
            .lcout(RTD_SCLK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40615),
            .ce(N__19746),
            .sr(_gnd_net_));
    defparam \CLK_DDS.bit_cnt_i0_LC_3_6_2 .C_ON=1'b0;
    defparam \CLK_DDS.bit_cnt_i0_LC_3_6_2 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.bit_cnt_i0_LC_3_6_2 .LUT_INIT=16'b0000010010101010;
    LogicCell40 \CLK_DDS.bit_cnt_i0_LC_3_6_2  (
            .in0(N__19509),
            .in1(N__29910),
            .in2(N__30045),
            .in3(N__29791),
            .lcout(bit_cnt_0_adj_1498),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55996),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.i1_3_lut_LC_3_6_4 .C_ON=1'b0;
    defparam \CLK_DDS.i1_3_lut_LC_3_6_4 .SEQ_MODE=4'b0000;
    defparam \CLK_DDS.i1_3_lut_LC_3_6_4 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \CLK_DDS.i1_3_lut_LC_3_6_4  (
            .in0(N__30016),
            .in1(N__29909),
            .in2(_gnd_net_),
            .in3(N__29790),
            .lcout(\CLK_DDS.n16974 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19325_2_lut_LC_3_6_7.C_ON=1'b0;
    defparam i19325_2_lut_LC_3_6_7.SEQ_MODE=4'b0000;
    defparam i19325_2_lut_LC_3_6_7.LUT_INIT=16'b1100110000000000;
    LogicCell40 i19325_2_lut_LC_3_6_7 (
            .in0(_gnd_net_),
            .in1(N__19508),
            .in2(_gnd_net_),
            .in3(N__19490),
            .lcout(n21625),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.i3_3_lut_4_lut_LC_3_7_0 .C_ON=1'b0;
    defparam \CLK_DDS.i3_3_lut_4_lut_LC_3_7_0 .SEQ_MODE=4'b0000;
    defparam \CLK_DDS.i3_3_lut_4_lut_LC_3_7_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \CLK_DDS.i3_3_lut_4_lut_LC_3_7_0  (
            .in0(N__29907),
            .in1(N__19477),
            .in2(N__30031),
            .in3(N__19455),
            .lcout(),
            .ltout(n8_adj_1680_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.dds_state_i0_LC_3_7_1 .C_ON=1'b0;
    defparam \CLK_DDS.dds_state_i0_LC_3_7_1 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.dds_state_i0_LC_3_7_1 .LUT_INIT=16'b1011000100010001;
    LogicCell40 \CLK_DDS.dds_state_i0_LC_3_7_1  (
            .in0(N__29820),
            .in1(N__29908),
            .in2(N__19437),
            .in3(N__19434),
            .lcout(dds_state_0_adj_1496),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56014),
            .ce(N__29718),
            .sr(_gnd_net_));
    defparam \RTD.i2_3_lut_LC_3_7_3 .C_ON=1'b0;
    defparam \RTD.i2_3_lut_LC_3_7_3 .SEQ_MODE=4'b0000;
    defparam \RTD.i2_3_lut_LC_3_7_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \RTD.i2_3_lut_LC_3_7_3  (
            .in0(N__19612),
            .in1(N__19577),
            .in2(_gnd_net_),
            .in3(N__19596),
            .lcout(\RTD.n18043 ),
            .ltout(\RTD.n18043_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i19370_3_lut_LC_3_7_4 .C_ON=1'b0;
    defparam \RTD.i19370_3_lut_LC_3_7_4 .SEQ_MODE=4'b0000;
    defparam \RTD.i19370_3_lut_LC_3_7_4 .LUT_INIT=16'b1111111101011111;
    LogicCell40 \RTD.i19370_3_lut_LC_3_7_4  (
            .in0(N__20580),
            .in1(_gnd_net_),
            .in2(N__19428),
            .in3(N__20711),
            .lcout(\RTD.n21494 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i19209_4_lut_LC_3_7_6 .C_ON=1'b0;
    defparam \RTD.i19209_4_lut_LC_3_7_6 .SEQ_MODE=4'b0000;
    defparam \RTD.i19209_4_lut_LC_3_7_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \RTD.i19209_4_lut_LC_3_7_6  (
            .in0(N__20579),
            .in1(N__20712),
            .in2(N__19872),
            .in3(N__20554),
            .lcout(),
            .ltout(\RTD.n21492_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adc_state_3__I_0_66_Mux_0_i7_4_lut_LC_3_7_7 .C_ON=1'b0;
    defparam \RTD.adc_state_3__I_0_66_Mux_0_i7_4_lut_LC_3_7_7 .SEQ_MODE=4'b0000;
    defparam \RTD.adc_state_3__I_0_66_Mux_0_i7_4_lut_LC_3_7_7 .LUT_INIT=16'b0111010100110001;
    LogicCell40 \RTD.adc_state_3__I_0_66_Mux_0_i7_4_lut_LC_3_7_7  (
            .in0(N__22379),
            .in1(N__22169),
            .in2(N__19629),
            .in3(N__20534),
            .lcout(\RTD.n7_adj_1435 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.bit_cnt_3769__i3_LC_3_8_0 .C_ON=1'b0;
    defparam \RTD.bit_cnt_3769__i3_LC_3_8_0 .SEQ_MODE=4'b1000;
    defparam \RTD.bit_cnt_3769__i3_LC_3_8_0 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \RTD.bit_cnt_3769__i3_LC_3_8_0  (
            .in0(N__19599),
            .in1(N__20582),
            .in2(N__19617),
            .in3(N__19581),
            .lcout(\RTD.bit_cnt_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40623),
            .ce(N__19806),
            .sr(N__19767));
    defparam \RTD.bit_cnt_3769__i2_LC_3_8_1 .C_ON=1'b0;
    defparam \RTD.bit_cnt_3769__i2_LC_3_8_1 .SEQ_MODE=4'b1000;
    defparam \RTD.bit_cnt_3769__i2_LC_3_8_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RTD.bit_cnt_3769__i2_LC_3_8_1  (
            .in0(N__19580),
            .in1(N__19613),
            .in2(_gnd_net_),
            .in3(N__19598),
            .lcout(\RTD.bit_cnt_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40623),
            .ce(N__19806),
            .sr(N__19767));
    defparam \RTD.i1_2_lut_LC_3_8_2 .C_ON=1'b0;
    defparam \RTD.i1_2_lut_LC_3_8_2 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_2_lut_LC_3_8_2 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \RTD.i1_2_lut_LC_3_8_2  (
            .in0(N__20555),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20581),
            .lcout(\RTD.adc_state_3_N_1114_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.bit_cnt_3769__i1_LC_3_8_3 .C_ON=1'b0;
    defparam \RTD.bit_cnt_3769__i1_LC_3_8_3 .SEQ_MODE=4'b1000;
    defparam \RTD.bit_cnt_3769__i1_LC_3_8_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \RTD.bit_cnt_3769__i1_LC_3_8_3  (
            .in0(N__19579),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19597),
            .lcout(\RTD.bit_cnt_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40623),
            .ce(N__19806),
            .sr(N__19767));
    defparam \RTD.bit_cnt_3769__i0_LC_3_8_4 .C_ON=1'b0;
    defparam \RTD.bit_cnt_3769__i0_LC_3_8_4 .SEQ_MODE=4'b1000;
    defparam \RTD.bit_cnt_3769__i0_LC_3_8_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \RTD.bit_cnt_3769__i0_LC_3_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19578),
            .lcout(\RTD.bit_cnt_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40623),
            .ce(N__19806),
            .sr(N__19767));
    defparam i15467_2_lut_3_lut_LC_3_8_6.C_ON=1'b0;
    defparam i15467_2_lut_3_lut_LC_3_8_6.SEQ_MODE=4'b0000;
    defparam i15467_2_lut_3_lut_LC_3_8_6.LUT_INIT=16'b0000000000100010;
    LogicCell40 i15467_2_lut_3_lut_LC_3_8_6 (
            .in0(N__45479),
            .in1(N__54893),
            .in2(_gnd_net_),
            .in3(N__54514),
            .lcout(n14_adj_1548),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.MOSI_59_LC_3_9_0 .C_ON=1'b0;
    defparam \RTD.MOSI_59_LC_3_9_0 .SEQ_MODE=4'b1000;
    defparam \RTD.MOSI_59_LC_3_9_0 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \RTD.MOSI_59_LC_3_9_0  (
            .in0(N__22097),
            .in1(N__22343),
            .in2(N__20454),
            .in3(N__22242),
            .lcout(RTD_SDI),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40616),
            .ce(N__19758),
            .sr(N__20810));
    defparam \RTD.i19122_3_lut_LC_3_9_1 .C_ON=1'b0;
    defparam \RTD.i19122_3_lut_LC_3_9_1 .SEQ_MODE=4'b0000;
    defparam \RTD.i19122_3_lut_LC_3_9_1 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \RTD.i19122_3_lut_LC_3_9_1  (
            .in0(N__22339),
            .in1(N__22512),
            .in2(_gnd_net_),
            .in3(N__20494),
            .lcout(),
            .ltout(\RTD.n21471_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_4_lut_adj_10_LC_3_9_2 .C_ON=1'b0;
    defparam \RTD.i1_4_lut_adj_10_LC_3_9_2 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_4_lut_adj_10_LC_3_9_2 .LUT_INIT=16'b0111010000000000;
    LogicCell40 \RTD.i1_4_lut_adj_10_LC_3_9_2  (
            .in0(N__22095),
            .in1(N__22639),
            .in2(N__19542),
            .in3(N__19868),
            .lcout(\RTD.n12_adj_1445 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i16510_3_lut_LC_3_9_3 .C_ON=1'b0;
    defparam \RTD.i16510_3_lut_LC_3_9_3 .SEQ_MODE=4'b0000;
    defparam \RTD.i16510_3_lut_LC_3_9_3 .LUT_INIT=16'b1010101011011101;
    LogicCell40 \RTD.i16510_3_lut_LC_3_9_3  (
            .in0(N__22342),
            .in1(N__19866),
            .in2(_gnd_net_),
            .in3(N__22096),
            .lcout(\RTD.n19032 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i2_3_lut_adj_19_LC_3_9_4 .C_ON=1'b0;
    defparam \RTD.i2_3_lut_adj_19_LC_3_9_4 .SEQ_MODE=4'b0000;
    defparam \RTD.i2_3_lut_adj_19_LC_3_9_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \RTD.i2_3_lut_adj_19_LC_3_9_4  (
            .in0(N__22094),
            .in1(N__22635),
            .in2(_gnd_net_),
            .in3(N__22338),
            .lcout(n1_adj_1592),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_2_lut_adj_4_LC_3_9_5 .C_ON=1'b0;
    defparam \RTD.i1_2_lut_adj_4_LC_3_9_5 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_2_lut_adj_4_LC_3_9_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \RTD.i1_2_lut_adj_4_LC_3_9_5  (
            .in0(N__22341),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20679),
            .lcout(),
            .ltout(\RTD.n4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i19032_4_lut_LC_3_9_6 .C_ON=1'b0;
    defparam \RTD.i19032_4_lut_LC_3_9_6 .SEQ_MODE=4'b0000;
    defparam \RTD.i19032_4_lut_LC_3_9_6 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \RTD.i19032_4_lut_LC_3_9_6  (
            .in0(N__22652),
            .in1(N__19867),
            .in2(N__19677),
            .in3(N__19661),
            .lcout(\RTD.n21387 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_2_lut_adj_21_LC_3_9_7 .C_ON=1'b0;
    defparam \RTD.i1_2_lut_adj_21_LC_3_9_7 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_2_lut_adj_21_LC_3_9_7 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \RTD.i1_2_lut_adj_21_LC_3_9_7  (
            .in0(N__22340),
            .in1(_gnd_net_),
            .in2(N__22677),
            .in3(_gnd_net_),
            .lcout(\RTD.n21061 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i18472_2_lut_LC_3_10_0 .C_ON=1'b0;
    defparam \RTD.i18472_2_lut_LC_3_10_0 .SEQ_MODE=4'b0000;
    defparam \RTD.i18472_2_lut_LC_3_10_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \RTD.i18472_2_lut_LC_3_10_0  (
            .in0(_gnd_net_),
            .in1(N__20671),
            .in2(_gnd_net_),
            .in3(N__22066),
            .lcout(\RTD.n21199 ),
            .ltout(\RTD.n21199_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i3_4_lut_LC_3_10_1 .C_ON=1'b0;
    defparam \RTD.i3_4_lut_LC_3_10_1 .SEQ_MODE=4'b0000;
    defparam \RTD.i3_4_lut_LC_3_10_1 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \RTD.i3_4_lut_LC_3_10_1  (
            .in0(N__22331),
            .in1(N__22605),
            .in2(N__19668),
            .in3(N__20345),
            .lcout(\RTD.n11868 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adc_state_3__I_0_66_Mux_1_i7_4_lut_4_lut_LC_3_10_2 .C_ON=1'b0;
    defparam \RTD.adc_state_3__I_0_66_Mux_1_i7_4_lut_4_lut_LC_3_10_2 .SEQ_MODE=4'b0000;
    defparam \RTD.adc_state_3__I_0_66_Mux_1_i7_4_lut_4_lut_LC_3_10_2 .LUT_INIT=16'b1111011011010110;
    LogicCell40 \RTD.adc_state_3__I_0_66_Mux_1_i7_4_lut_4_lut_LC_3_10_2  (
            .in0(N__20685),
            .in1(N__22336),
            .in2(N__22168),
            .in3(N__19665),
            .lcout(),
            .ltout(\RTD.n7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adc_state_i1_LC_3_10_3 .C_ON=1'b0;
    defparam \RTD.adc_state_i1_LC_3_10_3 .SEQ_MODE=4'b1000;
    defparam \RTD.adc_state_i1_LC_3_10_3 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \RTD.adc_state_i1_LC_3_10_3  (
            .in0(N__22337),
            .in1(N__22610),
            .in2(N__19650),
            .in3(N__22516),
            .lcout(\RTD.adc_state_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40538),
            .ce(N__19643),
            .sr(_gnd_net_));
    defparam \RTD.i27_4_lut_4_lut_LC_3_10_4 .C_ON=1'b0;
    defparam \RTD.i27_4_lut_4_lut_LC_3_10_4 .SEQ_MODE=4'b0000;
    defparam \RTD.i27_4_lut_4_lut_LC_3_10_4 .LUT_INIT=16'b1010101010000110;
    LogicCell40 \RTD.i27_4_lut_4_lut_LC_3_10_4  (
            .in0(N__22098),
            .in1(N__20673),
            .in2(N__22645),
            .in3(N__22332),
            .lcout(\RTD.n11860 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i19474_4_lut_4_lut_LC_3_10_5 .C_ON=1'b0;
    defparam \RTD.i19474_4_lut_4_lut_LC_3_10_5 .SEQ_MODE=4'b0000;
    defparam \RTD.i19474_4_lut_4_lut_LC_3_10_5 .LUT_INIT=16'b1011111111110111;
    LogicCell40 \RTD.i19474_4_lut_4_lut_LC_3_10_5  (
            .in0(N__22068),
            .in1(N__22609),
            .in2(N__22378),
            .in3(N__20687),
            .lcout(\RTD.n8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i31_4_lut_3_lut_LC_3_10_6 .C_ON=1'b0;
    defparam \RTD.i31_4_lut_3_lut_LC_3_10_6 .SEQ_MODE=4'b0000;
    defparam \RTD.i31_4_lut_3_lut_LC_3_10_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \RTD.i31_4_lut_3_lut_LC_3_10_6  (
            .in0(N__22603),
            .in1(N__22327),
            .in2(_gnd_net_),
            .in3(N__20672),
            .lcout(\RTD.n14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_2_lut_3_lut_4_lut_LC_3_10_7 .C_ON=1'b0;
    defparam \RTD.i1_2_lut_3_lut_4_lut_LC_3_10_7 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_2_lut_3_lut_4_lut_LC_3_10_7 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \RTD.i1_2_lut_3_lut_4_lut_LC_3_10_7  (
            .in0(N__22067),
            .in1(N__22604),
            .in2(N__22377),
            .in3(N__20686),
            .lcout(\RTD.n20370 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adress_i1_LC_5_7_0 .C_ON=1'b0;
    defparam \RTD.adress_i1_LC_5_7_0 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i1_LC_5_7_0 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \RTD.adress_i1_LC_5_7_0  (
            .in0(N__19733),
            .in1(N__19786),
            .in2(N__20409),
            .in3(N__20388),
            .lcout(adress_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40611),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adress_i2_LC_5_7_1 .C_ON=1'b0;
    defparam \RTD.adress_i2_LC_5_7_1 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i2_LC_5_7_1 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \RTD.adress_i2_LC_5_7_1  (
            .in0(N__20389),
            .in1(N__19718),
            .in2(N__19737),
            .in3(N__19795),
            .lcout(adress_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40611),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adress_i3_LC_5_7_2 .C_ON=1'b0;
    defparam \RTD.adress_i3_LC_5_7_2 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i3_LC_5_7_2 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \RTD.adress_i3_LC_5_7_2  (
            .in0(N__19706),
            .in1(N__19787),
            .in2(N__19722),
            .in3(N__20390),
            .lcout(adress_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40611),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adress_i4_LC_5_7_3 .C_ON=1'b0;
    defparam \RTD.adress_i4_LC_5_7_3 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i4_LC_5_7_3 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \RTD.adress_i4_LC_5_7_3  (
            .in0(N__20391),
            .in1(N__19694),
            .in2(N__19796),
            .in3(N__19707),
            .lcout(adress_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40611),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adress_i5_LC_5_7_4 .C_ON=1'b0;
    defparam \RTD.adress_i5_LC_5_7_4 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i5_LC_5_7_4 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \RTD.adress_i5_LC_5_7_4  (
            .in0(N__19838),
            .in1(N__19788),
            .in2(N__19698),
            .in3(N__20392),
            .lcout(adress_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40611),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adress_i6_LC_5_7_5 .C_ON=1'b0;
    defparam \RTD.adress_i6_LC_5_7_5 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i6_LC_5_7_5 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \RTD.adress_i6_LC_5_7_5  (
            .in0(N__20393),
            .in1(N__19839),
            .in2(N__19797),
            .in3(N__20516),
            .lcout(adress_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40611),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i0_LC_5_7_6 .C_ON=1'b0;
    defparam \RTD.read_buf_i0_LC_5_7_6 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i0_LC_5_7_6 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \RTD.read_buf_i0_LC_5_7_6  (
            .in0(N__21211),
            .in1(N__20968),
            .in2(N__19830),
            .in3(N__21045),
            .lcout(read_buf_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40611),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i11_LC_5_8_0 .C_ON=1'b0;
    defparam \RTD.read_buf_i11_LC_5_8_0 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i11_LC_5_8_0 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \RTD.read_buf_i11_LC_5_8_0  (
            .in0(N__19931),
            .in1(N__20950),
            .in2(N__20000),
            .in3(N__21042),
            .lcout(read_buf_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40609),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_2_lut_adj_8_LC_5_8_1 .C_ON=1'b0;
    defparam \RTD.i1_2_lut_adj_8_LC_5_8_1 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_2_lut_adj_8_LC_5_8_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \RTD.i1_2_lut_adj_8_LC_5_8_1  (
            .in0(_gnd_net_),
            .in1(N__20495),
            .in2(_gnd_net_),
            .in3(N__20427),
            .lcout(\RTD.n16766 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i14_LC_5_8_2 .C_ON=1'b0;
    defparam \RTD.read_buf_i14_LC_5_8_2 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i14_LC_5_8_2 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \RTD.read_buf_i14_LC_5_8_2  (
            .in0(N__21069),
            .in1(N__20951),
            .in2(N__19899),
            .in3(N__21043),
            .lcout(read_buf_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40609),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i19471_4_lut_4_lut_LC_5_8_3 .C_ON=1'b0;
    defparam \RTD.i19471_4_lut_4_lut_LC_5_8_3 .SEQ_MODE=4'b0000;
    defparam \RTD.i19471_4_lut_4_lut_LC_5_8_3 .LUT_INIT=16'b1110011000111100;
    LogicCell40 \RTD.i19471_4_lut_4_lut_LC_5_8_3  (
            .in0(N__22404),
            .in1(N__20748),
            .in2(N__22695),
            .in3(N__22188),
            .lcout(\RTD.n11915 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i10_LC_5_8_4 .C_ON=1'b0;
    defparam \RTD.read_buf_i10_LC_5_8_4 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i10_LC_5_8_4 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \RTD.read_buf_i10_LC_5_8_4  (
            .in0(N__19930),
            .in1(N__20949),
            .in2(N__20775),
            .in3(N__21041),
            .lcout(read_buf_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40609),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i12177_2_lut_LC_5_8_5 .C_ON=1'b0;
    defparam \RTD.i12177_2_lut_LC_5_8_5 .SEQ_MODE=4'b0000;
    defparam \RTD.i12177_2_lut_LC_5_8_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \RTD.i12177_2_lut_LC_5_8_5  (
            .in0(N__22687),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20744),
            .lcout(n14692),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_3_lut_4_lut_LC_5_8_6 .C_ON=1'b0;
    defparam \RTD.i1_3_lut_4_lut_LC_5_8_6 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_3_lut_4_lut_LC_5_8_6 .LUT_INIT=16'b1000101010010100;
    LogicCell40 \RTD.i1_3_lut_4_lut_LC_5_8_6  (
            .in0(N__22187),
            .in1(N__22691),
            .in2(N__20754),
            .in3(N__22405),
            .lcout(\RTD.n15280 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i6_LC_5_9_0 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i6_LC_5_9_0 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i6_LC_5_9_0 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \RTD.READ_DATA_i6_LC_5_9_0  (
            .in0(N__43472),
            .in1(N__21165),
            .in2(N__20880),
            .in3(N__22156),
            .lcout(buf_readRTD_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40610),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i10_LC_5_9_1 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i10_LC_5_9_1 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i10_LC_5_9_1 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \RTD.READ_DATA_i10_LC_5_9_1  (
            .in0(N__22153),
            .in1(N__19935),
            .in2(N__21173),
            .in3(N__23348),
            .lcout(buf_readRTD_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40610),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_4_lut_4_lut_LC_5_9_2 .C_ON=1'b0;
    defparam \RTD.i1_4_lut_4_lut_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_4_lut_4_lut_LC_5_9_2 .LUT_INIT=16'b1110010100000001;
    LogicCell40 \RTD.i1_4_lut_4_lut_LC_5_9_2  (
            .in0(N__20743),
            .in1(N__22375),
            .in2(N__22192),
            .in3(N__22670),
            .lcout(n13212),
            .ltout(n13212_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i15_LC_5_9_3 .C_ON=1'b0;
    defparam \RTD.read_buf_i15_LC_5_9_3 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i15_LC_5_9_3 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \RTD.read_buf_i15_LC_5_9_3  (
            .in0(N__19898),
            .in1(N__19910),
            .in2(N__19917),
            .in3(N__20921),
            .lcout(read_buf_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40610),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i15_LC_5_9_4 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i15_LC_5_9_4 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i15_LC_5_9_4 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \RTD.READ_DATA_i15_LC_5_9_4  (
            .in0(N__27149),
            .in1(N__21164),
            .in2(N__19914),
            .in3(N__22155),
            .lcout(buf_readRTD_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40610),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_4_lut_4_lut_adj_16_LC_5_9_5 .C_ON=1'b0;
    defparam \RTD.i1_4_lut_4_lut_adj_16_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_4_lut_4_lut_adj_16_LC_5_9_5 .LUT_INIT=16'b1110000010000000;
    LogicCell40 \RTD.i1_4_lut_4_lut_adj_16_LC_5_9_5  (
            .in0(N__22152),
            .in1(N__22376),
            .in2(N__22692),
            .in3(N__20742),
            .lcout(n11856),
            .ltout(n11856_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i14_LC_5_9_6 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i14_LC_5_9_6 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i14_LC_5_9_6 .LUT_INIT=16'b0011101000001010;
    LogicCell40 \RTD.READ_DATA_i14_LC_5_9_6  (
            .in0(N__22814),
            .in1(N__22154),
            .in2(N__19902),
            .in3(N__19897),
            .lcout(buf_readRTD_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40610),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.mode_53_LC_5_9_7 .C_ON=1'b0;
    defparam \RTD.mode_53_LC_5_9_7 .SEQ_MODE=4'b1000;
    defparam \RTD.mode_53_LC_5_9_7 .LUT_INIT=16'b1011101010101010;
    LogicCell40 \RTD.mode_53_LC_5_9_7  (
            .in0(N__19881),
            .in1(N__22527),
            .in2(N__22971),
            .in3(N__20430),
            .lcout(\RTD.mode ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40610),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i4_LC_5_10_0 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i4_LC_5_10_0 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i4_LC_5_10_0 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \RTD.READ_DATA_i4_LC_5_10_0  (
            .in0(N__22179),
            .in1(N__30620),
            .in2(N__20019),
            .in3(N__21161),
            .lcout(buf_readRTD_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40569),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i6_LC_5_10_1 .C_ON=1'b0;
    defparam \RTD.read_buf_i6_LC_5_10_1 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i6_LC_5_10_1 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \RTD.read_buf_i6_LC_5_10_1  (
            .in0(N__21029),
            .in1(N__19973),
            .in2(N__20975),
            .in3(N__20872),
            .lcout(read_buf_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40569),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i12_LC_5_10_2 .C_ON=1'b0;
    defparam \RTD.read_buf_i12_LC_5_10_2 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i12_LC_5_10_2 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \RTD.read_buf_i12_LC_5_10_2  (
            .in0(N__21082),
            .in1(N__20959),
            .in2(N__21044),
            .in3(N__19999),
            .lcout(read_buf_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40569),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i5_LC_5_10_3 .C_ON=1'b0;
    defparam \RTD.read_buf_i5_LC_5_10_3 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i5_LC_5_10_3 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \RTD.read_buf_i5_LC_5_10_3  (
            .in0(N__21028),
            .in1(N__19972),
            .in2(N__20974),
            .in3(N__20017),
            .lcout(read_buf_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40569),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i4_LC_5_10_4 .C_ON=1'b0;
    defparam \RTD.read_buf_i4_LC_5_10_4 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i4_LC_5_10_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \RTD.read_buf_i4_LC_5_10_4  (
            .in0(N__19954),
            .in1(N__20961),
            .in2(N__20018),
            .in3(N__21031),
            .lcout(read_buf_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40569),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i12_LC_5_10_5 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i12_LC_5_10_5 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i12_LC_5_10_5 .LUT_INIT=16'b0010111000100010;
    LogicCell40 \RTD.READ_DATA_i12_LC_5_10_5  (
            .in0(N__35021),
            .in1(N__21155),
            .in2(N__22215),
            .in3(N__21083),
            .lcout(buf_readRTD_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40569),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i3_LC_5_10_6 .C_ON=1'b0;
    defparam \RTD.read_buf_i3_LC_5_10_6 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i3_LC_5_10_6 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \RTD.read_buf_i3_LC_5_10_6  (
            .in0(N__21198),
            .in1(N__20960),
            .in2(N__19958),
            .in3(N__21030),
            .lcout(read_buf_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40569),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i11_LC_5_10_7 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i11_LC_5_10_7 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i11_LC_5_10_7 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \RTD.READ_DATA_i11_LC_5_10_7  (
            .in0(N__25907),
            .in1(N__21154),
            .in2(N__20001),
            .in3(N__22180),
            .lcout(buf_readRTD_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40569),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i5_LC_5_11_2 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i5_LC_5_11_2 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i5_LC_5_11_2 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \RTD.READ_DATA_i5_LC_5_11_2  (
            .in0(N__22181),
            .in1(N__19977),
            .in2(N__21174),
            .in3(N__28283),
            .lcout(buf_readRTD_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40612),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i3_LC_5_11_3 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i3_LC_5_11_3 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i3_LC_5_11_3 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \RTD.READ_DATA_i3_LC_5_11_3  (
            .in0(N__40805),
            .in1(N__21169),
            .in2(N__19959),
            .in3(N__22182),
            .lcout(buf_readRTD_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40612),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_6_i19_3_lut_LC_5_11_4.C_ON=1'b0;
    defparam mux_130_Mux_6_i19_3_lut_LC_5_11_4.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_6_i19_3_lut_LC_5_11_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_130_Mux_6_i19_3_lut_LC_5_11_4 (
            .in0(N__25404),
            .in1(N__23138),
            .in2(_gnd_net_),
            .in3(N__57151),
            .lcout(),
            .ltout(n19_adj_1600_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_6_i22_3_lut_LC_5_11_5.C_ON=1'b0;
    defparam mux_130_Mux_6_i22_3_lut_LC_5_11_5.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_6_i22_3_lut_LC_5_11_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 mux_130_Mux_6_i22_3_lut_LC_5_11_5 (
            .in0(_gnd_net_),
            .in1(N__20830),
            .in2(N__19938),
            .in3(N__47515),
            .lcout(n22_adj_1601),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i0_LC_5_12_0 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i0_LC_5_12_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i0_LC_5_12_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i0_LC_5_12_0  (
            .in0(N__27974),
            .in1(N__27804),
            .in2(N__21377),
            .in3(N__27259),
            .lcout(buf_adcdata_vac_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56059),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_7_i19_3_lut_LC_5_12_1.C_ON=1'b0;
    defparam mux_130_Mux_7_i19_3_lut_LC_5_12_1.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_7_i19_3_lut_LC_5_12_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_130_Mux_7_i19_3_lut_LC_5_12_1 (
            .in0(N__26766),
            .in1(N__20032),
            .in2(_gnd_net_),
            .in3(N__57260),
            .lcout(),
            .ltout(n19_adj_1597_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_7_i22_3_lut_LC_5_12_2.C_ON=1'b0;
    defparam mux_130_Mux_7_i22_3_lut_LC_5_12_2.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_7_i22_3_lut_LC_5_12_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 mux_130_Mux_7_i22_3_lut_LC_5_12_2 (
            .in0(_gnd_net_),
            .in1(N__21394),
            .in2(N__20043),
            .in3(N__47694),
            .lcout(n22_adj_1598),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i7_LC_5_12_3 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i7_LC_5_12_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i7_LC_5_12_3 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i7_LC_5_12_3  (
            .in0(N__27802),
            .in1(N__27977),
            .in2(N__23037),
            .in3(N__20033),
            .lcout(buf_adcdata_vac_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56059),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i4_LC_5_12_4 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i4_LC_5_12_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i4_LC_5_12_4 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC.ADC_DATA_i4_LC_5_12_4  (
            .in0(N__27976),
            .in1(N__27805),
            .in2(N__21287),
            .in3(N__21330),
            .lcout(buf_adcdata_vac_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56059),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i11_LC_5_12_5 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i11_LC_5_12_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i11_LC_5_12_5 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i11_LC_5_12_5  (
            .in0(N__27803),
            .in1(N__23284),
            .in2(N__22799),
            .in3(N__28244),
            .lcout(cmd_rdadctmp_11_adj_1481),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56059),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i13_LC_5_12_6 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i13_LC_5_12_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i13_LC_5_12_6 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i13_LC_5_12_6  (
            .in0(N__28245),
            .in1(N__21329),
            .in2(N__23227),
            .in3(N__27806),
            .lcout(cmd_rdadctmp_13_adj_1479),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56059),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i23_LC_5_12_7 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i23_LC_5_12_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i23_LC_5_12_7 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i23_LC_5_12_7  (
            .in0(N__27801),
            .in1(N__27975),
            .in2(N__21240),
            .in3(N__27100),
            .lcout(buf_adcdata_vac_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56059),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i3_LC_5_13_0 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i3_LC_5_13_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i3_LC_5_13_0 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i3_LC_5_13_0  (
            .in0(N__28213),
            .in1(N__20064),
            .in2(N__27758),
            .in3(N__21416),
            .lcout(cmd_rdadctmp_3_adj_1489),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56073),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i1_4_lut_LC_5_13_1 .C_ON=1'b0;
    defparam \ADC_VAC.i1_4_lut_LC_5_13_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i1_4_lut_LC_5_13_1 .LUT_INIT=16'b0000000100100010;
    LogicCell40 \ADC_VAC.i1_4_lut_LC_5_13_1  (
            .in0(N__21620),
            .in1(N__27655),
            .in2(N__21722),
            .in3(N__21556),
            .lcout(\ADC_VAC.n12803 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i8_LC_5_13_2 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i8_LC_5_13_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i8_LC_5_13_2 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i8_LC_5_13_2  (
            .in0(N__28215),
            .in1(N__20112),
            .in2(N__27759),
            .in3(N__21367),
            .lcout(cmd_rdadctmp_8_adj_1484),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56073),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i7_LC_5_13_3 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i7_LC_5_13_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i7_LC_5_13_3 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i7_LC_5_13_3  (
            .in0(N__20111),
            .in1(N__27658),
            .in2(N__24690),
            .in3(N__28214),
            .lcout(cmd_rdadctmp_7_adj_1485),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56073),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i0_LC_5_13_5 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i0_LC_5_13_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i0_LC_5_13_5 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i0_LC_5_13_5  (
            .in0(N__20084),
            .in1(N__27656),
            .in2(N__20103),
            .in3(N__28210),
            .lcout(cmd_rdadctmp_0_adj_1492),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56073),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i1_LC_5_13_6 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i1_LC_5_13_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i1_LC_5_13_6 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i1_LC_5_13_6  (
            .in0(N__28211),
            .in1(N__20072),
            .in2(N__27757),
            .in3(N__20085),
            .lcout(cmd_rdadctmp_1_adj_1491),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56073),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i2_LC_5_13_7 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i2_LC_5_13_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i2_LC_5_13_7 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i2_LC_5_13_7  (
            .in0(N__20063),
            .in1(N__27657),
            .in2(N__20076),
            .in3(N__28212),
            .lcout(cmd_rdadctmp_2_adj_1490),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56073),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.bit_cnt_i0_LC_5_14_0 .C_ON=1'b1;
    defparam \ADC_VAC.bit_cnt_i0_LC_5_14_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i0_LC_5_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i0_LC_5_14_0  (
            .in0(_gnd_net_),
            .in1(N__20184),
            .in2(_gnd_net_),
            .in3(N__20055),
            .lcout(\ADC_VAC.bit_cnt_0 ),
            .ltout(),
            .carryin(bfn_5_14_0_),
            .carryout(\ADC_VAC.n19835 ),
            .clk(N__56083),
            .ce(N__20142),
            .sr(N__20124));
    defparam \ADC_VAC.bit_cnt_i1_LC_5_14_1 .C_ON=1'b1;
    defparam \ADC_VAC.bit_cnt_i1_LC_5_14_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i1_LC_5_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i1_LC_5_14_1  (
            .in0(_gnd_net_),
            .in1(N__20225),
            .in2(_gnd_net_),
            .in3(N__20052),
            .lcout(\ADC_VAC.bit_cnt_1 ),
            .ltout(),
            .carryin(\ADC_VAC.n19835 ),
            .carryout(\ADC_VAC.n19836 ),
            .clk(N__56083),
            .ce(N__20142),
            .sr(N__20124));
    defparam \ADC_VAC.bit_cnt_i2_LC_5_14_2 .C_ON=1'b1;
    defparam \ADC_VAC.bit_cnt_i2_LC_5_14_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i2_LC_5_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i2_LC_5_14_2  (
            .in0(_gnd_net_),
            .in1(N__20211),
            .in2(_gnd_net_),
            .in3(N__20049),
            .lcout(\ADC_VAC.bit_cnt_2 ),
            .ltout(),
            .carryin(\ADC_VAC.n19836 ),
            .carryout(\ADC_VAC.n19837 ),
            .clk(N__56083),
            .ce(N__20142),
            .sr(N__20124));
    defparam \ADC_VAC.bit_cnt_i3_LC_5_14_3 .C_ON=1'b1;
    defparam \ADC_VAC.bit_cnt_i3_LC_5_14_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i3_LC_5_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i3_LC_5_14_3  (
            .in0(_gnd_net_),
            .in1(N__20238),
            .in2(_gnd_net_),
            .in3(N__20046),
            .lcout(\ADC_VAC.bit_cnt_3 ),
            .ltout(),
            .carryin(\ADC_VAC.n19837 ),
            .carryout(\ADC_VAC.n19838 ),
            .clk(N__56083),
            .ce(N__20142),
            .sr(N__20124));
    defparam \ADC_VAC.bit_cnt_i4_LC_5_14_4 .C_ON=1'b1;
    defparam \ADC_VAC.bit_cnt_i4_LC_5_14_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i4_LC_5_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i4_LC_5_14_4  (
            .in0(_gnd_net_),
            .in1(N__20250),
            .in2(_gnd_net_),
            .in3(N__20262),
            .lcout(\ADC_VAC.bit_cnt_4 ),
            .ltout(),
            .carryin(\ADC_VAC.n19838 ),
            .carryout(\ADC_VAC.n19839 ),
            .clk(N__56083),
            .ce(N__20142),
            .sr(N__20124));
    defparam \ADC_VAC.bit_cnt_i5_LC_5_14_5 .C_ON=1'b1;
    defparam \ADC_VAC.bit_cnt_i5_LC_5_14_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i5_LC_5_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i5_LC_5_14_5  (
            .in0(_gnd_net_),
            .in1(N__20157),
            .in2(_gnd_net_),
            .in3(N__20259),
            .lcout(\ADC_VAC.bit_cnt_5 ),
            .ltout(),
            .carryin(\ADC_VAC.n19839 ),
            .carryout(\ADC_VAC.n19840 ),
            .clk(N__56083),
            .ce(N__20142),
            .sr(N__20124));
    defparam \ADC_VAC.bit_cnt_i6_LC_5_14_6 .C_ON=1'b1;
    defparam \ADC_VAC.bit_cnt_i6_LC_5_14_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i6_LC_5_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i6_LC_5_14_6  (
            .in0(_gnd_net_),
            .in1(N__20198),
            .in2(_gnd_net_),
            .in3(N__20256),
            .lcout(\ADC_VAC.bit_cnt_6 ),
            .ltout(),
            .carryin(\ADC_VAC.n19840 ),
            .carryout(\ADC_VAC.n19841 ),
            .clk(N__56083),
            .ce(N__20142),
            .sr(N__20124));
    defparam \ADC_VAC.bit_cnt_i7_LC_5_14_7 .C_ON=1'b0;
    defparam \ADC_VAC.bit_cnt_i7_LC_5_14_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.bit_cnt_i7_LC_5_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VAC.bit_cnt_i7_LC_5_14_7  (
            .in0(_gnd_net_),
            .in1(N__20169),
            .in2(_gnd_net_),
            .in3(N__20253),
            .lcout(\ADC_VAC.bit_cnt_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56083),
            .ce(N__20142),
            .sr(N__20124));
    defparam \ADC_VAC.i18497_4_lut_LC_5_15_0 .C_ON=1'b0;
    defparam \ADC_VAC.i18497_4_lut_LC_5_15_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i18497_4_lut_LC_5_15_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VAC.i18497_4_lut_LC_5_15_0  (
            .in0(N__20249),
            .in1(N__20237),
            .in2(N__20226),
            .in3(N__20210),
            .lcout(),
            .ltout(\ADC_VAC.n21224_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i18507_4_lut_LC_5_15_1 .C_ON=1'b0;
    defparam \ADC_VAC.i18507_4_lut_LC_5_15_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i18507_4_lut_LC_5_15_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VAC.i18507_4_lut_LC_5_15_1  (
            .in0(N__20199),
            .in1(N__20183),
            .in2(N__20172),
            .in3(N__20168),
            .lcout(),
            .ltout(\ADC_VAC.n21234_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i19109_4_lut_LC_5_15_2 .C_ON=1'b0;
    defparam \ADC_VAC.i19109_4_lut_LC_5_15_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i19109_4_lut_LC_5_15_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \ADC_VAC.i19109_4_lut_LC_5_15_2  (
            .in0(N__27670),
            .in1(N__20156),
            .in2(N__20145),
            .in3(N__21552),
            .lcout(\ADC_VAC.n21468 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i12536_2_lut_LC_5_15_3 .C_ON=1'b0;
    defparam \ADC_VAC.i12536_2_lut_LC_5_15_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i12536_2_lut_LC_5_15_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \ADC_VAC.i12536_2_lut_LC_5_15_3  (
            .in0(N__21617),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20138),
            .lcout(\ADC_VAC.n15052 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i1_4_lut_adj_36_LC_5_15_4 .C_ON=1'b0;
    defparam \ADC_VAC.i1_4_lut_adj_36_LC_5_15_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i1_4_lut_adj_36_LC_5_15_4 .LUT_INIT=16'b1010101111101111;
    LogicCell40 \ADC_VAC.i1_4_lut_adj_36_LC_5_15_4  (
            .in0(N__27668),
            .in1(N__21616),
            .in2(N__21723),
            .in3(N__28713),
            .lcout(),
            .ltout(\ADC_VAC.n21157_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i1_2_lut_adj_37_LC_5_15_5 .C_ON=1'b0;
    defparam \ADC_VAC.i1_2_lut_adj_37_LC_5_15_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i1_2_lut_adj_37_LC_5_15_5 .LUT_INIT=16'b1111010111110101;
    LogicCell40 \ADC_VAC.i1_2_lut_adj_37_LC_5_15_5  (
            .in0(N__21553),
            .in1(_gnd_net_),
            .in2(N__20367),
            .in3(_gnd_net_),
            .lcout(\ADC_VAC.n21158 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i19419_2_lut_LC_5_15_7 .C_ON=1'b0;
    defparam \ADC_VAC.i19419_2_lut_LC_5_15_7 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i19419_2_lut_LC_5_15_7 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \ADC_VAC.i19419_2_lut_LC_5_15_7  (
            .in0(_gnd_net_),
            .in1(N__27669),
            .in2(_gnd_net_),
            .in3(N__21474),
            .lcout(\ADC_VAC.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.adc_state_i0_LC_5_16_0 .C_ON=1'b0;
    defparam \ADC_VAC.adc_state_i0_LC_5_16_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.adc_state_i0_LC_5_16_0 .LUT_INIT=16'b0101011100000010;
    LogicCell40 \ADC_VAC.adc_state_i0_LC_5_16_0  (
            .in0(N__21618),
            .in1(N__21555),
            .in2(N__27756),
            .in3(N__20364),
            .lcout(adc_state_0_adj_1460),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56095),
            .ce(N__20358),
            .sr(_gnd_net_));
    defparam \CLK_DDS.dds_state_i1_LC_6_6_0 .C_ON=1'b0;
    defparam \CLK_DDS.dds_state_i1_LC_6_6_0 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.dds_state_i1_LC_6_6_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \CLK_DDS.dds_state_i1_LC_6_6_0  (
            .in0(_gnd_net_),
            .in1(N__30103),
            .in2(_gnd_net_),
            .in3(N__29941),
            .lcout(dds_state_1_adj_1495),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55955),
            .ce(N__29711),
            .sr(N__29844));
    defparam \RTD.CS_52_LC_6_7_0 .C_ON=1'b0;
    defparam \RTD.CS_52_LC_6_7_0 .SEQ_MODE=4'b1000;
    defparam \RTD.CS_52_LC_6_7_0 .LUT_INIT=16'b0001000101011111;
    LogicCell40 \RTD.CS_52_LC_6_7_0  (
            .in0(N__22399),
            .in1(N__20729),
            .in2(N__20346),
            .in3(N__22685),
            .lcout(RTD_CS),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40614),
            .ce(N__20625),
            .sr(_gnd_net_));
    defparam \RTD.i18454_2_lut_LC_6_7_2 .C_ON=1'b0;
    defparam \RTD.i18454_2_lut_LC_6_7_2 .SEQ_MODE=4'b0000;
    defparam \RTD.i18454_2_lut_LC_6_7_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \RTD.i18454_2_lut_LC_6_7_2  (
            .in0(_gnd_net_),
            .in1(N__22683),
            .in2(_gnd_net_),
            .in3(N__20726),
            .lcout(),
            .ltout(\RTD.n21181_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i30_4_lut_LC_6_7_3 .C_ON=1'b0;
    defparam \RTD.i30_4_lut_LC_6_7_3 .SEQ_MODE=4'b0000;
    defparam \RTD.i30_4_lut_LC_6_7_3 .LUT_INIT=16'b1000101110001000;
    LogicCell40 \RTD.i30_4_lut_LC_6_7_3  (
            .in0(N__20298),
            .in1(N__22186),
            .in2(N__20286),
            .in3(N__22706),
            .lcout(\RTD.n13137 ),
            .ltout(\RTD.n13137_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i12599_2_lut_LC_6_7_4 .C_ON=1'b0;
    defparam \RTD.i12599_2_lut_LC_6_7_4 .SEQ_MODE=4'b0000;
    defparam \RTD.i12599_2_lut_LC_6_7_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \RTD.i12599_2_lut_LC_6_7_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20283),
            .in3(N__22684),
            .lcout(\RTD.n15115 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_2_lut_adj_9_LC_6_7_5 .C_ON=1'b0;
    defparam \RTD.i1_2_lut_adj_9_LC_6_7_5 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_2_lut_adj_9_LC_6_7_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \RTD.i1_2_lut_adj_9_LC_6_7_5  (
            .in0(N__20728),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22398),
            .lcout(\RTD.n7889 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_2_lut_3_lut_adj_22_LC_6_7_7 .C_ON=1'b0;
    defparam \RTD.i1_2_lut_3_lut_adj_22_LC_6_7_7 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_2_lut_3_lut_adj_22_LC_6_7_7 .LUT_INIT=16'b1101110111111111;
    LogicCell40 \RTD.i1_2_lut_3_lut_adj_22_LC_6_7_7  (
            .in0(N__20727),
            .in1(N__20589),
            .in2(_gnd_net_),
            .in3(N__20559),
            .lcout(\RTD.n19026 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adress_i7_LC_6_8_0 .C_ON=1'b0;
    defparam \RTD.adress_i7_LC_6_8_0 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i7_LC_6_8_0 .LUT_INIT=16'b1110001011000000;
    LogicCell40 \RTD.adress_i7_LC_6_8_0  (
            .in0(N__22403),
            .in1(N__20753),
            .in2(N__20517),
            .in3(N__20429),
            .lcout(\RTD.adress_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40608),
            .ce(N__20397),
            .sr(N__20814));
    defparam \RTD.i1_4_lut_LC_6_8_1 .C_ON=1'b0;
    defparam \RTD.i1_4_lut_LC_6_8_1 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_4_lut_LC_6_8_1 .LUT_INIT=16'b0111110110111110;
    LogicCell40 \RTD.i1_4_lut_LC_6_8_1  (
            .in0(N__25739),
            .in1(N__20786),
            .in2(N__27078),
            .in3(N__22902),
            .lcout(),
            .ltout(\RTD.n9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i7_4_lut_LC_6_8_2 .C_ON=1'b0;
    defparam \RTD.i7_4_lut_LC_6_8_2 .SEQ_MODE=4'b0000;
    defparam \RTD.i7_4_lut_LC_6_8_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \RTD.i7_4_lut_LC_6_8_2  (
            .in0(N__22476),
            .in1(N__22713),
            .in2(N__20502),
            .in3(N__22746),
            .lcout(\RTD.adress_7_N_1086_7 ),
            .ltout(\RTD.adress_7_N_1086_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i1_2_lut_adj_6_LC_6_8_3 .C_ON=1'b0;
    defparam \RTD.i1_2_lut_adj_6_LC_6_8_3 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_2_lut_adj_6_LC_6_8_3 .LUT_INIT=16'b1111000011111111;
    LogicCell40 \RTD.i1_2_lut_adj_6_LC_6_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20499),
            .in3(N__22400),
            .lcout(\RTD.n11 ),
            .ltout(\RTD.n11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i34_4_lut_LC_6_8_4 .C_ON=1'b0;
    defparam \RTD.i34_4_lut_LC_6_8_4 .SEQ_MODE=4'b0000;
    defparam \RTD.i34_4_lut_LC_6_8_4 .LUT_INIT=16'b1010101011110011;
    LogicCell40 \RTD.i34_4_lut_LC_6_8_4  (
            .in0(N__22401),
            .in1(N__20496),
            .in2(N__20460),
            .in3(N__20751),
            .lcout(),
            .ltout(\RTD.n19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i35_4_lut_LC_6_8_5 .C_ON=1'b0;
    defparam \RTD.i35_4_lut_LC_6_8_5 .SEQ_MODE=4'b0000;
    defparam \RTD.i35_4_lut_LC_6_8_5 .LUT_INIT=16'b1000100010111000;
    LogicCell40 \RTD.i35_4_lut_LC_6_8_5  (
            .in0(N__22544),
            .in1(N__22686),
            .in2(N__20457),
            .in3(N__22216),
            .lcout(n13054),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.adress_i0_LC_6_8_6 .C_ON=1'b0;
    defparam \RTD.adress_i0_LC_6_8_6 .SEQ_MODE=4'b1000;
    defparam \RTD.adress_i0_LC_6_8_6 .LUT_INIT=16'b1101000111110011;
    LogicCell40 \RTD.adress_i0_LC_6_8_6  (
            .in0(N__22402),
            .in1(N__20752),
            .in2(N__20450),
            .in3(N__20428),
            .lcout(adress_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40608),
            .ce(N__20397),
            .sr(N__20814));
    defparam \RTD.i1_2_lut_3_lut_LC_6_9_0 .C_ON=1'b0;
    defparam \RTD.i1_2_lut_3_lut_LC_6_9_0 .SEQ_MODE=4'b0000;
    defparam \RTD.i1_2_lut_3_lut_LC_6_9_0 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \RTD.i1_2_lut_3_lut_LC_6_9_0  (
            .in0(N__22352),
            .in1(N__20749),
            .in2(_gnd_net_),
            .in3(N__22175),
            .lcout(\RTD.n21036 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i8_LC_6_9_1 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i8_LC_6_9_1 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i8_LC_6_9_1 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \RTD.READ_DATA_i8_LC_6_9_1  (
            .in0(N__22177),
            .in1(N__25817),
            .in2(N__20609),
            .in3(N__21163),
            .lcout(buf_readRTD_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40613),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i9_LC_6_9_2 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i9_LC_6_9_2 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i9_LC_6_9_2 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \RTD.READ_DATA_i9_LC_6_9_2  (
            .in0(N__21162),
            .in1(N__22886),
            .in2(N__20774),
            .in3(N__22178),
            .lcout(buf_readRTD_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40613),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i6_LC_6_9_3 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i6_LC_6_9_3 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i6_LC_6_9_3 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \RTD.cfg_buf_i6_LC_6_9_3  (
            .in0(N__22960),
            .in1(N__23008),
            .in2(N__27070),
            .in3(N__20787),
            .lcout(\RTD.cfg_buf_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40613),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i1_LC_6_9_4 .C_ON=1'b0;
    defparam \RTD.read_buf_i1_LC_6_9_4 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i1_LC_6_9_4 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \RTD.read_buf_i1_LC_6_9_4  (
            .in0(N__21038),
            .in1(N__21218),
            .in2(N__21102),
            .in3(N__20922),
            .lcout(read_buf_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40613),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i9_LC_6_9_5 .C_ON=1'b0;
    defparam \RTD.read_buf_i9_LC_6_9_5 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i9_LC_6_9_5 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \RTD.read_buf_i9_LC_6_9_5  (
            .in0(N__20924),
            .in1(N__20767),
            .in2(N__20610),
            .in3(N__21040),
            .lcout(read_buf_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40613),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i19396_3_lut_3_lut_LC_6_9_6 .C_ON=1'b0;
    defparam \RTD.i19396_3_lut_3_lut_LC_6_9_6 .SEQ_MODE=4'b0000;
    defparam \RTD.i19396_3_lut_3_lut_LC_6_9_6 .LUT_INIT=16'b1010101000010001;
    LogicCell40 \RTD.i19396_3_lut_3_lut_LC_6_9_6  (
            .in0(N__22679),
            .in1(N__20750),
            .in2(_gnd_net_),
            .in3(N__22176),
            .lcout(\RTD.n11829 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i8_LC_6_9_7 .C_ON=1'b0;
    defparam \RTD.read_buf_i8_LC_6_9_7 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i8_LC_6_9_7 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \RTD.read_buf_i8_LC_6_9_7  (
            .in0(N__20923),
            .in1(N__20856),
            .in2(N__20608),
            .in3(N__21039),
            .lcout(read_buf_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40613),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i13_LC_6_10_0 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i13_LC_6_10_0 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i13_LC_6_10_0 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \RTD.READ_DATA_i13_LC_6_10_0  (
            .in0(N__22193),
            .in1(N__34892),
            .in2(N__21068),
            .in3(N__21152),
            .lcout(buf_readRTD_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40582),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i7_LC_6_10_1 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i7_LC_6_10_1 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i7_LC_6_10_1 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \RTD.READ_DATA_i7_LC_6_10_1  (
            .in0(N__21151),
            .in1(N__22196),
            .in2(N__23723),
            .in3(N__20855),
            .lcout(buf_readRTD_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40582),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i2_LC_6_10_2 .C_ON=1'b0;
    defparam \RTD.read_buf_i2_LC_6_10_2 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i2_LC_6_10_2 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \RTD.read_buf_i2_LC_6_10_2  (
            .in0(N__21101),
            .in1(N__20970),
            .in2(N__21196),
            .in3(N__21027),
            .lcout(read_buf_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40582),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i0_LC_6_10_3 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i0_LC_6_10_3 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i0_LC_6_10_3 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \RTD.READ_DATA_i0_LC_6_10_3  (
            .in0(N__21149),
            .in1(N__43697),
            .in2(N__21225),
            .in3(N__22197),
            .lcout(buf_readRTD_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40582),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i2_LC_6_10_4 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i2_LC_6_10_4 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i2_LC_6_10_4 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \RTD.READ_DATA_i2_LC_6_10_4  (
            .in0(N__22194),
            .in1(N__35159),
            .in2(N__21197),
            .in3(N__21153),
            .lcout(buf_readRTD_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40582),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.READ_DATA_i1_LC_6_10_5 .C_ON=1'b0;
    defparam \RTD.READ_DATA_i1_LC_6_10_5 .SEQ_MODE=4'b1000;
    defparam \RTD.READ_DATA_i1_LC_6_10_5 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \RTD.READ_DATA_i1_LC_6_10_5  (
            .in0(N__21150),
            .in1(N__22195),
            .in2(N__28337),
            .in3(N__21100),
            .lcout(buf_readRTD_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40582),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i13_LC_6_10_6 .C_ON=1'b0;
    defparam \RTD.read_buf_i13_LC_6_10_6 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i13_LC_6_10_6 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \RTD.read_buf_i13_LC_6_10_6  (
            .in0(N__21084),
            .in1(N__20969),
            .in2(N__21067),
            .in3(N__21026),
            .lcout(read_buf_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40582),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.read_buf_i7_LC_6_10_7 .C_ON=1'b0;
    defparam \RTD.read_buf_i7_LC_6_10_7 .SEQ_MODE=4'b1000;
    defparam \RTD.read_buf_i7_LC_6_10_7 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \RTD.read_buf_i7_LC_6_10_7  (
            .in0(N__21025),
            .in1(N__20854),
            .in2(N__20976),
            .in3(N__20876),
            .lcout(read_buf_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40582),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i0_LC_6_11_0 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i0_LC_6_11_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i0_LC_6_11_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i0_LC_6_11_0  (
            .in0(N__38590),
            .in1(N__38751),
            .in2(N__23496),
            .in3(N__27223),
            .lcout(buf_adcdata_iac_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56016),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i11_LC_6_11_2 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i11_LC_6_11_2 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i11_LC_6_11_2 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i11_LC_6_11_2  (
            .in0(N__38592),
            .in1(N__23527),
            .in2(N__24326),
            .in3(N__29392),
            .lcout(cmd_rdadctmp_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56016),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i6_LC_6_11_4 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i6_LC_6_11_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i6_LC_6_11_4 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i6_LC_6_11_4  (
            .in0(N__38591),
            .in1(N__38753),
            .in2(N__21497),
            .in3(N__20834),
            .lcout(buf_adcdata_iac_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56016),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i3_LC_6_11_5 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i3_LC_6_11_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i3_LC_6_11_5 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i3_LC_6_11_5  (
            .in0(N__38752),
            .in1(N__38594),
            .in2(N__23534),
            .in3(N__22846),
            .lcout(buf_adcdata_iac_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56016),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i14_LC_6_11_6 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i14_LC_6_11_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i14_LC_6_11_6 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i14_LC_6_11_6  (
            .in0(N__38593),
            .in1(N__24353),
            .in2(N__21496),
            .in3(N__29393),
            .lcout(cmd_rdadctmp_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56016),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i22_LC_6_11_7 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i22_LC_6_11_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i22_LC_6_11_7 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC.ADC_DATA_i22_LC_6_11_7  (
            .in0(N__27973),
            .in1(N__27800),
            .in2(N__23099),
            .in3(N__23202),
            .lcout(buf_adcdata_vac_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56016),
            .ce(),
            .sr(_gnd_net_));
    defparam i19316_2_lut_LC_6_12_0.C_ON=1'b0;
    defparam i19316_2_lut_LC_6_12_0.SEQ_MODE=4'b0000;
    defparam i19316_2_lut_LC_6_12_0.LUT_INIT=16'b0101010100000000;
    LogicCell40 i19316_2_lut_LC_6_12_0 (
            .in0(N__57187),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31974),
            .lcout(n21705),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_4_i19_3_lut_LC_6_12_2.C_ON=1'b0;
    defparam mux_130_Mux_4_i19_3_lut_LC_6_12_2.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_4_i19_3_lut_LC_6_12_2.LUT_INIT=16'b1010111110100000;
    LogicCell40 mux_130_Mux_4_i19_3_lut_LC_6_12_2 (
            .in0(N__25608),
            .in1(_gnd_net_),
            .in2(N__57259),
            .in3(N__21277),
            .lcout(),
            .ltout(n19_adj_1606_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_4_i22_3_lut_LC_6_12_3.C_ON=1'b0;
    defparam mux_130_Mux_4_i22_3_lut_LC_6_12_3.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_4_i22_3_lut_LC_6_12_3.LUT_INIT=16'b1111000010101010;
    LogicCell40 mux_130_Mux_4_i22_3_lut_LC_6_12_3 (
            .in0(N__21307),
            .in1(_gnd_net_),
            .in2(N__21261),
            .in3(N__47695),
            .lcout(),
            .ltout(n22_adj_1607_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_4_i30_3_lut_LC_6_12_4.C_ON=1'b0;
    defparam mux_130_Mux_4_i30_3_lut_LC_6_12_4.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_4_i30_3_lut_LC_6_12_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 mux_130_Mux_4_i30_3_lut_LC_6_12_4 (
            .in0(_gnd_net_),
            .in1(N__21258),
            .in2(N__21243),
            .in3(N__47091),
            .lcout(n30_adj_1608),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i31_LC_6_12_5 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i31_LC_6_12_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i31_LC_6_12_5 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i31_LC_6_12_5  (
            .in0(N__28191),
            .in1(N__23201),
            .in2(N__27847),
            .in3(N__21236),
            .lcout(cmd_rdadctmp_31_adj_1461),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56030),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i14_LC_6_12_6 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i14_LC_6_12_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i14_LC_6_12_6 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i14_LC_6_12_6  (
            .in0(N__23053),
            .in1(N__27796),
            .in2(N__23228),
            .in3(N__28190),
            .lcout(cmd_rdadctmp_14_adj_1478),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56030),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i7_LC_6_12_7 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i7_LC_6_12_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i7_LC_6_12_7 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i7_LC_6_12_7  (
            .in0(N__38764),
            .in1(N__38598),
            .in2(N__26301),
            .in3(N__21398),
            .lcout(buf_adcdata_iac_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56030),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i10_LC_6_13_0 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i10_LC_6_13_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i10_LC_6_13_0 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i10_LC_6_13_0  (
            .in0(N__22792),
            .in1(N__27723),
            .in2(N__23423),
            .in3(N__28187),
            .lcout(cmd_rdadctmp_10_adj_1482),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56046),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i9_LC_6_13_1 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i9_LC_6_13_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i9_LC_6_13_1 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i9_LC_6_13_1  (
            .in0(N__29383),
            .in1(N__36331),
            .in2(N__23489),
            .in3(N__38562),
            .lcout(cmd_rdadctmp_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56046),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i9_LC_6_13_2 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i9_LC_6_13_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i9_LC_6_13_2 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i9_LC_6_13_2  (
            .in0(N__23416),
            .in1(N__27725),
            .in2(N__21378),
            .in3(N__28189),
            .lcout(cmd_rdadctmp_9_adj_1483),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56046),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_7_i30_3_lut_LC_6_13_3.C_ON=1'b0;
    defparam mux_130_Mux_7_i30_3_lut_LC_6_13_3.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_7_i30_3_lut_LC_6_13_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_130_Mux_7_i30_3_lut_LC_6_13_3 (
            .in0(N__21351),
            .in1(N__21336),
            .in2(_gnd_net_),
            .in3(N__47048),
            .lcout(n30_adj_1599),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i12_LC_6_13_4 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i12_LC_6_13_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i12_LC_6_13_4 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i12_LC_6_13_4  (
            .in0(N__21328),
            .in1(N__27724),
            .in2(N__23297),
            .in3(N__28188),
            .lcout(cmd_rdadctmp_12_adj_1480),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56046),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i13_LC_6_13_6 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i13_LC_6_13_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i13_LC_6_13_6 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i13_LC_6_13_6  (
            .in0(N__38560),
            .in1(N__24346),
            .in2(N__23514),
            .in3(N__29384),
            .lcout(cmd_rdadctmp_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56046),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i4_LC_6_13_7 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i4_LC_6_13_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i4_LC_6_13_7 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_IAC.ADC_DATA_i4_LC_6_13_7  (
            .in0(N__38763),
            .in1(N__38561),
            .in2(N__21314),
            .in3(N__23513),
            .lcout(buf_adcdata_iac_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56046),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i4_LC_6_14_0.C_ON=1'b0;
    defparam buf_dds1_i4_LC_6_14_0.SEQ_MODE=4'b1000;
    defparam buf_dds1_i4_LC_6_14_0.LUT_INIT=16'b1110001000000000;
    LogicCell40 buf_dds1_i4_LC_6_14_0 (
            .in0(N__29452),
            .in1(N__46909),
            .in2(N__42714),
            .in3(N__46733),
            .lcout(buf_dds1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56060),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i3_LC_6_14_1.C_ON=1'b0;
    defparam comm_cmd_i3_LC_6_14_1.SEQ_MODE=4'b1000;
    defparam comm_cmd_i3_LC_6_14_1.LUT_INIT=16'b1011100000110000;
    LogicCell40 comm_cmd_i3_LC_6_14_1 (
            .in0(N__50982),
            .in1(N__37536),
            .in2(N__47131),
            .in3(N__49878),
            .lcout(comm_cmd_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56060),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i30_4_lut_LC_6_14_2 .C_ON=1'b0;
    defparam \ADC_VAC.i30_4_lut_LC_6_14_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i30_4_lut_LC_6_14_2 .LUT_INIT=16'b1011100000010001;
    LogicCell40 \ADC_VAC.i30_4_lut_LC_6_14_2  (
            .in0(N__28698),
            .in1(N__21621),
            .in2(N__21713),
            .in3(N__21557),
            .lcout(\ADC_VAC.n17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.DTRIG_39_LC_6_14_4 .C_ON=1'b0;
    defparam \ADC_VAC.DTRIG_39_LC_6_14_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.DTRIG_39_LC_6_14_4 .LUT_INIT=16'b1010101011101000;
    LogicCell40 \ADC_VAC.DTRIG_39_LC_6_14_4  (
            .in0(N__28846),
            .in1(N__21558),
            .in2(N__21627),
            .in3(N__27722),
            .lcout(acadc_dtrig_v),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56060),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i16_LC_6_14_7 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i16_LC_6_14_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i16_LC_6_14_7 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i16_LC_6_14_7  (
            .in0(N__27721),
            .in1(N__26181),
            .in2(N__27964),
            .in3(N__25762),
            .lcout(buf_adcdata_vac_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56060),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.CS_37_LC_6_15_0 .C_ON=1'b0;
    defparam \ADC_VAC.CS_37_LC_6_15_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.CS_37_LC_6_15_0 .LUT_INIT=16'b0011001100110001;
    LogicCell40 \ADC_VAC.CS_37_LC_6_15_0  (
            .in0(N__21729),
            .in1(N__21633),
            .in2(N__27755),
            .in3(N__21714),
            .lcout(VAC_CS),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56074),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i26_LC_6_15_1 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i26_LC_6_15_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i26_LC_6_15_1 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i26_LC_6_15_1  (
            .in0(N__21436),
            .in1(N__27645),
            .in2(N__26207),
            .in3(N__28130),
            .lcout(cmd_rdadctmp_26_adj_1466),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56074),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.SCLK_35_LC_6_15_2 .C_ON=1'b0;
    defparam \ADC_VAC.SCLK_35_LC_6_15_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.SCLK_35_LC_6_15_2 .LUT_INIT=16'b1101000011100100;
    LogicCell40 \ADC_VAC.SCLK_35_LC_6_15_2  (
            .in0(N__27644),
            .in1(N__21619),
            .in2(N__21458),
            .in3(N__21554),
            .lcout(VAC_SCLK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56074),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i27_LC_6_15_3 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i27_LC_6_15_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i27_LC_6_15_3 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i27_LC_6_15_3  (
            .in0(N__25996),
            .in1(N__27646),
            .in2(N__21441),
            .in3(N__28131),
            .lcout(cmd_rdadctmp_27_adj_1465),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56074),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i18_LC_6_15_4 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i18_LC_6_15_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i18_LC_6_15_4 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC.ADC_DATA_i18_LC_6_15_4  (
            .in0(N__27883),
            .in1(N__27650),
            .in2(N__24130),
            .in3(N__21440),
            .lcout(buf_adcdata_vac_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56074),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i4_LC_6_15_6 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i4_LC_6_15_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i4_LC_6_15_6 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i4_LC_6_15_6  (
            .in0(N__28132),
            .in1(N__24713),
            .in2(N__21426),
            .in3(N__27651),
            .lcout(cmd_rdadctmp_4_adj_1488),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56074),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i10_LC_6_15_7 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i10_LC_6_15_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i10_LC_6_15_7 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i10_LC_6_15_7  (
            .in0(N__24313),
            .in1(N__29380),
            .in2(N__36344),
            .in3(N__38563),
            .lcout(cmd_rdadctmp_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56074),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.adc_state_i2_LC_6_16_1 .C_ON=1'b0;
    defparam \ADC_VAC.adc_state_i2_LC_6_16_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.adc_state_i2_LC_6_16_1 .LUT_INIT=16'b0011001110001000;
    LogicCell40 \ADC_VAC.adc_state_i2_LC_6_16_1  (
            .in0(N__27630),
            .in1(N__21612),
            .in2(_gnd_net_),
            .in3(N__21542),
            .lcout(DTRIG_N_958_adj_1493),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56084),
            .ce(N__21738),
            .sr(_gnd_net_));
    defparam \ADC_VAC.adc_state_i1_LC_6_16_2 .C_ON=1'b0;
    defparam \ADC_VAC.adc_state_i1_LC_6_16_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.adc_state_i1_LC_6_16_2 .LUT_INIT=16'b0101000001010101;
    LogicCell40 \ADC_VAC.adc_state_i1_LC_6_16_2  (
            .in0(N__21543),
            .in1(_gnd_net_),
            .in2(N__21626),
            .in3(N__27631),
            .lcout(adc_state_1_adj_1459),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56084),
            .ce(N__21738),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i1_2_lut_LC_6_16_3 .C_ON=1'b0;
    defparam \ADC_VAC.i1_2_lut_LC_6_16_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i1_2_lut_LC_6_16_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \ADC_VAC.i1_2_lut_LC_6_16_3  (
            .in0(_gnd_net_),
            .in1(N__21607),
            .in2(_gnd_net_),
            .in3(N__21539),
            .lcout(n21050),
            .ltout(n21050_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.i1_3_lut_LC_6_16_4 .C_ON=1'b0;
    defparam \ADC_VAC.i1_3_lut_LC_6_16_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VAC.i1_3_lut_LC_6_16_4 .LUT_INIT=16'b1111000000110000;
    LogicCell40 \ADC_VAC.i1_3_lut_LC_6_16_4  (
            .in0(_gnd_net_),
            .in1(N__21715),
            .in2(N__21663),
            .in3(N__27628),
            .lcout(n12850),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_223_LC_6_16_6.C_ON=1'b0;
    defparam i1_4_lut_adj_223_LC_6_16_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_223_LC_6_16_6.LUT_INIT=16'b0010001100110010;
    LogicCell40 i1_4_lut_adj_223_LC_6_16_6 (
            .in0(N__21541),
            .in1(N__21650),
            .in2(N__21625),
            .in3(N__27629),
            .lcout(n14_adj_1657),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_61_LC_6_16_7.C_ON=1'b0;
    defparam i1_2_lut_adj_61_LC_6_16_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_61_LC_6_16_7.LUT_INIT=16'b0000000011001100;
    LogicCell40 i1_2_lut_adj_61_LC_6_16_7 (
            .in0(_gnd_net_),
            .in1(N__21608),
            .in2(_gnd_net_),
            .in3(N__21540),
            .lcout(n21076),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i15_LC_6_17_0 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i15_LC_6_17_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i15_LC_6_17_0 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i15_LC_6_17_0  (
            .in0(N__38408),
            .in1(N__26281),
            .in2(N__21501),
            .in3(N__29337),
            .lcout(cmd_rdadctmp_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56092),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i6_4_lut_LC_6_17_1 .C_ON=1'b0;
    defparam \ADC_IAC.i6_4_lut_LC_6_17_1 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i6_4_lut_LC_6_17_1 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \ADC_IAC.i6_4_lut_LC_6_17_1  (
            .in0(N__24828),
            .in1(N__21830),
            .in2(N__21963),
            .in3(N__38406),
            .lcout(\ADC_IAC.n16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i19194_4_lut_LC_6_17_5 .C_ON=1'b0;
    defparam \ADC_IAC.i19194_4_lut_LC_6_17_5 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i19194_4_lut_LC_6_17_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \ADC_IAC.i19194_4_lut_LC_6_17_5  (
            .in0(N__21770),
            .in1(N__21785),
            .in2(N__21756),
            .in3(N__21800),
            .lcout(),
            .ltout(\ADC_IAC.n21458_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i19307_4_lut_LC_6_17_6 .C_ON=1'b0;
    defparam \ADC_IAC.i19307_4_lut_LC_6_17_6 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i19307_4_lut_LC_6_17_6 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \ADC_IAC.i19307_4_lut_LC_6_17_6  (
            .in0(N__21941),
            .in1(N__21816),
            .in2(N__21840),
            .in3(N__21837),
            .lcout(\ADC_IAC.n21457 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i19411_2_lut_LC_6_17_7 .C_ON=1'b0;
    defparam \ADC_IAC.i19411_2_lut_LC_6_17_7 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i19411_2_lut_LC_6_17_7 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \ADC_IAC.i19411_2_lut_LC_6_17_7  (
            .in0(_gnd_net_),
            .in1(N__38407),
            .in2(_gnd_net_),
            .in3(N__23757),
            .lcout(\ADC_IAC.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.bit_cnt_i0_LC_6_18_0 .C_ON=1'b1;
    defparam \ADC_IAC.bit_cnt_i0_LC_6_18_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i0_LC_6_18_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i0_LC_6_18_0  (
            .in0(_gnd_net_),
            .in1(N__21831),
            .in2(_gnd_net_),
            .in3(N__21819),
            .lcout(\ADC_IAC.bit_cnt_0 ),
            .ltout(),
            .carryin(bfn_6_18_0_),
            .carryout(\ADC_IAC.n19828 ),
            .clk(N__56096),
            .ce(N__21930),
            .sr(N__21915));
    defparam \ADC_IAC.bit_cnt_i1_LC_6_18_1 .C_ON=1'b1;
    defparam \ADC_IAC.bit_cnt_i1_LC_6_18_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i1_LC_6_18_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i1_LC_6_18_1  (
            .in0(_gnd_net_),
            .in1(N__21815),
            .in2(_gnd_net_),
            .in3(N__21804),
            .lcout(\ADC_IAC.bit_cnt_1 ),
            .ltout(),
            .carryin(\ADC_IAC.n19828 ),
            .carryout(\ADC_IAC.n19829 ),
            .clk(N__56096),
            .ce(N__21930),
            .sr(N__21915));
    defparam \ADC_IAC.bit_cnt_i2_LC_6_18_2 .C_ON=1'b1;
    defparam \ADC_IAC.bit_cnt_i2_LC_6_18_2 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i2_LC_6_18_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i2_LC_6_18_2  (
            .in0(_gnd_net_),
            .in1(N__21801),
            .in2(_gnd_net_),
            .in3(N__21789),
            .lcout(\ADC_IAC.bit_cnt_2 ),
            .ltout(),
            .carryin(\ADC_IAC.n19829 ),
            .carryout(\ADC_IAC.n19830 ),
            .clk(N__56096),
            .ce(N__21930),
            .sr(N__21915));
    defparam \ADC_IAC.bit_cnt_i3_LC_6_18_3 .C_ON=1'b1;
    defparam \ADC_IAC.bit_cnt_i3_LC_6_18_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i3_LC_6_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i3_LC_6_18_3  (
            .in0(_gnd_net_),
            .in1(N__21786),
            .in2(_gnd_net_),
            .in3(N__21774),
            .lcout(\ADC_IAC.bit_cnt_3 ),
            .ltout(),
            .carryin(\ADC_IAC.n19830 ),
            .carryout(\ADC_IAC.n19831 ),
            .clk(N__56096),
            .ce(N__21930),
            .sr(N__21915));
    defparam \ADC_IAC.bit_cnt_i4_LC_6_18_4 .C_ON=1'b1;
    defparam \ADC_IAC.bit_cnt_i4_LC_6_18_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i4_LC_6_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i4_LC_6_18_4  (
            .in0(_gnd_net_),
            .in1(N__21771),
            .in2(_gnd_net_),
            .in3(N__21759),
            .lcout(\ADC_IAC.bit_cnt_4 ),
            .ltout(),
            .carryin(\ADC_IAC.n19831 ),
            .carryout(\ADC_IAC.n19832 ),
            .clk(N__56096),
            .ce(N__21930),
            .sr(N__21915));
    defparam \ADC_IAC.bit_cnt_i5_LC_6_18_5 .C_ON=1'b1;
    defparam \ADC_IAC.bit_cnt_i5_LC_6_18_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i5_LC_6_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i5_LC_6_18_5  (
            .in0(_gnd_net_),
            .in1(N__21755),
            .in2(_gnd_net_),
            .in3(N__21741),
            .lcout(\ADC_IAC.bit_cnt_5 ),
            .ltout(),
            .carryin(\ADC_IAC.n19832 ),
            .carryout(\ADC_IAC.n19833 ),
            .clk(N__56096),
            .ce(N__21930),
            .sr(N__21915));
    defparam \ADC_IAC.bit_cnt_i6_LC_6_18_6 .C_ON=1'b1;
    defparam \ADC_IAC.bit_cnt_i6_LC_6_18_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i6_LC_6_18_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i6_LC_6_18_6  (
            .in0(_gnd_net_),
            .in1(N__21962),
            .in2(_gnd_net_),
            .in3(N__21948),
            .lcout(\ADC_IAC.bit_cnt_6 ),
            .ltout(),
            .carryin(\ADC_IAC.n19833 ),
            .carryout(\ADC_IAC.n19834 ),
            .clk(N__56096),
            .ce(N__21930),
            .sr(N__21915));
    defparam \ADC_IAC.bit_cnt_i7_LC_6_18_7 .C_ON=1'b0;
    defparam \ADC_IAC.bit_cnt_i7_LC_6_18_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.bit_cnt_i7_LC_6_18_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_IAC.bit_cnt_i7_LC_6_18_7  (
            .in0(_gnd_net_),
            .in1(N__21942),
            .in2(_gnd_net_),
            .in3(N__21945),
            .lcout(\ADC_IAC.bit_cnt_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56096),
            .ce(N__21930),
            .sr(N__21915));
    defparam \ADC_IAC.i1_4_lut_LC_6_19_1 .C_ON=1'b0;
    defparam \ADC_IAC.i1_4_lut_LC_6_19_1 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i1_4_lut_LC_6_19_1 .LUT_INIT=16'b0000000101000100;
    LogicCell40 \ADC_IAC.i1_4_lut_LC_6_19_1  (
            .in0(N__38457),
            .in1(N__24935),
            .in2(N__24615),
            .in3(N__24852),
            .lcout(\ADC_IAC.n12698 ),
            .ltout(\ADC_IAC.n12698_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i12498_2_lut_LC_6_19_2 .C_ON=1'b0;
    defparam \ADC_IAC.i12498_2_lut_LC_6_19_2 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i12498_2_lut_LC_6_19_2 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \ADC_IAC.i12498_2_lut_LC_6_19_2  (
            .in0(N__24939),
            .in1(_gnd_net_),
            .in2(N__21918),
            .in3(_gnd_net_),
            .lcout(\ADC_IAC.n15014 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_rst_I_0_1_lut_LC_6_19_3.C_ON=1'b0;
    defparam acadc_rst_I_0_1_lut_LC_6_19_3.SEQ_MODE=4'b0000;
    defparam acadc_rst_I_0_1_lut_LC_6_19_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 acadc_rst_I_0_1_lut_LC_6_19_3 (
            .in0(N__35731),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(AC_ADC_SYNC),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_225_LC_6_19_4.C_ON=1'b0;
    defparam i1_4_lut_adj_225_LC_6_19_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_225_LC_6_19_4.LUT_INIT=16'b0010001100110010;
    LogicCell40 i1_4_lut_adj_225_LC_6_19_4 (
            .in0(N__24853),
            .in1(N__21869),
            .in2(N__24942),
            .in3(N__38458),
            .lcout(),
            .ltout(n14_adj_1662_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.CS_37_LC_6_19_5 .C_ON=1'b0;
    defparam \ADC_IAC.CS_37_LC_6_19_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.CS_37_LC_6_19_5 .LUT_INIT=16'b0000111000001111;
    LogicCell40 \ADC_IAC.CS_37_LC_6_19_5  (
            .in0(N__38459),
            .in1(N__24606),
            .in2(N__21882),
            .in3(N__23799),
            .lcout(IAC_CS),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56099),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i3_LC_7_5_0 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i3_LC_7_5_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i3_LC_7_5_0 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \ADC_VDC.ADC_DATA_i3_LC_7_5_0  (
            .in0(N__24057),
            .in1(N__51413),
            .in2(N__22874),
            .in3(N__31626),
            .lcout(buf_adcdata_vdc_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42373),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.CS_28_LC_7_6_3 .C_ON=1'b0;
    defparam \CLK_DDS.CS_28_LC_7_6_3 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.CS_28_LC_7_6_3 .LUT_INIT=16'b0010001001110111;
    LogicCell40 \CLK_DDS.CS_28_LC_7_6_3  (
            .in0(N__30102),
            .in1(N__29767),
            .in2(_gnd_net_),
            .in3(N__29942),
            .lcout(DDS_CS1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55951),
            .ce(N__30123),
            .sr(_gnd_net_));
    defparam \RTD.cfg_tmp_i1_LC_7_7_0 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i1_LC_7_7_0 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i1_LC_7_7_0 .LUT_INIT=16'b1110101001000000;
    LogicCell40 \RTD.cfg_tmp_i1_LC_7_7_0  (
            .in0(N__22217),
            .in1(N__22412),
            .in2(N__39600),
            .in3(N__21981),
            .lcout(\RTD.cfg_tmp_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40622),
            .ce(N__21975),
            .sr(N__21969));
    defparam \RTD.cfg_tmp_i2_LC_7_7_1 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i2_LC_7_7_1 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i2_LC_7_7_1 .LUT_INIT=16'b1100110010100000;
    LogicCell40 \RTD.cfg_tmp_i2_LC_7_7_1  (
            .in0(N__22410),
            .in1(N__22461),
            .in2(N__23334),
            .in3(N__22223),
            .lcout(\RTD.cfg_tmp_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40622),
            .ce(N__21975),
            .sr(N__21969));
    defparam \RTD.cfg_tmp_i3_LC_7_7_2 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i3_LC_7_7_2 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i3_LC_7_7_2 .LUT_INIT=16'b1110010010100000;
    LogicCell40 \RTD.cfg_tmp_i3_LC_7_7_2  (
            .in0(N__22218),
            .in1(N__22413),
            .in2(N__22455),
            .in3(N__25946),
            .lcout(\RTD.cfg_tmp_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40622),
            .ce(N__21975),
            .sr(N__21969));
    defparam \RTD.cfg_tmp_i4_LC_7_7_3 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i4_LC_7_7_3 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i4_LC_7_7_3 .LUT_INIT=16'b1100110010100000;
    LogicCell40 \RTD.cfg_tmp_i4_LC_7_7_3  (
            .in0(N__35010),
            .in1(N__22446),
            .in2(N__22421),
            .in3(N__22224),
            .lcout(\RTD.cfg_tmp_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40622),
            .ce(N__21975),
            .sr(N__21969));
    defparam \RTD.cfg_tmp_i5_LC_7_7_4 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i5_LC_7_7_4 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i5_LC_7_7_4 .LUT_INIT=16'b1101100010001000;
    LogicCell40 \RTD.cfg_tmp_i5_LC_7_7_4  (
            .in0(N__22221),
            .in1(N__22440),
            .in2(N__22422),
            .in3(N__34939),
            .lcout(\RTD.cfg_tmp_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40622),
            .ce(N__21975),
            .sr(N__21969));
    defparam \RTD.cfg_tmp_i6_LC_7_7_5 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i6_LC_7_7_5 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i6_LC_7_7_5 .LUT_INIT=16'b1110110000100000;
    LogicCell40 \RTD.cfg_tmp_i6_LC_7_7_5  (
            .in0(N__22411),
            .in1(N__22220),
            .in2(N__27077),
            .in3(N__22434),
            .lcout(\RTD.cfg_tmp_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40622),
            .ce(N__21975),
            .sr(N__21969));
    defparam \RTD.cfg_tmp_i7_LC_7_7_6 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i7_LC_7_7_6 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i7_LC_7_7_6 .LUT_INIT=16'b1110101001000000;
    LogicCell40 \RTD.cfg_tmp_i7_LC_7_7_6  (
            .in0(N__22219),
            .in1(N__22414),
            .in2(N__27024),
            .in3(N__22428),
            .lcout(\RTD.cfg_tmp_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40622),
            .ce(N__21975),
            .sr(N__21969));
    defparam \RTD.cfg_tmp_i0_LC_7_7_7 .C_ON=1'b0;
    defparam \RTD.cfg_tmp_i0_LC_7_7_7 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_tmp_i0_LC_7_7_7 .LUT_INIT=16'b1100110010100000;
    LogicCell40 \RTD.cfg_tmp_i0_LC_7_7_7  (
            .in0(N__22409),
            .in1(N__22235),
            .in2(N__25740),
            .in3(N__22222),
            .lcout(\RTD.cfg_tmp_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40622),
            .ce(N__21975),
            .sr(N__21969));
    defparam \RTD.cfg_buf_i4_LC_7_8_0 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i4_LC_7_8_0 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i4_LC_7_8_0 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \RTD.cfg_buf_i4_LC_7_8_0  (
            .in0(N__22731),
            .in1(N__22949),
            .in2(N__23009),
            .in3(N__35008),
            .lcout(\RTD.cfg_buf_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40607),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i5_LC_7_8_1 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i5_LC_7_8_1 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i5_LC_7_8_1 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \RTD.cfg_buf_i5_LC_7_8_1  (
            .in0(N__22755),
            .in1(N__23005),
            .in2(N__22968),
            .in3(N__34940),
            .lcout(\RTD.cfg_buf_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40607),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i3_4_lut_adj_7_LC_7_8_2 .C_ON=1'b0;
    defparam \RTD.i3_4_lut_adj_7_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \RTD.i3_4_lut_adj_7_LC_7_8_2 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \RTD.i3_4_lut_adj_7_LC_7_8_2  (
            .in0(N__34941),
            .in1(N__22754),
            .in2(N__25947),
            .in3(N__22739),
            .lcout(\RTD.n11_adj_1444 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i3_LC_7_8_3 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i3_LC_7_8_3 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i3_LC_7_8_3 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \RTD.cfg_buf_i3_LC_7_8_3  (
            .in0(N__22740),
            .in1(N__22998),
            .in2(N__22967),
            .in3(N__25942),
            .lcout(\RTD.cfg_buf_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40607),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i2_LC_7_8_4 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i2_LC_7_8_4 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i2_LC_7_8_4 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \RTD.cfg_buf_i2_LC_7_8_4  (
            .in0(N__22722),
            .in1(N__22950),
            .in2(N__23010),
            .in3(N__23323),
            .lcout(\RTD.cfg_buf_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40607),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i2_4_lut_LC_7_8_5 .C_ON=1'b0;
    defparam \RTD.i2_4_lut_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \RTD.i2_4_lut_LC_7_8_5 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \RTD.i2_4_lut_LC_7_8_5  (
            .in0(N__35009),
            .in1(N__22730),
            .in2(N__23330),
            .in3(N__22721),
            .lcout(\RTD.n10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i22_4_lut_LC_7_8_6 .C_ON=1'b0;
    defparam \RTD.i22_4_lut_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \RTD.i22_4_lut_LC_7_8_6 .LUT_INIT=16'b1100000011100010;
    LogicCell40 \RTD.i22_4_lut_LC_7_8_6  (
            .in0(N__22707),
            .in1(N__22694),
            .in2(N__22545),
            .in3(N__22526),
            .lcout(\RTD.n13090 ),
            .ltout(\RTD.n13090_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i1_LC_7_8_7 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i1_LC_7_8_7 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i1_LC_7_8_7 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \RTD.cfg_buf_i1_LC_7_8_7  (
            .in0(N__22948),
            .in1(N__39596),
            .in2(N__22491),
            .in3(N__22488),
            .lcout(\RTD.cfg_buf_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40607),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.i4_4_lut_LC_7_9_0 .C_ON=1'b0;
    defparam \RTD.i4_4_lut_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \RTD.i4_4_lut_LC_7_9_0 .LUT_INIT=16'b0110111111110110;
    LogicCell40 \RTD.i4_4_lut_LC_7_9_0  (
            .in0(N__27017),
            .in1(N__22469),
            .in2(N__39595),
            .in3(N__22487),
            .lcout(\RTD.n12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i7_LC_7_9_1 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i7_LC_7_9_1 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i7_LC_7_9_1 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \RTD.cfg_buf_i7_LC_7_9_1  (
            .in0(N__22470),
            .in1(N__27016),
            .in2(N__22970),
            .in3(N__23007),
            .lcout(\RTD.cfg_buf_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40621),
            .ce(),
            .sr(_gnd_net_));
    defparam \RTD.cfg_buf_i0_LC_7_9_2 .C_ON=1'b0;
    defparam \RTD.cfg_buf_i0_LC_7_9_2 .SEQ_MODE=4'b1000;
    defparam \RTD.cfg_buf_i0_LC_7_9_2 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \RTD.cfg_buf_i0_LC_7_9_2  (
            .in0(N__25735),
            .in1(N__23006),
            .in2(N__22969),
            .in3(N__22901),
            .lcout(\RTD.cfg_buf_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__40621),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_1_i20_3_lut_LC_7_9_3.C_ON=1'b0;
    defparam mux_128_Mux_1_i20_3_lut_LC_7_9_3.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_1_i20_3_lut_LC_7_9_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_128_Mux_1_i20_3_lut_LC_7_9_3 (
            .in0(N__22887),
            .in1(N__39585),
            .in2(_gnd_net_),
            .in3(N__57196),
            .lcout(n20_adj_1693),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_3_i19_3_lut_LC_7_9_4.C_ON=1'b0;
    defparam mux_130_Mux_3_i19_3_lut_LC_7_9_4.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_3_i19_3_lut_LC_7_9_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_130_Mux_3_i19_3_lut_LC_7_9_4 (
            .in0(N__57198),
            .in1(N__22875),
            .in2(_gnd_net_),
            .in3(N__23258),
            .lcout(),
            .ltout(n19_adj_1609_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_3_i22_3_lut_LC_7_9_5.C_ON=1'b0;
    defparam mux_130_Mux_3_i22_3_lut_LC_7_9_5.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_3_i22_3_lut_LC_7_9_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 mux_130_Mux_3_i22_3_lut_LC_7_9_5 (
            .in0(_gnd_net_),
            .in1(N__22853),
            .in2(N__22824),
            .in3(N__47500),
            .lcout(n22_adj_1610),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22407_bdd_4_lut_LC_7_9_6.C_ON=1'b0;
    defparam n22407_bdd_4_lut_LC_7_9_6.SEQ_MODE=4'b0000;
    defparam n22407_bdd_4_lut_LC_7_9_6.LUT_INIT=16'b1111101001000100;
    LogicCell40 n22407_bdd_4_lut_LC_7_9_6 (
            .in0(N__47501),
            .in1(N__23706),
            .in2(N__23697),
            .in3(N__23175),
            .lcout(n22410),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19857_LC_7_9_7.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19857_LC_7_9_7.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19857_LC_7_9_7.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_cmd_0__bdd_4_lut_19857_LC_7_9_7 (
            .in0(N__27060),
            .in1(N__57197),
            .in2(N__22821),
            .in3(N__46256),
            .lcout(n22629),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i2_LC_7_10_0 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i2_LC_7_10_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i2_LC_7_10_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i2_LC_7_10_0  (
            .in0(N__28001),
            .in1(N__27850),
            .in2(N__22803),
            .in3(N__23159),
            .lcout(buf_adcdata_vac_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55987),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_1_i19_3_lut_LC_7_10_1.C_ON=1'b0;
    defparam mux_129_Mux_1_i19_3_lut_LC_7_10_1.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_1_i19_3_lut_LC_7_10_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_129_Mux_1_i19_3_lut_LC_7_10_1 (
            .in0(N__25437),
            .in1(N__23561),
            .in2(_gnd_net_),
            .in3(N__57091),
            .lcout(n19_adj_1652),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.MOSI_31_LC_7_10_2 .C_ON=1'b0;
    defparam \CLK_DDS.MOSI_31_LC_7_10_2 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.MOSI_31_LC_7_10_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \CLK_DDS.MOSI_31_LC_7_10_2  (
            .in0(N__24396),
            .in1(N__22766),
            .in2(_gnd_net_),
            .in3(N__29822),
            .lcout(DDS_MOSI1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55987),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19678_LC_7_10_3.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19678_LC_7_10_3.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19678_LC_7_10_3.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_19678_LC_7_10_3 (
            .in0(N__24099),
            .in1(N__46257),
            .in2(N__23184),
            .in3(N__47451),
            .lcout(n22407),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_2_i19_3_lut_LC_7_10_4.C_ON=1'b0;
    defparam mux_130_Mux_2_i19_3_lut_LC_7_10_4.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_2_i19_3_lut_LC_7_10_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_130_Mux_2_i19_3_lut_LC_7_10_4 (
            .in0(N__57092),
            .in1(N__25647),
            .in2(_gnd_net_),
            .in3(N__23158),
            .lcout(),
            .ltout(n19_adj_1612_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_2_i22_3_lut_LC_7_10_5.C_ON=1'b0;
    defparam mux_130_Mux_2_i22_3_lut_LC_7_10_5.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_2_i22_3_lut_LC_7_10_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 mux_130_Mux_2_i22_3_lut_LC_7_10_5 (
            .in0(_gnd_net_),
            .in1(N__24283),
            .in2(N__23145),
            .in3(N__47452),
            .lcout(n22_adj_1613),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i6_LC_7_10_6 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i6_LC_7_10_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i6_LC_7_10_6 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i6_LC_7_10_6  (
            .in0(N__28002),
            .in1(N__27851),
            .in2(N__23064),
            .in3(N__23137),
            .lcout(buf_adcdata_vac_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55987),
            .ce(),
            .sr(_gnd_net_));
    defparam i15464_2_lut_3_lut_LC_7_11_0.C_ON=1'b0;
    defparam i15464_2_lut_3_lut_LC_7_11_0.SEQ_MODE=4'b0000;
    defparam i15464_2_lut_3_lut_LC_7_11_0.LUT_INIT=16'b0000000000100010;
    LogicCell40 i15464_2_lut_3_lut_LC_7_11_0 (
            .in0(N__45848),
            .in1(N__54884),
            .in2(_gnd_net_),
            .in3(N__54555),
            .lcout(n14_adj_1574),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22629_bdd_4_lut_LC_7_11_1.C_ON=1'b0;
    defparam n22629_bdd_4_lut_LC_7_11_1.SEQ_MODE=4'b0000;
    defparam n22629_bdd_4_lut_LC_7_11_1.LUT_INIT=16'b1100110011100010;
    LogicCell40 n22629_bdd_4_lut_LC_7_11_1 (
            .in0(N__23092),
            .in1(N__23073),
            .in2(N__25686),
            .in3(N__46159),
            .lcout(n21237),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i2_LC_7_11_2.C_ON=1'b0;
    defparam buf_cfgRTD_i2_LC_7_11_2.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i2_LC_7_11_2.LUT_INIT=16'b0011000010101010;
    LogicCell40 buf_cfgRTD_i2_LC_7_11_2 (
            .in0(N__23314),
            .in1(N__49312),
            .in2(N__45868),
            .in3(N__39663),
            .lcout(buf_cfgRTD_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56000),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i16_LC_7_11_3 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i16_LC_7_11_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i16_LC_7_11_3 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i16_LC_7_11_3  (
            .in0(N__27848),
            .in1(N__26221),
            .in2(N__23030),
            .in3(N__28268),
            .lcout(cmd_rdadctmp_16_adj_1476),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56000),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i15_LC_7_11_4 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i15_LC_7_11_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i15_LC_7_11_4 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i15_LC_7_11_4  (
            .in0(N__28267),
            .in1(N__23023),
            .in2(N__23060),
            .in3(N__27849),
            .lcout(cmd_rdadctmp_15_adj_1477),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56000),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_6_i30_3_lut_LC_7_11_5.C_ON=1'b0;
    defparam mux_130_Mux_6_i30_3_lut_LC_7_11_5.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_6_i30_3_lut_LC_7_11_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_130_Mux_6_i30_3_lut_LC_7_11_5 (
            .in0(N__47158),
            .in1(N__23403),
            .in2(_gnd_net_),
            .in3(N__23388),
            .lcout(n30_adj_1602),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_2_i30_3_lut_LC_7_11_6.C_ON=1'b0;
    defparam mux_130_Mux_2_i30_3_lut_LC_7_11_6.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_2_i30_3_lut_LC_7_11_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_130_Mux_2_i30_3_lut_LC_7_11_6 (
            .in0(N__23379),
            .in1(N__23358),
            .in2(_gnd_net_),
            .in3(N__47159),
            .lcout(n30_adj_1614),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_2_i20_3_lut_LC_7_11_7.C_ON=1'b0;
    defparam mux_128_Mux_2_i20_3_lut_LC_7_11_7.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_2_i20_3_lut_LC_7_11_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_128_Mux_2_i20_3_lut_LC_7_11_7 (
            .in0(N__56937),
            .in1(N__23352),
            .in2(_gnd_net_),
            .in3(N__23313),
            .lcout(n20_adj_1684),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i17_LC_7_12_0 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i17_LC_7_12_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i17_LC_7_12_0 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i17_LC_7_12_0  (
            .in0(N__23461),
            .in1(N__27794),
            .in2(N__26234),
            .in3(N__28246),
            .lcout(cmd_rdadctmp_17_adj_1475),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56017),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i3_LC_7_12_1 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i3_LC_7_12_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i3_LC_7_12_1 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i3_LC_7_12_1  (
            .in0(N__27791),
            .in1(N__27989),
            .in2(N__23298),
            .in3(N__23257),
            .lcout(buf_adcdata_vac_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56017),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i5_LC_7_12_2 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i5_LC_7_12_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i5_LC_7_12_2 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i5_LC_7_12_2  (
            .in0(N__27990),
            .in1(N__27792),
            .in2(N__23235),
            .in3(N__24257),
            .lcout(buf_adcdata_vac_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56017),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i1_LC_7_12_3.C_ON=1'b0;
    defparam comm_cmd_i1_LC_7_12_3.SEQ_MODE=4'b1000;
    defparam comm_cmd_i1_LC_7_12_3.LUT_INIT=16'b1011001110000000;
    LogicCell40 comm_cmd_i1_LC_7_12_3 (
            .in0(N__50981),
            .in1(N__37522),
            .in2(N__49745),
            .in3(N__46224),
            .lcout(comm_cmd_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56017),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i30_LC_7_12_4 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i30_LC_7_12_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i30_LC_7_12_4 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i30_LC_7_12_4  (
            .in0(N__23200),
            .in1(N__27795),
            .in2(N__23448),
            .in3(N__28247),
            .lcout(cmd_rdadctmp_30_adj_1462),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56017),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i21_LC_7_12_5 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i21_LC_7_12_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i21_LC_7_12_5 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC.ADC_DATA_i21_LC_7_12_5  (
            .in0(N__27790),
            .in1(N__27988),
            .in2(N__27421),
            .in3(N__23447),
            .lcout(buf_adcdata_vac_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56017),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i9_LC_7_12_6 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i9_LC_7_12_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i9_LC_7_12_6 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i9_LC_7_12_6  (
            .in0(N__27991),
            .in1(N__27793),
            .in2(N__23466),
            .in3(N__23560),
            .lcout(buf_adcdata_vac_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56017),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i12_LC_7_13_0 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i12_LC_7_13_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i12_LC_7_13_0 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i12_LC_7_13_0  (
            .in0(N__38558),
            .in1(N__23509),
            .in2(N__23538),
            .in3(N__29363),
            .lcout(cmd_rdadctmp_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56031),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i8_LC_7_13_1 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i8_LC_7_13_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i8_LC_7_13_1 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i8_LC_7_13_1  (
            .in0(N__29362),
            .in1(N__23482),
            .in2(N__23667),
            .in3(N__38559),
            .lcout(cmd_rdadctmp_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56031),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_dtrig_i_I_0_2_lut_LC_7_13_2.C_ON=1'b0;
    defparam acadc_dtrig_i_I_0_2_lut_LC_7_13_2.SEQ_MODE=4'b0000;
    defparam acadc_dtrig_i_I_0_2_lut_LC_7_13_2.LUT_INIT=16'b1100110000000000;
    LogicCell40 acadc_dtrig_i_I_0_2_lut_LC_7_13_2 (
            .in0(_gnd_net_),
            .in1(N__28826),
            .in2(_gnd_net_),
            .in3(N__28785),
            .lcout(iac_raw_buf_N_776),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i18_LC_7_13_3 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i18_LC_7_13_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i18_LC_7_13_3 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i18_LC_7_13_3  (
            .in0(N__27821),
            .in1(N__23465),
            .in2(N__26126),
            .in3(N__28254),
            .lcout(cmd_rdadctmp_18_adj_1474),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56031),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.DTRIG_39_LC_7_13_4 .C_ON=1'b0;
    defparam \ADC_IAC.DTRIG_39_LC_7_13_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.DTRIG_39_LC_7_13_4 .LUT_INIT=16'b1111111001000000;
    LogicCell40 \ADC_IAC.DTRIG_39_LC_7_13_4  (
            .in0(N__38557),
            .in1(N__24854),
            .in2(N__24940),
            .in3(N__28786),
            .lcout(acadc_dtrig_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56031),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i29_LC_7_13_5 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i29_LC_7_13_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i29_LC_7_13_5 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i29_LC_7_13_5  (
            .in0(N__27822),
            .in1(N__24412),
            .in2(N__23443),
            .in3(N__28256),
            .lcout(cmd_rdadctmp_29_adj_1463),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56031),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i28_LC_7_13_6 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i28_LC_7_13_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i28_LC_7_13_6 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i28_LC_7_13_6  (
            .in0(N__28255),
            .in1(N__27823),
            .in2(N__24416),
            .in3(N__26003),
            .lcout(cmd_rdadctmp_28_adj_1464),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56031),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i1_LC_7_13_7 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i1_LC_7_13_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i1_LC_7_13_7 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i1_LC_7_13_7  (
            .in0(N__27820),
            .in1(N__27965),
            .in2(N__23424),
            .in3(N__32162),
            .lcout(buf_adcdata_vac_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56031),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i10_LC_7_14_0 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i10_LC_7_14_0 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i10_LC_7_14_0 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \CLK_DDS.tmp_buf_i10_LC_7_14_0  (
            .in0(N__30094),
            .in1(N__29845),
            .in2(N__23586),
            .in3(N__30873),
            .lcout(\CLK_DDS.tmp_buf_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56047),
            .ce(N__30147),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i11_LC_7_14_1 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i11_LC_7_14_1 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i11_LC_7_14_1 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLK_DDS.tmp_buf_i11_LC_7_14_1  (
            .in0(N__29846),
            .in1(N__30098),
            .in2(N__23634),
            .in3(N__26442),
            .lcout(\CLK_DDS.tmp_buf_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56047),
            .ce(N__30147),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i12_LC_7_14_2 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i12_LC_7_14_2 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i12_LC_7_14_2 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \CLK_DDS.tmp_buf_i12_LC_7_14_2  (
            .in0(N__30095),
            .in1(N__29847),
            .in2(N__23625),
            .in3(N__36287),
            .lcout(\CLK_DDS.tmp_buf_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56047),
            .ce(N__30147),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i13_LC_7_14_3 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i13_LC_7_14_3 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i13_LC_7_14_3 .LUT_INIT=16'b0000110010101010;
    LogicCell40 \CLK_DDS.tmp_buf_i13_LC_7_14_3  (
            .in0(N__34960),
            .in1(N__23616),
            .in2(N__29872),
            .in3(N__30101),
            .lcout(\CLK_DDS.tmp_buf_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56047),
            .ce(N__30147),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i14_LC_7_14_4 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i14_LC_7_14_4 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i14_LC_7_14_4 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \CLK_DDS.tmp_buf_i14_LC_7_14_4  (
            .in0(N__30096),
            .in1(N__29851),
            .in2(N__23607),
            .in3(N__35637),
            .lcout(\CLK_DDS.tmp_buf_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56047),
            .ce(N__30147),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i15_LC_7_14_5 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i15_LC_7_14_5 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i15_LC_7_14_5 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLK_DDS.tmp_buf_i15_LC_7_14_5  (
            .in0(N__29852),
            .in1(N__30099),
            .in2(N__23595),
            .in3(N__30897),
            .lcout(tmp_buf_15_adj_1497),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56047),
            .ce(N__30147),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i9_LC_7_14_6 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i9_LC_7_14_6 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i9_LC_7_14_6 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \CLK_DDS.tmp_buf_i9_LC_7_14_6  (
            .in0(N__30097),
            .in1(N__29854),
            .in2(N__23577),
            .in3(N__32526),
            .lcout(\CLK_DDS.tmp_buf_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56047),
            .ce(N__30147),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i8_LC_7_14_7 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i8_LC_7_14_7 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i8_LC_7_14_7 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLK_DDS.tmp_buf_i8_LC_7_14_7  (
            .in0(N__29853),
            .in1(N__30100),
            .in2(N__24540),
            .in3(N__39103),
            .lcout(\CLK_DDS.tmp_buf_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56047),
            .ce(N__30147),
            .sr(_gnd_net_));
    defparam \SIG_DDS.bit_cnt_i3_LC_7_15_0 .C_ON=1'b0;
    defparam \SIG_DDS.bit_cnt_i3_LC_7_15_0 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.bit_cnt_i3_LC_7_15_0 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \SIG_DDS.bit_cnt_i3_LC_7_15_0  (
            .in0(N__24474),
            .in1(N__24441),
            .in2(N__24498),
            .in3(N__36605),
            .lcout(\SIG_DDS.bit_cnt_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56061),
            .ce(N__44517),
            .sr(N__24645));
    defparam \SIG_DDS.bit_cnt_i1_LC_7_15_1 .C_ON=1'b0;
    defparam \SIG_DDS.bit_cnt_i1_LC_7_15_1 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.bit_cnt_i1_LC_7_15_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \SIG_DDS.bit_cnt_i1_LC_7_15_1  (
            .in0(N__24439),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24497),
            .lcout(\SIG_DDS.bit_cnt_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56061),
            .ce(N__44517),
            .sr(N__24645));
    defparam i18636_3_lut_LC_7_15_3.C_ON=1'b0;
    defparam i18636_3_lut_LC_7_15_3.SEQ_MODE=4'b0000;
    defparam i18636_3_lut_LC_7_15_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 i18636_3_lut_LC_7_15_3 (
            .in0(N__23733),
            .in1(N__28389),
            .in2(_gnd_net_),
            .in3(N__46258),
            .lcout(n21363),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.bit_cnt_i2_LC_7_15_4 .C_ON=1'b0;
    defparam \SIG_DDS.bit_cnt_i2_LC_7_15_4 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.bit_cnt_i2_LC_7_15_4 .LUT_INIT=16'b0110011010101010;
    LogicCell40 \SIG_DDS.bit_cnt_i2_LC_7_15_4  (
            .in0(N__24473),
            .in1(N__24493),
            .in2(_gnd_net_),
            .in3(N__24440),
            .lcout(\SIG_DDS.bit_cnt_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56061),
            .ce(N__44517),
            .sr(N__24645));
    defparam mux_128_Mux_1_i16_3_lut_LC_7_15_5.C_ON=1'b0;
    defparam mux_128_Mux_1_i16_3_lut_LC_7_15_5.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_1_i16_3_lut_LC_7_15_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_128_Mux_1_i16_3_lut_LC_7_15_5 (
            .in0(N__57269),
            .in1(N__32525),
            .in2(_gnd_net_),
            .in3(N__31253),
            .lcout(n16_adj_1690),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_1_i17_3_lut_LC_7_15_6.C_ON=1'b0;
    defparam mux_128_Mux_1_i17_3_lut_LC_7_15_6.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_1_i17_3_lut_LC_7_15_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_128_Mux_1_i17_3_lut_LC_7_15_6 (
            .in0(N__24749),
            .in1(N__26090),
            .in2(_gnd_net_),
            .in3(N__57268),
            .lcout(n17_adj_1691),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.adc_state_i2_LC_7_16_1 .C_ON=1'b0;
    defparam \ADC_IAC.adc_state_i2_LC_7_16_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.adc_state_i2_LC_7_16_1 .LUT_INIT=16'b0011001110001000;
    LogicCell40 \ADC_IAC.adc_state_i2_LC_7_16_1  (
            .in0(N__38447),
            .in1(N__24908),
            .in2(_gnd_net_),
            .in3(N__24840),
            .lcout(DTRIG_N_958),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56075),
            .ce(N__23682),
            .sr(_gnd_net_));
    defparam \ADC_IAC.adc_state_i1_LC_7_16_2 .C_ON=1'b0;
    defparam \ADC_IAC.adc_state_i1_LC_7_16_2 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.adc_state_i1_LC_7_16_2 .LUT_INIT=16'b0101000001010101;
    LogicCell40 \ADC_IAC.adc_state_i1_LC_7_16_2  (
            .in0(N__24841),
            .in1(_gnd_net_),
            .in2(N__24927),
            .in3(N__38448),
            .lcout(adc_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56075),
            .ce(N__23682),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_52_LC_7_16_7.C_ON=1'b0;
    defparam i1_2_lut_adj_52_LC_7_16_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_52_LC_7_16_7.LUT_INIT=16'b0000000011001100;
    LogicCell40 i1_2_lut_adj_52_LC_7_16_7 (
            .in0(_gnd_net_),
            .in1(N__24904),
            .in2(_gnd_net_),
            .in3(N__24839),
            .lcout(n21079),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.adc_state_i0_LC_7_17_4 .C_ON=1'b0;
    defparam \ADC_IAC.adc_state_i0_LC_7_17_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.adc_state_i0_LC_7_17_4 .LUT_INIT=16'b0001111100010000;
    LogicCell40 \ADC_IAC.adc_state_i0_LC_7_17_4  (
            .in0(N__38446),
            .in1(N__24846),
            .in2(N__24928),
            .in3(N__23673),
            .lcout(adc_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56085),
            .ce(N__25008),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i7_LC_7_18_0 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i7_LC_7_18_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i7_LC_7_18_0 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i7_LC_7_18_0  (
            .in0(N__23657),
            .in1(N__29328),
            .in2(N__23646),
            .in3(N__38401),
            .lcout(cmd_rdadctmp_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56093),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i6_LC_7_18_1 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i6_LC_7_18_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i6_LC_7_18_1 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i6_LC_7_18_1  (
            .in0(N__38399),
            .in1(N__23642),
            .in2(N__29374),
            .in3(N__23766),
            .lcout(cmd_rdadctmp_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56093),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i3_LC_7_18_2 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i3_LC_7_18_2 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i3_LC_7_18_2 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i3_LC_7_18_2  (
            .in0(N__23789),
            .in1(N__29326),
            .in2(N__38564),
            .in3(N__24989),
            .lcout(cmd_rdadctmp_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56093),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_226_LC_7_18_3.C_ON=1'b0;
    defparam i1_2_lut_adj_226_LC_7_18_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_226_LC_7_18_3.LUT_INIT=16'b0011001100000000;
    LogicCell40 i1_2_lut_adj_226_LC_7_18_3 (
            .in0(_gnd_net_),
            .in1(N__24918),
            .in2(_gnd_net_),
            .in3(N__24850),
            .lcout(n21082),
            .ltout(n21082_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i1_3_lut_LC_7_18_4 .C_ON=1'b0;
    defparam \ADC_IAC.i1_3_lut_LC_7_18_4 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i1_3_lut_LC_7_18_4 .LUT_INIT=16'b1111000000110000;
    LogicCell40 \ADC_IAC.i1_3_lut_LC_7_18_4  (
            .in0(_gnd_net_),
            .in1(N__24616),
            .in2(N__23793),
            .in3(N__38397),
            .lcout(n12771),
            .ltout(n12771_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i4_LC_7_18_5 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i4_LC_7_18_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i4_LC_7_18_5 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i4_LC_7_18_5  (
            .in0(N__38398),
            .in1(N__23790),
            .in2(N__23781),
            .in3(N__23774),
            .lcout(cmd_rdadctmp_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56093),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i5_LC_7_18_6 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i5_LC_7_18_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i5_LC_7_18_6 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i5_LC_7_18_6  (
            .in0(N__23765),
            .in1(N__29327),
            .in2(N__23778),
            .in3(N__38400),
            .lcout(cmd_rdadctmp_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56093),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i30_4_lut_LC_7_18_7 .C_ON=1'b0;
    defparam \ADC_IAC.i30_4_lut_LC_7_18_7 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i30_4_lut_LC_7_18_7 .LUT_INIT=16'b1100100001010001;
    LogicCell40 \ADC_IAC.i30_4_lut_LC_7_18_7  (
            .in0(N__24926),
            .in1(N__24851),
            .in2(N__24623),
            .in3(N__28708),
            .lcout(\ADC_IAC.n17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pll_main.i19991_1_lut_LC_8_1_5 .C_ON=1'b0;
    defparam \pll_main.i19991_1_lut_LC_8_1_5 .SEQ_MODE=4'b0000;
    defparam \pll_main.i19991_1_lut_LC_8_1_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \pll_main.i19991_1_lut_LC_8_1_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50810),
            .lcout(DDS_MCLK1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i18_LC_8_4_4 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i18_LC_8_4_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i18_LC_8_4_4 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \ADC_VDC.ADC_DATA_i18_LC_8_4_4  (
            .in0(N__51476),
            .in1(N__31620),
            .in2(N__24155),
            .in3(N__24198),
            .lcout(buf_adcdata_vdc_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42413),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i16_LC_8_5_0 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i16_LC_8_5_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i16_LC_8_5_0 .LUT_INIT=16'b0100111001000100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i16_LC_8_5_0  (
            .in0(N__29082),
            .in1(N__24029),
            .in2(N__51758),
            .in3(N__25469),
            .lcout(cmd_rdadctmp_16_adj_1507),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42365),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i17_LC_8_5_1 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i17_LC_8_5_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i17_LC_8_5_1 .LUT_INIT=16'b0011101100001000;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i17_LC_8_5_1  (
            .in0(N__24028),
            .in1(N__29084),
            .in2(N__51708),
            .in3(N__24004),
            .lcout(cmd_rdadctmp_17_adj_1506),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42365),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i19_LC_8_5_2 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i19_LC_8_5_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i19_LC_8_5_2 .LUT_INIT=16'b0010111100100000;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i19_LC_8_5_2  (
            .in0(N__23974),
            .in1(N__51640),
            .in2(N__29117),
            .in3(N__25258),
            .lcout(cmd_rdadctmp_19_adj_1504),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42365),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i6_LC_8_5_3 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i6_LC_8_5_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i6_LC_8_5_3 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i6_LC_8_5_3  (
            .in0(N__51639),
            .in1(N__25301),
            .in2(N__23909),
            .in3(N__29093),
            .lcout(cmd_rdadctmp_6_adj_1517),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42365),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i1_LC_8_5_4 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i1_LC_8_5_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i1_LC_8_5_4 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i1_LC_8_5_4  (
            .in0(N__29083),
            .in1(N__23831),
            .in2(N__25074),
            .in3(N__51648),
            .lcout(cmd_rdadctmp_1_adj_1522),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42365),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i0_LC_8_5_5 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i0_LC_8_5_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i0_LC_8_5_5 .LUT_INIT=16'b0000110010101010;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i0_LC_8_5_5  (
            .in0(N__23830),
            .in1(N__51942),
            .in2(N__51707),
            .in3(N__29091),
            .lcout(cmd_rdadctmp_0_adj_1523),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42365),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i7_LC_8_5_6 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i7_LC_8_5_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i7_LC_8_5_6 .LUT_INIT=16'b0010111100100000;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i7_LC_8_5_6  (
            .in0(N__23902),
            .in1(N__51641),
            .in2(N__29118),
            .in3(N__25277),
            .lcout(cmd_rdadctmp_7_adj_1516),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42365),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i18_LC_8_5_7 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i18_LC_8_5_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i18_LC_8_5_7 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i18_LC_8_5_7  (
            .in0(N__51638),
            .in1(N__24005),
            .in2(N__23981),
            .in3(N__29092),
            .lcout(cmd_rdadctmp_18_adj_1505),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42365),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadcbuf_i0_LC_8_6_0 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i0_LC_8_6_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i0_LC_8_6_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i0_LC_8_6_0  (
            .in0(_gnd_net_),
            .in1(N__23814),
            .in2(N__23835),
            .in3(_gnd_net_),
            .lcout(\ADC_VDC.cmd_rdadcbuf_0 ),
            .ltout(),
            .carryin(bfn_8_6_0_),
            .carryout(\ADC_VDC.n19842 ),
            .clk(N__42394),
            .ce(N__26908),
            .sr(N__26856));
    defparam \ADC_VDC.cmd_rdadcbuf_i1_LC_8_6_1 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i1_LC_8_6_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i1_LC_8_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i1_LC_8_6_1  (
            .in0(_gnd_net_),
            .in1(N__23808),
            .in2(N__25072),
            .in3(N__23802),
            .lcout(\ADC_VDC.cmd_rdadcbuf_1 ),
            .ltout(),
            .carryin(\ADC_VDC.n19842 ),
            .carryout(\ADC_VDC.n19843 ),
            .clk(N__42394),
            .ce(N__26908),
            .sr(N__26856));
    defparam \ADC_VDC.cmd_rdadcbuf_i2_LC_8_6_2 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i2_LC_8_6_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i2_LC_8_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i2_LC_8_6_2  (
            .in0(_gnd_net_),
            .in1(N__23952),
            .in2(N__25047),
            .in3(N__23946),
            .lcout(\ADC_VDC.cmd_rdadcbuf_2 ),
            .ltout(),
            .carryin(\ADC_VDC.n19843 ),
            .carryout(\ADC_VDC.n19844 ),
            .clk(N__42394),
            .ce(N__26908),
            .sr(N__26856));
    defparam \ADC_VDC.cmd_rdadcbuf_i3_LC_8_6_3 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i3_LC_8_6_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i3_LC_8_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i3_LC_8_6_3  (
            .in0(_gnd_net_),
            .in1(N__23943),
            .in2(N__25029),
            .in3(N__23937),
            .lcout(\ADC_VDC.cmd_rdadcbuf_3 ),
            .ltout(),
            .carryin(\ADC_VDC.n19844 ),
            .carryout(\ADC_VDC.n19845 ),
            .clk(N__42394),
            .ce(N__26908),
            .sr(N__26856));
    defparam \ADC_VDC.cmd_rdadcbuf_i4_LC_8_6_4 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i4_LC_8_6_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i4_LC_8_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i4_LC_8_6_4  (
            .in0(_gnd_net_),
            .in1(N__25315),
            .in2(N__23934),
            .in3(N__23922),
            .lcout(\ADC_VDC.cmd_rdadcbuf_4 ),
            .ltout(),
            .carryin(\ADC_VDC.n19845 ),
            .carryout(\ADC_VDC.n19846 ),
            .clk(N__42394),
            .ce(N__26908),
            .sr(N__26856));
    defparam \ADC_VDC.cmd_rdadcbuf_i5_LC_8_6_5 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i5_LC_8_6_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i5_LC_8_6_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i5_LC_8_6_5  (
            .in0(_gnd_net_),
            .in1(N__23919),
            .in2(N__25302),
            .in3(N__23913),
            .lcout(\ADC_VDC.cmd_rdadcbuf_5 ),
            .ltout(),
            .carryin(\ADC_VDC.n19846 ),
            .carryout(\ADC_VDC.n19847 ),
            .clk(N__42394),
            .ce(N__26908),
            .sr(N__26856));
    defparam \ADC_VDC.cmd_rdadcbuf_i6_LC_8_6_6 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i6_LC_8_6_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i6_LC_8_6_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i6_LC_8_6_6  (
            .in0(_gnd_net_),
            .in1(N__23883),
            .in2(N__23910),
            .in3(N__23877),
            .lcout(\ADC_VDC.cmd_rdadcbuf_6 ),
            .ltout(),
            .carryin(\ADC_VDC.n19847 ),
            .carryout(\ADC_VDC.n19848 ),
            .clk(N__42394),
            .ce(N__26908),
            .sr(N__26856));
    defparam \ADC_VDC.cmd_rdadcbuf_i7_LC_8_6_7 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i7_LC_8_6_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i7_LC_8_6_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i7_LC_8_6_7  (
            .in0(_gnd_net_),
            .in1(N__25276),
            .in2(N__23874),
            .in3(N__23865),
            .lcout(\ADC_VDC.cmd_rdadcbuf_7 ),
            .ltout(),
            .carryin(\ADC_VDC.n19848 ),
            .carryout(\ADC_VDC.n19849 ),
            .clk(N__42394),
            .ce(N__26908),
            .sr(N__26856));
    defparam \ADC_VDC.cmd_rdadcbuf_i8_LC_8_7_0 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i8_LC_8_7_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i8_LC_8_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i8_LC_8_7_0  (
            .in0(_gnd_net_),
            .in1(N__23862),
            .in2(N__25238),
            .in3(N__23856),
            .lcout(\ADC_VDC.cmd_rdadcbuf_8 ),
            .ltout(),
            .carryin(bfn_8_7_0_),
            .carryout(\ADC_VDC.n19850 ),
            .clk(N__42411),
            .ce(N__26946),
            .sr(N__26853));
    defparam \ADC_VDC.cmd_rdadcbuf_i9_LC_8_7_1 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i9_LC_8_7_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i9_LC_8_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i9_LC_8_7_1  (
            .in0(_gnd_net_),
            .in1(N__23853),
            .in2(N__25215),
            .in3(N__23847),
            .lcout(\ADC_VDC.cmd_rdadcbuf_9 ),
            .ltout(),
            .carryin(\ADC_VDC.n19850 ),
            .carryout(\ADC_VDC.n19851 ),
            .clk(N__42411),
            .ce(N__26946),
            .sr(N__26853));
    defparam \ADC_VDC.cmd_rdadcbuf_i10_LC_8_7_2 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i10_LC_8_7_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i10_LC_8_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i10_LC_8_7_2  (
            .in0(_gnd_net_),
            .in1(N__23844),
            .in2(N__25194),
            .in3(N__23838),
            .lcout(\ADC_VDC.cmd_rdadcbuf_10 ),
            .ltout(),
            .carryin(\ADC_VDC.n19851 ),
            .carryout(\ADC_VDC.n19852 ),
            .clk(N__42411),
            .ce(N__26946),
            .sr(N__26853));
    defparam \ADC_VDC.cmd_rdadcbuf_i11_LC_8_7_3 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i11_LC_8_7_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i11_LC_8_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i11_LC_8_7_3  (
            .in0(_gnd_net_),
            .in1(N__25379),
            .in2(N__25167),
            .in3(N__24066),
            .lcout(cmd_rdadcbuf_11),
            .ltout(),
            .carryin(\ADC_VDC.n19852 ),
            .carryout(\ADC_VDC.n19853 ),
            .clk(N__42411),
            .ce(N__26946),
            .sr(N__26853));
    defparam \ADC_VDC.cmd_rdadcbuf_i12_LC_8_7_4 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i12_LC_8_7_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i12_LC_8_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i12_LC_8_7_4  (
            .in0(_gnd_net_),
            .in1(N__25147),
            .in2(N__31493),
            .in3(N__24063),
            .lcout(cmd_rdadcbuf_12),
            .ltout(),
            .carryin(\ADC_VDC.n19853 ),
            .carryout(\ADC_VDC.n19854 ),
            .clk(N__42411),
            .ce(N__26946),
            .sr(N__26853));
    defparam \ADC_VDC.cmd_rdadcbuf_i13_LC_8_7_5 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i13_LC_8_7_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i13_LC_8_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i13_LC_8_7_5  (
            .in0(_gnd_net_),
            .in1(N__25658),
            .in2(N__25126),
            .in3(N__24060),
            .lcout(cmd_rdadcbuf_13),
            .ltout(),
            .carryin(\ADC_VDC.n19854 ),
            .carryout(\ADC_VDC.n19855 ),
            .clk(N__42411),
            .ce(N__26946),
            .sr(N__26853));
    defparam \ADC_VDC.cmd_rdadcbuf_i14_LC_8_7_6 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i14_LC_8_7_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i14_LC_8_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i14_LC_8_7_6  (
            .in0(_gnd_net_),
            .in1(N__24050),
            .in2(N__25488),
            .in3(N__24039),
            .lcout(cmd_rdadcbuf_14),
            .ltout(),
            .carryin(\ADC_VDC.n19855 ),
            .carryout(\ADC_VDC.n19856 ),
            .clk(N__42411),
            .ce(N__26946),
            .sr(N__26853));
    defparam \ADC_VDC.cmd_rdadcbuf_i15_LC_8_7_7 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i15_LC_8_7_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i15_LC_8_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i15_LC_8_7_7  (
            .in0(_gnd_net_),
            .in1(N__25619),
            .in2(N__25470),
            .in3(N__24036),
            .lcout(cmd_rdadcbuf_15),
            .ltout(),
            .carryin(\ADC_VDC.n19856 ),
            .carryout(\ADC_VDC.n19857 ),
            .clk(N__42411),
            .ce(N__26946),
            .sr(N__26853));
    defparam \ADC_VDC.cmd_rdadcbuf_i16_LC_8_8_0 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i16_LC_8_8_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i16_LC_8_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i16_LC_8_8_0  (
            .in0(_gnd_net_),
            .in1(N__25586),
            .in2(N__24033),
            .in3(N__24012),
            .lcout(cmd_rdadcbuf_16),
            .ltout(),
            .carryin(bfn_8_8_0_),
            .carryout(\ADC_VDC.n19858 ),
            .clk(N__42384),
            .ce(N__26930),
            .sr(N__26854));
    defparam \ADC_VDC.cmd_rdadcbuf_i17_LC_8_8_1 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i17_LC_8_8_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i17_LC_8_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i17_LC_8_8_1  (
            .in0(_gnd_net_),
            .in1(N__25419),
            .in2(N__24009),
            .in3(N__23988),
            .lcout(cmd_rdadcbuf_17),
            .ltout(),
            .carryin(\ADC_VDC.n19858 ),
            .carryout(\ADC_VDC.n19859 ),
            .clk(N__42384),
            .ce(N__26930),
            .sr(N__26854));
    defparam \ADC_VDC.cmd_rdadcbuf_i18_LC_8_8_2 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i18_LC_8_8_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i18_LC_8_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i18_LC_8_8_2  (
            .in0(_gnd_net_),
            .in1(N__26777),
            .in2(N__23985),
            .in3(N__23955),
            .lcout(cmd_rdadcbuf_18),
            .ltout(),
            .carryin(\ADC_VDC.n19859 ),
            .carryout(\ADC_VDC.n19860 ),
            .clk(N__42384),
            .ce(N__26930),
            .sr(N__26854));
    defparam \ADC_VDC.cmd_rdadcbuf_i19_LC_8_8_3 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i19_LC_8_8_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i19_LC_8_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i19_LC_8_8_3  (
            .in0(_gnd_net_),
            .in1(N__25260),
            .in2(N__29666),
            .in3(N__24093),
            .lcout(cmd_rdadcbuf_19),
            .ltout(),
            .carryin(\ADC_VDC.n19860 ),
            .carryout(\ADC_VDC.n19861 ),
            .clk(N__42384),
            .ce(N__26930),
            .sr(N__26854));
    defparam \ADC_VDC.cmd_rdadcbuf_i20_LC_8_8_4 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i20_LC_8_8_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i20_LC_8_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i20_LC_8_8_4  (
            .in0(_gnd_net_),
            .in1(N__25448),
            .in2(N__25554),
            .in3(N__24090),
            .lcout(cmd_rdadcbuf_20),
            .ltout(),
            .carryin(\ADC_VDC.n19861 ),
            .carryout(\ADC_VDC.n19862 ),
            .clk(N__42384),
            .ce(N__26930),
            .sr(N__26854));
    defparam \ADC_VDC.cmd_rdadcbuf_i21_LC_8_8_5 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i21_LC_8_8_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i21_LC_8_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i21_LC_8_8_5  (
            .in0(_gnd_net_),
            .in1(N__25343),
            .in2(N__25529),
            .in3(N__24087),
            .lcout(cmd_rdadcbuf_21),
            .ltout(),
            .carryin(\ADC_VDC.n19862 ),
            .carryout(\ADC_VDC.n19863 ),
            .clk(N__42384),
            .ce(N__26930),
            .sr(N__26854));
    defparam \ADC_VDC.cmd_rdadcbuf_i22_LC_8_8_6 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i22_LC_8_8_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i22_LC_8_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i22_LC_8_8_6  (
            .in0(_gnd_net_),
            .in1(N__26705),
            .in2(N__30279),
            .in3(N__24084),
            .lcout(cmd_rdadcbuf_22),
            .ltout(),
            .carryin(\ADC_VDC.n19863 ),
            .carryout(\ADC_VDC.n19864 ),
            .clk(N__42384),
            .ce(N__26930),
            .sr(N__26854));
    defparam \ADC_VDC.cmd_rdadcbuf_i23_LC_8_8_7 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i23_LC_8_8_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i23_LC_8_8_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i23_LC_8_8_7  (
            .in0(_gnd_net_),
            .in1(N__26792),
            .in2(N__30243),
            .in3(N__24081),
            .lcout(cmd_rdadcbuf_23),
            .ltout(),
            .carryin(\ADC_VDC.n19864 ),
            .carryout(\ADC_VDC.n19865 ),
            .clk(N__42384),
            .ce(N__26930),
            .sr(N__26854));
    defparam \ADC_VDC.cmd_rdadcbuf_i24_LC_8_9_0 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i24_LC_8_9_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i24_LC_8_9_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i24_LC_8_9_0  (
            .in0(_gnd_net_),
            .in1(N__29642),
            .in2(_gnd_net_),
            .in3(N__24078),
            .lcout(cmd_rdadcbuf_24),
            .ltout(),
            .carryin(bfn_8_9_0_),
            .carryout(\ADC_VDC.n19866 ),
            .clk(N__42412),
            .ce(N__26941),
            .sr(N__26868));
    defparam \ADC_VDC.cmd_rdadcbuf_i25_LC_8_9_1 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i25_LC_8_9_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i25_LC_8_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i25_LC_8_9_1  (
            .in0(_gnd_net_),
            .in1(N__26720),
            .in2(_gnd_net_),
            .in3(N__24075),
            .lcout(cmd_rdadcbuf_25),
            .ltout(),
            .carryin(\ADC_VDC.n19866 ),
            .carryout(\ADC_VDC.n19867 ),
            .clk(N__42412),
            .ce(N__26941),
            .sr(N__26868));
    defparam \ADC_VDC.cmd_rdadcbuf_i26_LC_8_9_2 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i26_LC_8_9_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i26_LC_8_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i26_LC_8_9_2  (
            .in0(_gnd_net_),
            .in1(N__26738),
            .in2(_gnd_net_),
            .in3(N__24072),
            .lcout(cmd_rdadcbuf_26),
            .ltout(),
            .carryin(\ADC_VDC.n19867 ),
            .carryout(\ADC_VDC.n19868 ),
            .clk(N__42412),
            .ce(N__26941),
            .sr(N__26868));
    defparam \ADC_VDC.cmd_rdadcbuf_i27_LC_8_9_3 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i27_LC_8_9_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i27_LC_8_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i27_LC_8_9_3  (
            .in0(_gnd_net_),
            .in1(N__25100),
            .in2(_gnd_net_),
            .in3(N__24069),
            .lcout(cmd_rdadcbuf_27),
            .ltout(),
            .carryin(\ADC_VDC.n19868 ),
            .carryout(\ADC_VDC.n19869 ),
            .clk(N__42412),
            .ce(N__26941),
            .sr(N__26868));
    defparam \ADC_VDC.cmd_rdadcbuf_i28_LC_8_9_4 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i28_LC_8_9_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i28_LC_8_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i28_LC_8_9_4  (
            .in0(_gnd_net_),
            .in1(N__29564),
            .in2(_gnd_net_),
            .in3(N__24201),
            .lcout(cmd_rdadcbuf_28),
            .ltout(),
            .carryin(\ADC_VDC.n19869 ),
            .carryout(\ADC_VDC.n19870 ),
            .clk(N__42412),
            .ce(N__26941),
            .sr(N__26868));
    defparam \ADC_VDC.cmd_rdadcbuf_i29_LC_8_9_5 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i29_LC_8_9_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i29_LC_8_9_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i29_LC_8_9_5  (
            .in0(_gnd_net_),
            .in1(N__24191),
            .in2(_gnd_net_),
            .in3(N__24180),
            .lcout(cmd_rdadcbuf_29),
            .ltout(),
            .carryin(\ADC_VDC.n19870 ),
            .carryout(\ADC_VDC.n19871 ),
            .clk(N__42412),
            .ce(N__26941),
            .sr(N__26868));
    defparam \ADC_VDC.cmd_rdadcbuf_i30_LC_8_9_6 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i30_LC_8_9_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i30_LC_8_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i30_LC_8_9_6  (
            .in0(_gnd_net_),
            .in1(N__29600),
            .in2(_gnd_net_),
            .in3(N__24177),
            .lcout(cmd_rdadcbuf_30),
            .ltout(),
            .carryin(\ADC_VDC.n19871 ),
            .carryout(\ADC_VDC.n19872 ),
            .clk(N__42412),
            .ce(N__26941),
            .sr(N__26868));
    defparam \ADC_VDC.cmd_rdadcbuf_i31_LC_8_9_7 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i31_LC_8_9_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i31_LC_8_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i31_LC_8_9_7  (
            .in0(_gnd_net_),
            .in1(N__29474),
            .in2(_gnd_net_),
            .in3(N__24174),
            .lcout(cmd_rdadcbuf_31),
            .ltout(),
            .carryin(\ADC_VDC.n19872 ),
            .carryout(\ADC_VDC.n19873 ),
            .clk(N__42412),
            .ce(N__26941),
            .sr(N__26868));
    defparam \ADC_VDC.cmd_rdadcbuf_i32_LC_8_10_0 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i32_LC_8_10_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i32_LC_8_10_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i32_LC_8_10_0  (
            .in0(_gnd_net_),
            .in1(N__29519),
            .in2(_gnd_net_),
            .in3(N__24171),
            .lcout(cmd_rdadcbuf_32),
            .ltout(),
            .carryin(bfn_8_10_0_),
            .carryout(\ADC_VDC.n19874 ),
            .clk(N__42434),
            .ce(N__26945),
            .sr(N__26855));
    defparam \ADC_VDC.cmd_rdadcbuf_i33_LC_8_10_1 .C_ON=1'b1;
    defparam \ADC_VDC.cmd_rdadcbuf_i33_LC_8_10_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i33_LC_8_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i33_LC_8_10_1  (
            .in0(_gnd_net_),
            .in1(N__25328),
            .in2(_gnd_net_),
            .in3(N__24168),
            .lcout(cmd_rdadcbuf_33),
            .ltout(),
            .carryin(\ADC_VDC.n19874 ),
            .carryout(\ADC_VDC.n19875 ),
            .clk(N__42434),
            .ce(N__26945),
            .sr(N__26855));
    defparam \ADC_VDC.add_23_36_lut_LC_8_10_2 .C_ON=1'b0;
    defparam \ADC_VDC.add_23_36_lut_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.add_23_36_lut_LC_8_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.add_23_36_lut_LC_8_10_2  (
            .in0(_gnd_net_),
            .in1(N__25861),
            .in2(_gnd_net_),
            .in3(N__24165),
            .lcout(\ADC_VDC.cmd_rdadcbuf_35_N_1296_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_2_i19_3_lut_LC_8_11_0.C_ON=1'b0;
    defparam mux_128_Mux_2_i19_3_lut_LC_8_11_0.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_2_i19_3_lut_LC_8_11_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_128_Mux_2_i19_3_lut_LC_8_11_0 (
            .in0(N__57148),
            .in1(N__24162),
            .in2(_gnd_net_),
            .in3(N__24131),
            .lcout(n19_adj_1683),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_1_i19_3_lut_LC_8_11_1.C_ON=1'b0;
    defparam mux_128_Mux_1_i19_3_lut_LC_8_11_1.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_1_i19_3_lut_LC_8_11_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_128_Mux_1_i19_3_lut_LC_8_11_1 (
            .in0(N__29553),
            .in1(N__24521),
            .in2(_gnd_net_),
            .in3(N__57149),
            .lcout(n19_adj_1692),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i5_LC_8_11_2 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i5_LC_8_11_2 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i5_LC_8_11_2 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \ADC_IAC.ADC_DATA_i5_LC_8_11_2  (
            .in0(N__24227),
            .in1(N__24357),
            .in2(N__38607),
            .in3(N__38775),
            .lcout(buf_adcdata_iac_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55988),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i2_LC_8_11_3 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i2_LC_8_11_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i2_LC_8_11_3 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_IAC.ADC_DATA_i2_LC_8_11_3  (
            .in0(N__38774),
            .in1(N__38602),
            .in2(N__24290),
            .in3(N__24330),
            .lcout(buf_adcdata_iac_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55988),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_5_i19_3_lut_LC_8_11_4.C_ON=1'b0;
    defparam mux_130_Mux_5_i19_3_lut_LC_8_11_4.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_5_i19_3_lut_LC_8_11_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_130_Mux_5_i19_3_lut_LC_8_11_4 (
            .in0(N__57150),
            .in1(N__25575),
            .in2(_gnd_net_),
            .in3(N__24253),
            .lcout(),
            .ltout(n19_adj_1603_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_5_i22_3_lut_LC_8_11_5.C_ON=1'b0;
    defparam mux_130_Mux_5_i22_3_lut_LC_8_11_5.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_5_i22_3_lut_LC_8_11_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 mux_130_Mux_5_i22_3_lut_LC_8_11_5 (
            .in0(_gnd_net_),
            .in1(N__24226),
            .in2(N__24213),
            .in3(N__47453),
            .lcout(n22_adj_1604),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i20_LC_8_11_6 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i20_LC_8_11_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i20_LC_8_11_6 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i20_LC_8_11_6  (
            .in0(N__27500),
            .in1(N__27458),
            .in2(N__27858),
            .in3(N__28269),
            .lcout(cmd_rdadctmp_20_adj_1472),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55988),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i2_LC_8_11_7.C_ON=1'b0;
    defparam comm_cmd_i2_LC_8_11_7.SEQ_MODE=4'b1000;
    defparam comm_cmd_i2_LC_8_11_7.LUT_INIT=16'b1011100000110000;
    LogicCell40 comm_cmd_i2_LC_8_11_7 (
            .in0(N__50994),
            .in1(N__37532),
            .in2(N__47537),
            .in3(N__50157),
            .lcout(comm_cmd_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55988),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.dds_state_i0_LC_8_12_1 .C_ON=1'b0;
    defparam \SIG_DDS.dds_state_i0_LC_8_12_1 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.dds_state_i0_LC_8_12_1 .LUT_INIT=16'b1010000000110011;
    LogicCell40 \SIG_DDS.dds_state_i0_LC_8_12_1  (
            .in0(N__36591),
            .in1(N__44702),
            .in2(N__24453),
            .in3(N__44516),
            .lcout(dds_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56001),
            .ce(N__44550),
            .sr(_gnd_net_));
    defparam comm_cmd_2__bdd_4_lut_19668_LC_8_12_3.C_ON=1'b0;
    defparam comm_cmd_2__bdd_4_lut_19668_LC_8_12_3.SEQ_MODE=4'b0000;
    defparam comm_cmd_2__bdd_4_lut_19668_LC_8_12_3.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_2__bdd_4_lut_19668_LC_8_12_3 (
            .in0(N__30558),
            .in1(N__47190),
            .in2(N__32580),
            .in3(N__47457),
            .lcout(),
            .ltout(n22377_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22377_bdd_4_lut_LC_8_12_4.C_ON=1'b0;
    defparam n22377_bdd_4_lut_LC_8_12_4.SEQ_MODE=4'b0000;
    defparam n22377_bdd_4_lut_LC_8_12_4.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22377_bdd_4_lut_LC_8_12_4 (
            .in0(N__47191),
            .in1(N__30735),
            .in2(N__24210),
            .in3(N__24207),
            .lcout(n22380),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i1_LC_8_13_0.C_ON=1'b0;
    defparam comm_buf_6__i1_LC_8_13_0.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i1_LC_8_13_0.LUT_INIT=16'b0011000010101010;
    LogicCell40 comm_buf_6__i1_LC_8_13_0 (
            .in0(N__49973),
            .in1(N__55461),
            .in2(N__49746),
            .in3(N__53141),
            .lcout(comm_buf_6_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56018),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i13_LC_8_13_2.C_ON=1'b0;
    defparam buf_dds1_i13_LC_8_13_2.SEQ_MODE=4'b1000;
    defparam buf_dds1_i13_LC_8_13_2.LUT_INIT=16'b1011100011111100;
    LogicCell40 buf_dds1_i13_LC_8_13_2 (
            .in0(N__30723),
            .in1(N__46916),
            .in2(N__34967),
            .in3(N__55462),
            .lcout(buf_dds1_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56018),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i5_LC_8_13_3.C_ON=1'b0;
    defparam buf_dds1_i5_LC_8_13_3.SEQ_MODE=4'b1000;
    defparam buf_dds1_i5_LC_8_13_3.LUT_INIT=16'b1111010111001100;
    LogicCell40 buf_dds1_i5_LC_8_13_3 (
            .in0(N__55460),
            .in1(N__25364),
            .in2(N__37257),
            .in3(N__46915),
            .lcout(buf_dds1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56018),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i10_LC_8_13_4 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i10_LC_8_13_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i10_LC_8_13_4 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC.ADC_DATA_i10_LC_8_13_4  (
            .in0(N__27966),
            .in1(N__27827),
            .in2(N__27325),
            .in3(N__26122),
            .lcout(buf_adcdata_vac_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56018),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i20_LC_8_13_5 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i20_LC_8_13_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i20_LC_8_13_5 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i20_LC_8_13_5  (
            .in0(N__27826),
            .in1(N__27967),
            .in2(N__24417),
            .in3(N__31859),
            .lcout(buf_adcdata_vac_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56018),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i14_LC_8_13_6 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i14_LC_8_13_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i14_LC_8_13_6 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \ADC_IAC.ADC_DATA_i14_LC_8_13_6  (
            .in0(N__38750),
            .in1(N__43378),
            .in2(N__24669),
            .in3(N__38606),
            .lcout(buf_adcdata_iac_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56018),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i0_LC_8_14_0 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i0_LC_8_14_0 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i0_LC_8_14_0 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \CLK_DDS.tmp_buf_i0_LC_8_14_0  (
            .in0(N__29873),
            .in1(N__30108),
            .in2(N__41736),
            .in3(N__24392),
            .lcout(\CLK_DDS.tmp_buf_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56032),
            .ce(N__30143),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i1_LC_8_14_1 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i1_LC_8_14_1 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i1_LC_8_14_1 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \CLK_DDS.tmp_buf_i1_LC_8_14_1  (
            .in0(N__30104),
            .in1(N__29874),
            .in2(N__24381),
            .in3(N__35607),
            .lcout(\CLK_DDS.tmp_buf_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56032),
            .ce(N__30143),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i2_LC_8_14_2 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i2_LC_8_14_2 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i2_LC_8_14_2 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \CLK_DDS.tmp_buf_i2_LC_8_14_2  (
            .in0(N__29875),
            .in1(N__24372),
            .in2(N__30114),
            .in3(N__26265),
            .lcout(\CLK_DDS.tmp_buf_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56032),
            .ce(N__30143),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i3_LC_8_14_3 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i3_LC_8_14_3 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i3_LC_8_14_3 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \CLK_DDS.tmp_buf_i3_LC_8_14_3  (
            .in0(N__30105),
            .in1(N__29876),
            .in2(N__24366),
            .in3(N__32688),
            .lcout(\CLK_DDS.tmp_buf_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56032),
            .ce(N__30143),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i4_LC_8_14_4 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i4_LC_8_14_4 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i4_LC_8_14_4 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLK_DDS.tmp_buf_i4_LC_8_14_4  (
            .in0(N__29877),
            .in1(N__30109),
            .in2(N__24576),
            .in3(N__29456),
            .lcout(\CLK_DDS.tmp_buf_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56032),
            .ce(N__30143),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i5_LC_8_14_5 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i5_LC_8_14_5 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i5_LC_8_14_5 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \CLK_DDS.tmp_buf_i5_LC_8_14_5  (
            .in0(N__30106),
            .in1(N__29878),
            .in2(N__24567),
            .in3(N__25363),
            .lcout(\CLK_DDS.tmp_buf_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56032),
            .ce(N__30143),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i6_LC_8_14_6 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i6_LC_8_14_6 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i6_LC_8_14_6 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \CLK_DDS.tmp_buf_i6_LC_8_14_6  (
            .in0(N__29879),
            .in1(N__30110),
            .in2(N__24558),
            .in3(N__46965),
            .lcout(\CLK_DDS.tmp_buf_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56032),
            .ce(N__30143),
            .sr(_gnd_net_));
    defparam \CLK_DDS.tmp_buf_i7_LC_8_14_7 .C_ON=1'b0;
    defparam \CLK_DDS.tmp_buf_i7_LC_8_14_7 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.tmp_buf_i7_LC_8_14_7 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \CLK_DDS.tmp_buf_i7_LC_8_14_7  (
            .in0(N__30107),
            .in1(N__29880),
            .in2(N__24549),
            .in3(N__36576),
            .lcout(\CLK_DDS.tmp_buf_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56032),
            .ce(N__30143),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i17_LC_8_15_0 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i17_LC_8_15_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i17_LC_8_15_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i17_LC_8_15_0  (
            .in0(N__27978),
            .in1(N__27824),
            .in2(N__26208),
            .in3(N__24520),
            .lcout(buf_adcdata_vac_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56048),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.i4_4_lut_LC_8_15_1 .C_ON=1'b0;
    defparam \SIG_DDS.i4_4_lut_LC_8_15_1 .SEQ_MODE=4'b0000;
    defparam \SIG_DDS.i4_4_lut_LC_8_15_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \SIG_DDS.i4_4_lut_LC_8_15_1  (
            .in0(N__24492),
            .in1(N__24437),
            .in2(N__24472),
            .in3(N__44709),
            .lcout(\SIG_DDS.n10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.bit_cnt_i0_LC_8_15_2 .C_ON=1'b0;
    defparam \SIG_DDS.bit_cnt_i0_LC_8_15_2 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.bit_cnt_i0_LC_8_15_2 .LUT_INIT=16'b0000010100001010;
    LogicCell40 \SIG_DDS.bit_cnt_i0_LC_8_15_2  (
            .in0(N__44508),
            .in1(_gnd_net_),
            .in2(N__24641),
            .in3(N__24438),
            .lcout(bit_cnt_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56048),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i8_LC_8_15_3.C_ON=1'b0;
    defparam buf_dds1_i8_LC_8_15_3.SEQ_MODE=4'b1000;
    defparam buf_dds1_i8_LC_8_15_3.LUT_INIT=16'b1110001000000000;
    LogicCell40 buf_dds1_i8_LC_8_15_3 (
            .in0(N__39104),
            .in1(N__46914),
            .in2(N__45647),
            .in3(N__46754),
            .lcout(buf_dds1_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56048),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i22_LC_8_15_4 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i22_LC_8_15_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i22_LC_8_15_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i22_LC_8_15_4  (
            .in0(N__28089),
            .in1(N__27825),
            .in2(N__26347),
            .in3(N__28237),
            .lcout(cmd_rdadctmp_22_adj_1470),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56048),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_adj_292_LC_8_15_6.C_ON=1'b0;
    defparam i2_3_lut_adj_292_LC_8_15_6.SEQ_MODE=4'b0000;
    defparam i2_3_lut_adj_292_LC_8_15_6.LUT_INIT=16'b0000000001000100;
    LogicCell40 i2_3_lut_adj_292_LC_8_15_6 (
            .in0(N__46454),
            .in1(N__47193),
            .in2(_gnd_net_),
            .in3(N__47532),
            .lcout(n69),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i5_LC_8_16_1 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i5_LC_8_16_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i5_LC_8_16_1 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i5_LC_8_16_1  (
            .in0(N__24698),
            .in1(N__24720),
            .in2(N__27855),
            .in3(N__28185),
            .lcout(cmd_rdadctmp_5_adj_1487),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56062),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i22_LC_8_16_2 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i22_LC_8_16_2 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i22_LC_8_16_2 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i22_LC_8_16_2  (
            .in0(N__24658),
            .in1(N__29386),
            .in2(N__33114),
            .in3(N__38456),
            .lcout(cmd_rdadctmp_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56062),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i6_LC_8_16_3 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i6_LC_8_16_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i6_LC_8_16_3 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i6_LC_8_16_3  (
            .in0(N__24680),
            .in1(N__27778),
            .in2(N__24702),
            .in3(N__28186),
            .lcout(cmd_rdadctmp_6_adj_1486),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56062),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i22_LC_8_16_4 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i22_LC_8_16_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i22_LC_8_16_4 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_IAC.ADC_DATA_i22_LC_8_16_4  (
            .in0(N__38640),
            .in1(N__38455),
            .in2(N__30778),
            .in3(N__26585),
            .lcout(buf_adcdata_iac_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56062),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i23_LC_8_16_5 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i23_LC_8_16_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i23_LC_8_16_5 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i23_LC_8_16_5  (
            .in0(N__38454),
            .in1(N__24659),
            .in2(N__29394),
            .in3(N__28738),
            .lcout(cmd_rdadctmp_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56062),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.i12572_3_lut_LC_8_16_6 .C_ON=1'b0;
    defparam \SIG_DDS.i12572_3_lut_LC_8_16_6 .SEQ_MODE=4'b0000;
    defparam \SIG_DDS.i12572_3_lut_LC_8_16_6 .LUT_INIT=16'b1011101100000000;
    LogicCell40 \SIG_DDS.i12572_3_lut_LC_8_16_6  (
            .in0(N__44667),
            .in1(N__44708),
            .in2(_gnd_net_),
            .in3(N__44504),
            .lcout(n15092),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i28_LC_8_17_2 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i28_LC_8_17_2 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i28_LC_8_17_2 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i28_LC_8_17_2  (
            .in0(N__38403),
            .in1(N__28900),
            .in2(N__26408),
            .in3(N__29325),
            .lcout(cmd_rdadctmp_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56076),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i29_LC_8_17_3 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i29_LC_8_17_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i29_LC_8_17_3 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i29_LC_8_17_3  (
            .in0(N__29323),
            .in1(N__28960),
            .in2(N__28907),
            .in3(N__38404),
            .lcout(cmd_rdadctmp_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56076),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i1_4_lut_adj_3_LC_8_17_5 .C_ON=1'b0;
    defparam \ADC_IAC.i1_4_lut_adj_3_LC_8_17_5 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i1_4_lut_adj_3_LC_8_17_5 .LUT_INIT=16'b1100110111101111;
    LogicCell40 \ADC_IAC.i1_4_lut_adj_3_LC_8_17_5  (
            .in0(N__24903),
            .in1(N__38402),
            .in2(N__24624),
            .in3(N__28709),
            .lcout(),
            .ltout(\ADC_IAC.n21159_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.i1_2_lut_LC_8_17_6 .C_ON=1'b0;
    defparam \ADC_IAC.i1_2_lut_LC_8_17_6 .SEQ_MODE=4'b0000;
    defparam \ADC_IAC.i1_2_lut_LC_8_17_6 .LUT_INIT=16'b1111000011111111;
    LogicCell40 \ADC_IAC.i1_2_lut_LC_8_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25011),
            .in3(N__24842),
            .lcout(\ADC_IAC.n21160 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i30_LC_8_17_7 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i30_LC_8_17_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i30_LC_8_17_7 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i30_LC_8_17_7  (
            .in0(N__29324),
            .in1(N__38405),
            .in2(N__26586),
            .in3(N__28961),
            .lcout(cmd_rdadctmp_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56076),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i19_LC_8_18_0 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i19_LC_8_18_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i19_LC_8_18_0 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i19_LC_8_18_0  (
            .in0(N__38449),
            .in1(N__26383),
            .in2(N__38265),
            .in3(N__29334),
            .lcout(cmd_rdadctmp_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56086),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i1_LC_8_18_1 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i1_LC_8_18_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i1_LC_8_18_1 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i1_LC_8_18_1  (
            .in0(N__24998),
            .in1(N__29333),
            .in2(N__24954),
            .in3(N__38453),
            .lcout(cmd_rdadctmp_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56086),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i2_LC_8_18_2 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i2_LC_8_18_2 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i2_LC_8_18_2 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i2_LC_8_18_2  (
            .in0(N__38451),
            .in1(N__24999),
            .in2(N__24990),
            .in3(N__29336),
            .lcout(cmd_rdadctmp_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56086),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i0_LC_8_18_3 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i0_LC_8_18_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i0_LC_8_18_3 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i0_LC_8_18_3  (
            .in0(N__24950),
            .in1(N__29332),
            .in2(N__24975),
            .in3(N__38452),
            .lcout(cmd_rdadctmp_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56086),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i20_LC_8_18_4 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i20_LC_8_18_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i20_LC_8_18_4 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i20_LC_8_18_4  (
            .in0(N__38450),
            .in1(N__26384),
            .in2(N__29429),
            .in3(N__29335),
            .lcout(cmd_rdadctmp_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56086),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.SCLK_35_LC_8_19_4 .C_ON=1'b0;
    defparam \ADC_IAC.SCLK_35_LC_8_19_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.SCLK_35_LC_8_19_4 .LUT_INIT=16'b1101000011100100;
    LogicCell40 \ADC_IAC.SCLK_35_LC_8_19_4  (
            .in0(N__38588),
            .in1(N__24941),
            .in2(N__24776),
            .in3(N__24855),
            .lcout(IAC_SCLK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56094),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i17_LC_8_19_5 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i17_LC_8_19_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i17_LC_8_19_5 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i17_LC_8_19_5  (
            .in0(N__38762),
            .in1(N__38589),
            .in2(N__28887),
            .in3(N__24742),
            .lcout(buf_adcdata_iac_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56094),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i16_LC_9_3_0 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i16_LC_9_3_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i16_LC_9_3_0 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \ADC_VDC.ADC_DATA_i16_LC_9_3_0  (
            .in0(N__51489),
            .in1(N__31625),
            .in2(N__25799),
            .in3(N__25107),
            .lcout(buf_adcdata_vdc_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42429),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i7791_3_lut_4_lut_LC_9_3_4 .C_ON=1'b0;
    defparam \ADC_VDC.i7791_3_lut_4_lut_LC_9_3_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i7791_3_lut_4_lut_LC_9_3_4 .LUT_INIT=16'b0101001011011010;
    LogicCell40 \ADC_VDC.i7791_3_lut_4_lut_LC_9_3_4  (
            .in0(N__51908),
            .in1(N__51174),
            .in2(N__52004),
            .in3(N__31661),
            .lcout(),
            .ltout(\ADC_VDC.n10309_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_4_lut_4_lut_adj_29_LC_9_3_5 .C_ON=1'b0;
    defparam \ADC_VDC.i1_4_lut_4_lut_adj_29_LC_9_3_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_4_lut_4_lut_adj_29_LC_9_3_5 .LUT_INIT=16'b1101110011111110;
    LogicCell40 \ADC_VDC.i1_4_lut_4_lut_adj_29_LC_9_3_5  (
            .in0(N__51637),
            .in1(N__51488),
            .in2(N__25089),
            .in3(N__29688),
            .lcout(\ADC_VDC.n13276 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.adc_state_i3_LC_9_4_3 .C_ON=1'b0;
    defparam \ADC_VDC.adc_state_i3_LC_9_4_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.adc_state_i3_LC_9_4_3 .LUT_INIT=16'b0001100000110000;
    LogicCell40 \ADC_VDC.adc_state_i3_LC_9_4_3  (
            .in0(N__51894),
            .in1(N__51500),
            .in2(N__51709),
            .in3(N__51179),
            .lcout(adc_state_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42399),
            .ce(N__25086),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i22_LC_9_5_0 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i22_LC_9_5_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i22_LC_9_5_0 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i22_LC_9_5_0  (
            .in0(N__51696),
            .in1(N__29080),
            .in2(N__30274),
            .in3(N__25530),
            .lcout(cmd_rdadctmp_22_adj_1501),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42301),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i10_LC_9_5_2 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i10_LC_9_5_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i10_LC_9_5_2 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i10_LC_9_5_2  (
            .in0(N__25213),
            .in1(N__29070),
            .in2(N__25193),
            .in3(N__51602),
            .lcout(cmd_rdadctmp_10_adj_1513),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42301),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i3_LC_9_5_3 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i3_LC_9_5_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i3_LC_9_5_3 .LUT_INIT=16'b0010111100100000;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i3_LC_9_5_3  (
            .in0(N__25046),
            .in1(N__51698),
            .in2(N__29114),
            .in3(N__25027),
            .lcout(cmd_rdadctmp_3_adj_1520),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42301),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i2_LC_9_5_4 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i2_LC_9_5_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i2_LC_9_5_4 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i2_LC_9_5_4  (
            .in0(N__51697),
            .in1(N__25045),
            .in2(N__25073),
            .in3(N__29081),
            .lcout(cmd_rdadctmp_2_adj_1521),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42301),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i4_LC_9_5_5 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i4_LC_9_5_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i4_LC_9_5_5 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i4_LC_9_5_5  (
            .in0(N__51600),
            .in1(N__25316),
            .in2(N__29115),
            .in3(N__25028),
            .lcout(cmd_rdadctmp_4_adj_1519),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42301),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_4_lut_4_lut_4_lut_LC_9_5_6 .C_ON=1'b0;
    defparam \ADC_VDC.i1_4_lut_4_lut_4_lut_LC_9_5_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_4_lut_4_lut_4_lut_LC_9_5_6 .LUT_INIT=16'b1010110010001000;
    LogicCell40 \ADC_VDC.i1_4_lut_4_lut_4_lut_LC_9_5_6  (
            .in0(N__51412),
            .in1(N__51599),
            .in2(N__51910),
            .in3(N__51145),
            .lcout(\ADC_VDC.n13463 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i5_LC_9_5_7 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i5_LC_9_5_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i5_LC_9_5_7 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i5_LC_9_5_7  (
            .in0(N__51601),
            .in1(N__25300),
            .in2(N__29116),
            .in3(N__25317),
            .lcout(cmd_rdadctmp_5_adj_1518),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42301),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i8_LC_9_6_0 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i8_LC_9_6_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i8_LC_9_6_0 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i8_LC_9_6_0  (
            .in0(N__51704),
            .in1(N__25234),
            .in2(N__25281),
            .in3(N__29136),
            .lcout(cmd_rdadctmp_8_adj_1515),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42424),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i20_LC_9_6_1 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i20_LC_9_6_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i20_LC_9_6_1 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i20_LC_9_6_1  (
            .in0(N__51701),
            .in1(N__25549),
            .in2(N__29142),
            .in3(N__25259),
            .lcout(cmd_rdadctmp_20_adj_1503),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42424),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i9_LC_9_6_2 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i9_LC_9_6_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i9_LC_9_6_2 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i9_LC_9_6_2  (
            .in0(N__51705),
            .in1(N__25214),
            .in2(N__25239),
            .in3(N__29137),
            .lcout(cmd_rdadctmp_9_adj_1514),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42424),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i11_LC_9_6_3 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i11_LC_9_6_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i11_LC_9_6_3 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i11_LC_9_6_3  (
            .in0(N__51699),
            .in1(N__25165),
            .in2(N__29139),
            .in3(N__25189),
            .lcout(cmd_rdadctmp_11_adj_1512),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42424),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i14_LC_9_6_4 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i14_LC_9_6_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i14_LC_9_6_4 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i14_LC_9_6_4  (
            .in0(N__51703),
            .in1(N__25487),
            .in2(N__25134),
            .in3(N__29135),
            .lcout(cmd_rdadctmp_14_adj_1509),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42424),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i12_LC_9_6_5 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i12_LC_9_6_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i12_LC_9_6_5 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i12_LC_9_6_5  (
            .in0(N__51700),
            .in1(N__25149),
            .in2(N__29140),
            .in3(N__25166),
            .lcout(cmd_rdadctmp_12_adj_1511),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42424),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i13_LC_9_6_6 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i13_LC_9_6_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i13_LC_9_6_6 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i13_LC_9_6_6  (
            .in0(N__25148),
            .in1(N__51702),
            .in2(N__25133),
            .in3(N__29134),
            .lcout(cmd_rdadctmp_13_adj_1510),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42424),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i15_LC_9_6_7 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i15_LC_9_6_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i15_LC_9_6_7 .LUT_INIT=16'b0010111100100000;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i15_LC_9_6_7  (
            .in0(N__25486),
            .in1(N__51706),
            .in2(N__29141),
            .in3(N__25468),
            .lcout(cmd_rdadctmp_15_adj_1508),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42424),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i7_4_lut_LC_9_7_0 .C_ON=1'b0;
    defparam \ADC_VDC.i7_4_lut_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i7_4_lut_LC_9_7_0 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \ADC_VDC.i7_4_lut_LC_9_7_0  (
            .in0(N__26975),
            .in1(N__26516),
            .in2(N__26631),
            .in3(N__26957),
            .lcout(\ADC_VDC.n19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i9_LC_9_7_1 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i9_LC_9_7_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i9_LC_9_7_1 .LUT_INIT=16'b0010111100100000;
    LogicCell40 \ADC_VDC.ADC_DATA_i9_LC_9_7_1  (
            .in0(N__25449),
            .in1(N__51475),
            .in2(N__31624),
            .in3(N__25430),
            .lcout(buf_adcdata_vdc_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42410),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i6_LC_9_7_2 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i6_LC_9_7_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i6_LC_9_7_2 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \ADC_VDC.ADC_DATA_i6_LC_9_7_2  (
            .in0(N__51473),
            .in1(N__31610),
            .in2(N__25397),
            .in3(N__25418),
            .lcout(buf_adcdata_vdc_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42410),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i0_LC_9_7_3 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i0_LC_9_7_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i0_LC_9_7_3 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i0_LC_9_7_3  (
            .in0(N__31609),
            .in1(N__51474),
            .in2(N__27293),
            .in3(N__25380),
            .lcout(buf_adcdata_vdc_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42410),
            .ce(),
            .sr(_gnd_net_));
    defparam n22473_bdd_4_lut_LC_9_7_4.C_ON=1'b0;
    defparam n22473_bdd_4_lut_LC_9_7_4.SEQ_MODE=4'b0000;
    defparam n22473_bdd_4_lut_LC_9_7_4.LUT_INIT=16'b1100111011000010;
    LogicCell40 n22473_bdd_4_lut_LC_9_7_4 (
            .in0(N__25970),
            .in1(N__25896),
            .in2(N__46469),
            .in3(N__29589),
            .lcout(n22476),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_5_i16_3_lut_LC_9_7_5.C_ON=1'b0;
    defparam mux_129_Mux_5_i16_3_lut_LC_9_7_5.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_5_i16_3_lut_LC_9_7_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_129_Mux_5_i16_3_lut_LC_9_7_5 (
            .in0(N__25368),
            .in1(N__33027),
            .in2(_gnd_net_),
            .in3(N__57105),
            .lcout(n16_adj_1628),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i12698_2_lut_LC_9_7_7 .C_ON=1'b0;
    defparam \ADC_VDC.i12698_2_lut_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i12698_2_lut_LC_9_7_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ADC_VDC.i12698_2_lut_LC_9_7_7  (
            .in0(N__51690),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26900),
            .lcout(\ADC_VDC.n15175 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i10_LC_9_8_0 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i10_LC_9_8_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i10_LC_9_8_0 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i10_LC_9_8_0  (
            .in0(N__31580),
            .in1(N__51496),
            .in2(N__27350),
            .in3(N__25344),
            .lcout(buf_adcdata_vdc_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42383),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i22_LC_9_8_2 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i22_LC_9_8_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i22_LC_9_8_2 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \ADC_VDC.ADC_DATA_i22_LC_9_8_2  (
            .in0(N__25332),
            .in1(N__51498),
            .in2(N__25676),
            .in3(N__31585),
            .lcout(buf_adcdata_vdc_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42383),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i2_LC_9_8_3 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i2_LC_9_8_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i2_LC_9_8_3 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \ADC_VDC.ADC_DATA_i2_LC_9_8_3  (
            .in0(N__51494),
            .in1(N__31583),
            .in2(N__25643),
            .in3(N__25659),
            .lcout(buf_adcdata_vdc_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42383),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i4_LC_9_8_4 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i4_LC_9_8_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i4_LC_9_8_4 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i4_LC_9_8_4  (
            .in0(N__31582),
            .in1(N__51497),
            .in2(N__25604),
            .in3(N__25620),
            .lcout(buf_adcdata_vdc_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42383),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i5_LC_9_8_5 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i5_LC_9_8_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i5_LC_9_8_5 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \ADC_VDC.ADC_DATA_i5_LC_9_8_5  (
            .in0(N__51495),
            .in1(N__25587),
            .in2(N__25571),
            .in3(N__31584),
            .lcout(buf_adcdata_vdc_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42383),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i23_LC_9_8_6 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i23_LC_9_8_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i23_LC_9_8_6 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i23_LC_9_8_6  (
            .in0(N__31581),
            .in1(N__51499),
            .in2(N__27138),
            .in3(N__25863),
            .lcout(buf_adcdata_vdc_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42383),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i21_LC_9_8_7 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i21_LC_9_8_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i21_LC_9_8_7 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i21_LC_9_8_7  (
            .in0(N__51746),
            .in1(N__25525),
            .in2(N__29138),
            .in3(N__25553),
            .lcout(cmd_rdadctmp_21_adj_1502),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42383),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadcbuf_i34_LC_9_9_0 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadcbuf_i34_LC_9_9_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadcbuf_i34_LC_9_9_0 .LUT_INIT=16'b0000010111001100;
    LogicCell40 \ADC_VDC.cmd_rdadcbuf_i34_LC_9_9_0  (
            .in0(N__51478),
            .in1(N__25506),
            .in2(N__25842),
            .in3(N__51744),
            .lcout(cmd_rdadcbuf_34),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42430),
            .ce(N__25833),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i9_4_lut_LC_9_9_2 .C_ON=1'b0;
    defparam \ADC_VDC.i9_4_lut_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i9_4_lut_LC_9_9_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.i9_4_lut_LC_9_9_2  (
            .in0(N__26649),
            .in1(N__26610),
            .in2(N__26673),
            .in3(N__26694),
            .lcout(),
            .ltout(\ADC_VDC.n21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i11_3_lut_LC_9_9_3 .C_ON=1'b0;
    defparam \ADC_VDC.i11_3_lut_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i11_3_lut_LC_9_9_3 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \ADC_VDC.i11_3_lut_LC_9_9_3  (
            .in0(_gnd_net_),
            .in1(N__25500),
            .in2(N__25491),
            .in3(N__30159),
            .lcout(\ADC_VDC.n18780 ),
            .ltout(\ADC_VDC.n18780_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_3_lut_LC_9_9_4 .C_ON=1'b0;
    defparam \ADC_VDC.i1_3_lut_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_3_lut_LC_9_9_4 .LUT_INIT=16'b1111111100111100;
    LogicCell40 \ADC_VDC.i1_3_lut_LC_9_9_4  (
            .in0(_gnd_net_),
            .in1(N__25862),
            .in2(N__25845),
            .in3(N__51212),
            .lcout(\ADC_VDC.n4_adj_1451 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_3_lut_4_lut_LC_9_9_5 .C_ON=1'b0;
    defparam \ADC_VDC.i1_3_lut_4_lut_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_3_lut_4_lut_LC_9_9_5 .LUT_INIT=16'b1100100011110000;
    LogicCell40 \ADC_VDC.i1_3_lut_4_lut_LC_9_9_5  (
            .in0(N__51211),
            .in1(N__51477),
            .in2(N__51759),
            .in3(N__51911),
            .lcout(\ADC_VDC.n13503 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19823_LC_9_10_0.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19823_LC_9_10_0.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19823_LC_9_10_0.LUT_INIT=16'b1101101011010000;
    LogicCell40 comm_cmd_0__bdd_4_lut_19823_LC_9_10_0 (
            .in0(N__46301),
            .in1(N__25824),
            .in2(N__56960),
            .in3(N__25715),
            .lcout(),
            .ltout(n22575_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22575_bdd_4_lut_LC_9_10_1.C_ON=1'b0;
    defparam n22575_bdd_4_lut_LC_9_10_1.SEQ_MODE=4'b0000;
    defparam n22575_bdd_4_lut_LC_9_10_1.LUT_INIT=16'b1111000010101100;
    LogicCell40 n22575_bdd_4_lut_LC_9_10_1 (
            .in0(N__25806),
            .in1(N__25778),
            .in2(N__25743),
            .in3(N__46302),
            .lcout(n22578),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i0_LC_9_10_2.C_ON=1'b0;
    defparam buf_cfgRTD_i0_LC_9_10_2.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i0_LC_9_10_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 buf_cfgRTD_i0_LC_9_10_2 (
            .in0(N__40448),
            .in1(N__39639),
            .in2(_gnd_net_),
            .in3(N__25716),
            .lcout(buf_cfgRTD_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55964),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_3_lut_LC_9_10_3.C_ON=1'b0;
    defparam i2_2_lut_3_lut_LC_9_10_3.SEQ_MODE=4'b0000;
    defparam i2_2_lut_3_lut_LC_9_10_3.LUT_INIT=16'b1101110111111111;
    LogicCell40 i2_2_lut_3_lut_LC_9_10_3 (
            .in0(N__47450),
            .in1(N__56787),
            .in2(_gnd_net_),
            .in3(N__46300),
            .lcout(),
            .ltout(n10902_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_279_LC_9_10_4.C_ON=1'b0;
    defparam i1_4_lut_adj_279_LC_9_10_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_279_LC_9_10_4.LUT_INIT=16'b1010101100000000;
    LogicCell40 i1_4_lut_adj_279_LC_9_10_4 (
            .in0(N__49383),
            .in1(N__30477),
            .in2(N__25692),
            .in3(N__55430),
            .lcout(n12624),
            .ltout(n12624_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i3_LC_9_10_5.C_ON=1'b0;
    defparam buf_cfgRTD_i3_LC_9_10_5.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i3_LC_9_10_5.LUT_INIT=16'b0000101011001010;
    LogicCell40 buf_cfgRTD_i3_LC_9_10_5 (
            .in0(N__25928),
            .in1(N__45348),
            .in2(N__25689),
            .in3(N__49384),
            .lcout(buf_cfgRTD_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55964),
            .ce(),
            .sr(_gnd_net_));
    defparam i36_4_lut_4_lut_LC_9_10_6.C_ON=1'b0;
    defparam i36_4_lut_4_lut_LC_9_10_6.SEQ_MODE=4'b0000;
    defparam i36_4_lut_4_lut_LC_9_10_6.LUT_INIT=16'b0100001011001110;
    LogicCell40 i36_4_lut_4_lut_LC_9_10_6 (
            .in0(N__46299),
            .in1(N__47165),
            .in2(N__56959),
            .in3(N__47449),
            .lcout(n30_adj_1499),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19809_LC_9_10_7.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19809_LC_9_10_7.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19809_LC_9_10_7.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_cmd_0__bdd_4_lut_19809_LC_9_10_7 (
            .in0(N__25927),
            .in1(N__56783),
            .in2(N__25914),
            .in3(N__46298),
            .lcout(n22473),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_idxvec_i0_LC_9_11_0.C_ON=1'b1;
    defparam data_idxvec_i0_LC_9_11_0.SEQ_MODE=4'b1000;
    defparam data_idxvec_i0_LC_9_11_0.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i0_LC_9_11_0 (
            .in0(N__43206),
            .in1(N__55402),
            .in2(N__43865),
            .in3(N__25887),
            .lcout(data_idxvec_0),
            .ltout(),
            .carryin(bfn_9_11_0_),
            .carryout(n19813),
            .clk(N__55975),
            .ce(N__26156),
            .sr(_gnd_net_));
    defparam data_idxvec_i1_LC_9_11_1.C_ON=1'b1;
    defparam data_idxvec_i1_LC_9_11_1.SEQ_MODE=4'b1000;
    defparam data_idxvec_i1_LC_9_11_1.LUT_INIT=16'b1010001110101100;
    LogicCell40 data_idxvec_i1_LC_9_11_1 (
            .in0(N__36170),
            .in1(N__44213),
            .in2(N__55465),
            .in3(N__25884),
            .lcout(data_idxvec_1),
            .ltout(),
            .carryin(n19813),
            .carryout(n19814),
            .clk(N__55975),
            .ce(N__26156),
            .sr(_gnd_net_));
    defparam data_idxvec_i2_LC_9_11_2.C_ON=1'b1;
    defparam data_idxvec_i2_LC_9_11_2.SEQ_MODE=4'b1000;
    defparam data_idxvec_i2_LC_9_11_2.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i2_LC_9_11_2 (
            .in0(N__34859),
            .in1(N__55406),
            .in2(N__35423),
            .in3(N__25881),
            .lcout(data_idxvec_2),
            .ltout(),
            .carryin(n19814),
            .carryout(n19815),
            .clk(N__55975),
            .ce(N__26156),
            .sr(_gnd_net_));
    defparam data_idxvec_i3_LC_9_11_3.C_ON=1'b1;
    defparam data_idxvec_i3_LC_9_11_3.SEQ_MODE=4'b1000;
    defparam data_idxvec_i3_LC_9_11_3.LUT_INIT=16'b1010001110101100;
    LogicCell40 data_idxvec_i3_LC_9_11_3 (
            .in0(N__36486),
            .in1(N__41237),
            .in2(N__55466),
            .in3(N__25878),
            .lcout(data_idxvec_3),
            .ltout(),
            .carryin(n19815),
            .carryout(n19816),
            .clk(N__55975),
            .ce(N__26156),
            .sr(_gnd_net_));
    defparam data_idxvec_i4_LC_9_11_4.C_ON=1'b1;
    defparam data_idxvec_i4_LC_9_11_4.SEQ_MODE=4'b1000;
    defparam data_idxvec_i4_LC_9_11_4.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i4_LC_9_11_4 (
            .in0(N__36198),
            .in1(N__55410),
            .in2(N__30677),
            .in3(N__25875),
            .lcout(data_idxvec_4),
            .ltout(),
            .carryin(n19816),
            .carryout(n19817),
            .clk(N__55975),
            .ce(N__26156),
            .sr(_gnd_net_));
    defparam data_idxvec_i5_LC_9_11_5.C_ON=1'b1;
    defparam data_idxvec_i5_LC_9_11_5.SEQ_MODE=4'b1000;
    defparam data_idxvec_i5_LC_9_11_5.LUT_INIT=16'b1010001110101100;
    LogicCell40 data_idxvec_i5_LC_9_11_5 (
            .in0(N__37249),
            .in1(N__32327),
            .in2(N__55467),
            .in3(N__25872),
            .lcout(data_idxvec_5),
            .ltout(),
            .carryin(n19817),
            .carryout(n19818),
            .clk(N__55975),
            .ce(N__26156),
            .sr(_gnd_net_));
    defparam data_idxvec_i6_LC_9_11_6.C_ON=1'b1;
    defparam data_idxvec_i6_LC_9_11_6.SEQ_MODE=4'b1000;
    defparam data_idxvec_i6_LC_9_11_6.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i6_LC_9_11_6 (
            .in0(N__31727),
            .in1(N__55414),
            .in2(N__43457),
            .in3(N__25869),
            .lcout(data_idxvec_6),
            .ltout(),
            .carryin(n19818),
            .carryout(n19819),
            .clk(N__55975),
            .ce(N__26156),
            .sr(_gnd_net_));
    defparam data_idxvec_i7_LC_9_11_7.C_ON=1'b1;
    defparam data_idxvec_i7_LC_9_11_7.SEQ_MODE=4'b1000;
    defparam data_idxvec_i7_LC_9_11_7.LUT_INIT=16'b1010001110101100;
    LogicCell40 data_idxvec_i7_LC_9_11_7 (
            .in0(N__32274),
            .in1(N__46544),
            .in2(N__55468),
            .in3(N__25866),
            .lcout(data_idxvec_7),
            .ltout(),
            .carryin(n19819),
            .carryout(n19820),
            .clk(N__55975),
            .ce(N__26156),
            .sr(_gnd_net_));
    defparam data_idxvec_i8_LC_9_12_0.C_ON=1'b1;
    defparam data_idxvec_i8_LC_9_12_0.SEQ_MODE=4'b1000;
    defparam data_idxvec_i8_LC_9_12_0.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i8_LC_9_12_0 (
            .in0(N__40452),
            .in1(N__55420),
            .in2(N__40925),
            .in3(N__26034),
            .lcout(data_idxvec_8),
            .ltout(),
            .carryin(bfn_9_12_0_),
            .carryout(n19821),
            .clk(N__55989),
            .ce(N__26160),
            .sr(_gnd_net_));
    defparam data_idxvec_i9_LC_9_12_1.C_ON=1'b1;
    defparam data_idxvec_i9_LC_9_12_1.SEQ_MODE=4'b1000;
    defparam data_idxvec_i9_LC_9_12_1.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i9_LC_9_12_1 (
            .in0(N__37452),
            .in1(N__55427),
            .in2(N__43106),
            .in3(N__26031),
            .lcout(data_idxvec_9),
            .ltout(),
            .carryin(n19821),
            .carryout(n19822),
            .clk(N__55989),
            .ce(N__26160),
            .sr(_gnd_net_));
    defparam data_idxvec_i10_LC_9_12_2.C_ON=1'b1;
    defparam data_idxvec_i10_LC_9_12_2.SEQ_MODE=4'b1000;
    defparam data_idxvec_i10_LC_9_12_2.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i10_LC_9_12_2 (
            .in0(N__32042),
            .in1(N__55421),
            .in2(N__40703),
            .in3(N__26028),
            .lcout(data_idxvec_10),
            .ltout(),
            .carryin(n19822),
            .carryout(n19823),
            .clk(N__55989),
            .ce(N__26160),
            .sr(_gnd_net_));
    defparam data_idxvec_i11_LC_9_12_3.C_ON=1'b1;
    defparam data_idxvec_i11_LC_9_12_3.SEQ_MODE=4'b1000;
    defparam data_idxvec_i11_LC_9_12_3.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i11_LC_9_12_3 (
            .in0(N__35253),
            .in1(N__55428),
            .in2(N__26061),
            .in3(N__26025),
            .lcout(data_idxvec_11),
            .ltout(),
            .carryin(n19823),
            .carryout(n19824),
            .clk(N__55989),
            .ce(N__26160),
            .sr(_gnd_net_));
    defparam data_idxvec_i12_LC_9_12_4.C_ON=1'b1;
    defparam data_idxvec_i12_LC_9_12_4.SEQ_MODE=4'b1000;
    defparam data_idxvec_i12_LC_9_12_4.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i12_LC_9_12_4 (
            .in0(N__37206),
            .in1(N__55422),
            .in2(N__40379),
            .in3(N__26022),
            .lcout(data_idxvec_12),
            .ltout(),
            .carryin(n19824),
            .carryout(n19825),
            .clk(N__55989),
            .ce(N__26160),
            .sr(_gnd_net_));
    defparam data_idxvec_i13_LC_9_12_5.C_ON=1'b1;
    defparam data_idxvec_i13_LC_9_12_5.SEQ_MODE=4'b1000;
    defparam data_idxvec_i13_LC_9_12_5.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i13_LC_9_12_5 (
            .in0(N__30721),
            .in1(N__55429),
            .in2(N__32411),
            .in3(N__26019),
            .lcout(data_idxvec_13),
            .ltout(),
            .carryin(n19825),
            .carryout(n19826),
            .clk(N__55989),
            .ce(N__26160),
            .sr(_gnd_net_));
    defparam data_idxvec_i14_LC_9_12_6.C_ON=1'b1;
    defparam data_idxvec_i14_LC_9_12_6.SEQ_MODE=4'b1000;
    defparam data_idxvec_i14_LC_9_12_6.LUT_INIT=16'b1000101110111000;
    LogicCell40 data_idxvec_i14_LC_9_12_6 (
            .in0(N__30359),
            .in1(N__55423),
            .in2(N__32600),
            .in3(N__26016),
            .lcout(data_idxvec_14),
            .ltout(),
            .carryin(n19826),
            .carryout(n19827),
            .clk(N__55989),
            .ce(N__26160),
            .sr(_gnd_net_));
    defparam data_idxvec_i15_LC_9_12_7.C_ON=1'b0;
    defparam data_idxvec_i15_LC_9_12_7.SEQ_MODE=4'b1000;
    defparam data_idxvec_i15_LC_9_12_7.LUT_INIT=16'b1010001110101100;
    LogicCell40 data_idxvec_i15_LC_9_12_7 (
            .in0(N__37472),
            .in1(N__28481),
            .in2(N__55469),
            .in3(N__26013),
            .lcout(data_idxvec_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55989),
            .ce(N__26160),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i19_LC_9_13_0 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i19_LC_9_13_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i19_LC_9_13_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i19_LC_9_13_0  (
            .in0(N__27999),
            .in1(N__27839),
            .in2(N__26010),
            .in3(N__25969),
            .lcout(buf_adcdata_vac_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56002),
            .ce(),
            .sr(_gnd_net_));
    defparam i15_4_lut_adj_295_LC_9_13_1.C_ON=1'b0;
    defparam i15_4_lut_adj_295_LC_9_13_1.SEQ_MODE=4'b0000;
    defparam i15_4_lut_adj_295_LC_9_13_1.LUT_INIT=16'b1010001011110111;
    LogicCell40 i15_4_lut_adj_295_LC_9_13_1 (
            .in0(N__55419),
            .in1(N__41124),
            .in2(N__49389),
            .in3(N__38946),
            .lcout(n12493),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15461_2_lut_3_lut_LC_9_13_2.C_ON=1'b0;
    defparam i15461_2_lut_3_lut_LC_9_13_2.SEQ_MODE=4'b0000;
    defparam i15461_2_lut_3_lut_LC_9_13_2.LUT_INIT=16'b0000000001000100;
    LogicCell40 i15461_2_lut_3_lut_LC_9_13_2 (
            .in0(N__54863),
            .in1(N__49567),
            .in2(_gnd_net_),
            .in3(N__54573),
            .lcout(n14_adj_1571),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22509_bdd_4_lut_LC_9_13_4.C_ON=1'b0;
    defparam n22509_bdd_4_lut_LC_9_13_4.SEQ_MODE=4'b0000;
    defparam n22509_bdd_4_lut_LC_9_13_4.LUT_INIT=16'b1110111000110000;
    LogicCell40 n22509_bdd_4_lut_LC_9_13_4 (
            .in0(N__26139),
            .in1(N__47536),
            .in2(N__32538),
            .in3(N__26040),
            .lcout(n22512),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i7_LC_9_13_5.C_ON=1'b0;
    defparam buf_device_acadc_i7_LC_9_13_5.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i7_LC_9_13_5.LUT_INIT=16'b0000101011001100;
    LogicCell40 buf_device_acadc_i7_LC_9_13_5 (
            .in0(N__49568),
            .in1(N__30806),
            .in2(N__49390),
            .in3(N__39515),
            .lcout(VAC_FLT0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56002),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i19_LC_9_13_6 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i19_LC_9_13_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i19_LC_9_13_6 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i19_LC_9_13_6  (
            .in0(N__28265),
            .in1(N__27445),
            .in2(N__26127),
            .in3(N__27840),
            .lcout(cmd_rdadctmp_19_adj_1473),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56002),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i2_LC_9_13_7.C_ON=1'b0;
    defparam buf_device_acadc_i2_LC_9_13_7.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i2_LC_9_13_7.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_device_acadc_i2_LC_9_13_7 (
            .in0(N__49365),
            .in1(N__39514),
            .in2(N__53458),
            .in3(N__26080),
            .lcout(IAC_OSR1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56002),
            .ce(),
            .sr(_gnd_net_));
    defparam i15228_2_lut_LC_9_14_0.C_ON=1'b0;
    defparam i15228_2_lut_LC_9_14_0.SEQ_MODE=4'b0000;
    defparam i15228_2_lut_LC_9_14_0.LUT_INIT=16'b1111111111001100;
    LogicCell40 i15228_2_lut_LC_9_14_0 (
            .in0(_gnd_net_),
            .in1(N__28839),
            .in2(_gnd_net_),
            .in3(N__28801),
            .lcout(n17728),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i2_LC_9_14_1.C_ON=1'b0;
    defparam buf_dds1_i2_LC_9_14_1.SEQ_MODE=4'b1000;
    defparam buf_dds1_i2_LC_9_14_1.LUT_INIT=16'b1110001000000000;
    LogicCell40 buf_dds1_i2_LC_9_14_1 (
            .in0(N__26264),
            .in1(N__46889),
            .in2(N__45480),
            .in3(N__46766),
            .lcout(buf_dds1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56019),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_3_i26_3_lut_LC_9_14_2.C_ON=1'b0;
    defparam mux_128_Mux_3_i26_3_lut_LC_9_14_2.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_3_i26_3_lut_LC_9_14_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_128_Mux_3_i26_3_lut_LC_9_14_2 (
            .in0(N__56913),
            .in1(N__26060),
            .in2(_gnd_net_),
            .in3(N__37955),
            .lcout(),
            .ltout(n26_adj_1678_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19760_LC_9_14_3.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19760_LC_9_14_3.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19760_LC_9_14_3.LUT_INIT=16'b1011101111000000;
    LogicCell40 comm_cmd_1__bdd_4_lut_19760_LC_9_14_3 (
            .in0(N__45753),
            .in1(N__47563),
            .in2(N__26043),
            .in3(N__46317),
            .lcout(n22509),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i2_LC_9_14_4.C_ON=1'b0;
    defparam buf_dds0_i2_LC_9_14_4.SEQ_MODE=4'b1000;
    defparam buf_dds0_i2_LC_9_14_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 buf_dds0_i2_LC_9_14_4 (
            .in0(N__34855),
            .in1(N__31448),
            .in2(_gnd_net_),
            .in3(N__41666),
            .lcout(buf_dds0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56019),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_2_i16_3_lut_LC_9_14_6.C_ON=1'b0;
    defparam mux_129_Mux_2_i16_3_lut_LC_9_14_6.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_2_i16_3_lut_LC_9_14_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_129_Mux_2_i16_3_lut_LC_9_14_6 (
            .in0(N__56914),
            .in1(N__26263),
            .in2(_gnd_net_),
            .in3(N__31447),
            .lcout(n16_adj_1645),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18607_3_lut_LC_9_14_7.C_ON=1'b0;
    defparam i18607_3_lut_LC_9_14_7.SEQ_MODE=4'b0000;
    defparam i18607_3_lut_LC_9_14_7.LUT_INIT=16'b1110111000100010;
    LogicCell40 i18607_3_lut_LC_9_14_7 (
            .in0(N__26418),
            .in1(N__47564),
            .in2(_gnd_net_),
            .in3(N__26250),
            .lcout(n21334),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i8_LC_9_15_0 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i8_LC_9_15_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i8_LC_9_15_0 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC.ADC_DATA_i8_LC_9_15_0  (
            .in0(N__27981),
            .in1(N__27833),
            .in2(N__43741),
            .in3(N__26238),
            .lcout(buf_adcdata_vac_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56033),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i25_LC_9_15_1 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i25_LC_9_15_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i25_LC_9_15_1 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i25_LC_9_15_1  (
            .in0(N__28240),
            .in1(N__26174),
            .in2(N__27856),
            .in3(N__26194),
            .lcout(cmd_rdadctmp_25_adj_1467),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56033),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i23_LC_9_15_2 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i23_LC_9_15_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i23_LC_9_15_2 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i23_LC_9_15_2  (
            .in0(N__26323),
            .in1(N__27834),
            .in2(N__26354),
            .in3(N__28238),
            .lcout(cmd_rdadctmp_23_adj_1469),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56033),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_rst_327_LC_9_15_3.C_ON=1'b0;
    defparam acadc_rst_327_LC_9_15_3.SEQ_MODE=4'b1000;
    defparam acadc_rst_327_LC_9_15_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 acadc_rst_327_LC_9_15_3 (
            .in0(N__45870),
            .in1(N__28046),
            .in2(_gnd_net_),
            .in3(N__35706),
            .lcout(acadc_rst),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56033),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i24_LC_9_15_4 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i24_LC_9_15_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i24_LC_9_15_4 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i24_LC_9_15_4  (
            .in0(N__26173),
            .in1(N__27835),
            .in2(N__26328),
            .in3(N__28239),
            .lcout(cmd_rdadctmp_24_adj_1468),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56033),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i9_LC_9_15_5.C_ON=1'b0;
    defparam buf_dds0_i9_LC_9_15_5.SEQ_MODE=4'b1000;
    defparam buf_dds0_i9_LC_9_15_5.LUT_INIT=16'b0101000011001100;
    LogicCell40 buf_dds0_i9_LC_9_15_5 (
            .in0(N__49369),
            .in1(N__31252),
            .in2(N__53462),
            .in3(N__41663),
            .lcout(buf_dds0_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56033),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i14_LC_9_15_6 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i14_LC_9_15_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i14_LC_9_15_6 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i14_LC_9_15_6  (
            .in0(N__27979),
            .in1(N__27832),
            .in2(N__26355),
            .in3(N__32461),
            .lcout(buf_adcdata_vac_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56033),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i15_LC_9_15_7 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i15_LC_9_15_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i15_LC_9_15_7 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC.ADC_DATA_i15_LC_9_15_7  (
            .in0(N__27831),
            .in1(N__27980),
            .in2(N__28432),
            .in3(N__26327),
            .lcout(buf_adcdata_vac_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56033),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_293_LC_9_16_0.C_ON=1'b0;
    defparam i1_4_lut_adj_293_LC_9_16_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_293_LC_9_16_0.LUT_INIT=16'b1100000011001000;
    LogicCell40 i1_4_lut_adj_293_LC_9_16_0 (
            .in0(N__26313),
            .in1(N__55464),
            .in2(N__49370),
            .in3(N__44114),
            .lcout(n12654),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i11_LC_9_16_2.C_ON=1'b0;
    defparam buf_dds1_i11_LC_9_16_2.SEQ_MODE=4'b1000;
    defparam buf_dds1_i11_LC_9_16_2.LUT_INIT=16'b1110001000000000;
    LogicCell40 buf_dds1_i11_LC_9_16_2 (
            .in0(N__26441),
            .in1(N__46885),
            .in2(N__45357),
            .in3(N__46732),
            .lcout(buf_dds1_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56049),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i16_LC_9_16_4 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i16_LC_9_16_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i16_LC_9_16_4 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i16_LC_9_16_4  (
            .in0(N__33796),
            .in1(N__29385),
            .in2(N__26300),
            .in3(N__38553),
            .lcout(cmd_rdadctmp_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56049),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i6_LC_9_16_6.C_ON=1'b0;
    defparam buf_device_acadc_i6_LC_9_16_6.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i6_LC_9_16_6.LUT_INIT=16'b0011000010101010;
    LogicCell40 buf_device_acadc_i6_LC_9_16_6 (
            .in0(N__27373),
            .in1(N__49305),
            .in2(N__52290),
            .in3(N__39538),
            .lcout(VAC_OSR1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56049),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i10_LC_9_16_7.C_ON=1'b0;
    defparam buf_dds0_i10_LC_9_16_7.SEQ_MODE=4'b1000;
    defparam buf_dds0_i10_LC_9_16_7.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_dds0_i10_LC_9_16_7 (
            .in0(N__49304),
            .in1(N__41664),
            .in2(N__45879),
            .in3(N__31081),
            .lcout(buf_dds0_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56049),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i19_LC_9_17_0 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i19_LC_9_17_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i19_LC_9_17_0 .LUT_INIT=16'b1101111110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i19_LC_9_17_0  (
            .in0(N__38500),
            .in1(N__26409),
            .in2(N__38770),
            .in3(N__26461),
            .lcout(buf_adcdata_iac_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56063),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i17_LC_9_17_2 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i17_LC_9_17_2 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i17_LC_9_17_2 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i17_LC_9_17_2  (
            .in0(N__38501),
            .in1(N__33803),
            .in2(N__33776),
            .in3(N__29382),
            .lcout(cmd_rdadctmp_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56063),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i4_LC_9_17_3.C_ON=1'b0;
    defparam buf_device_acadc_i4_LC_9_17_3.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i4_LC_9_17_3.LUT_INIT=16'b0000110010101010;
    LogicCell40 buf_device_acadc_i4_LC_9_17_3 (
            .in0(N__26486),
            .in1(N__45352),
            .in2(N__49391),
            .in3(N__39539),
            .lcout(IAC_FLT1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56063),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_start_329_LC_9_17_4.C_ON=1'b0;
    defparam eis_start_329_LC_9_17_4.SEQ_MODE=4'b1000;
    defparam eis_start_329_LC_9_17_4.LUT_INIT=16'b1011101110001000;
    LogicCell40 eis_start_329_LC_9_17_4 (
            .in0(N__45648),
            .in1(N__28050),
            .in2(_gnd_net_),
            .in3(N__31028),
            .lcout(eis_start),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56063),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19842_LC_9_17_5.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19842_LC_9_17_5.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19842_LC_9_17_5.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_cmd_0__bdd_4_lut_19842_LC_9_17_5 (
            .in0(N__26485),
            .in1(N__57097),
            .in2(N__26465),
            .in3(N__46406),
            .lcout(),
            .ltout(n22605_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22605_bdd_4_lut_LC_9_17_6.C_ON=1'b0;
    defparam n22605_bdd_4_lut_LC_9_17_6.SEQ_MODE=4'b0000;
    defparam n22605_bdd_4_lut_LC_9_17_6.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22605_bdd_4_lut_LC_9_17_6 (
            .in0(N__46407),
            .in1(N__31366),
            .in2(N__26445),
            .in3(N__26431),
            .lcout(n22608),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i18_LC_9_17_7 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i18_LC_9_17_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i18_LC_9_17_7 .LUT_INIT=16'b1101100001010000;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i18_LC_9_17_7  (
            .in0(N__29381),
            .in1(N__38502),
            .in2(N__38264),
            .in3(N__33772),
            .lcout(cmd_rdadctmp_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56063),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i27_LC_9_18_0 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i27_LC_9_18_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i27_LC_9_18_0 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i27_LC_9_18_0  (
            .in0(N__38583),
            .in1(N__26401),
            .in2(N__32786),
            .in3(N__29372),
            .lcout(cmd_rdadctmp_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56077),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i11_LC_9_18_1 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i11_LC_9_18_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i11_LC_9_18_1 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \ADC_IAC.ADC_DATA_i11_LC_9_18_1  (
            .in0(N__38742),
            .in1(N__26385),
            .in2(N__41296),
            .in3(N__38584),
            .lcout(buf_adcdata_iac_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56077),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i25_LC_9_18_3 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i25_LC_9_18_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i25_LC_9_18_3 .LUT_INIT=16'b1110001000100010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i25_LC_9_18_3  (
            .in0(N__28879),
            .in1(N__29373),
            .in2(N__26370),
            .in3(N__38586),
            .lcout(cmd_rdadctmp_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56077),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i16_LC_9_18_4 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i16_LC_9_18_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i16_LC_9_18_4 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_IAC.ADC_DATA_i16_LC_9_18_4  (
            .in0(N__38582),
            .in1(N__38743),
            .in2(N__39142),
            .in3(N__26369),
            .lcout(buf_adcdata_iac_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56077),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i24_LC_9_18_5 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i24_LC_9_18_5 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i24_LC_9_18_5 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i24_LC_9_18_5  (
            .in0(N__26365),
            .in1(N__38585),
            .in2(N__29390),
            .in3(N__28745),
            .lcout(cmd_rdadctmp_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56077),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i31_LC_9_18_7 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i31_LC_9_18_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i31_LC_9_18_7 .LUT_INIT=16'b1100101000001010;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i31_LC_9_18_7  (
            .in0(N__29213),
            .in1(N__38587),
            .in2(N__29391),
            .in3(N__26584),
            .lcout(cmd_rdadctmp_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56077),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i16257_3_lut_LC_10_4_1 .C_ON=1'b0;
    defparam \ADC_VDC.i16257_3_lut_LC_10_4_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i16257_3_lut_LC_10_4_1 .LUT_INIT=16'b0111011101100110;
    LogicCell40 \ADC_VDC.i16257_3_lut_LC_10_4_1  (
            .in0(N__51154),
            .in1(N__51882),
            .in2(_gnd_net_),
            .in3(N__26565),
            .lcout(),
            .ltout(\ADC_VDC.n18783_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.adc_state_i1_LC_10_4_2 .C_ON=1'b0;
    defparam \ADC_VDC.adc_state_i1_LC_10_4_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.adc_state_i1_LC_10_4_2 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \ADC_VDC.adc_state_i1_LC_10_4_2  (
            .in0(N__51329),
            .in1(N__51636),
            .in2(N__26553),
            .in3(N__29148),
            .lcout(\ADC_VDC.adc_state_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42398),
            .ce(N__26550),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i19425_4_lut_LC_10_4_3 .C_ON=1'b0;
    defparam \ADC_VDC.i19425_4_lut_LC_10_4_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i19425_4_lut_LC_10_4_3 .LUT_INIT=16'b1100111011011111;
    LogicCell40 \ADC_VDC.i19425_4_lut_LC_10_4_3  (
            .in0(N__51635),
            .in1(N__51328),
            .in2(N__31398),
            .in3(N__26544),
            .lcout(\ADC_VDC.n16_adj_1450 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i39_3_lut_4_lut_LC_10_4_5 .C_ON=1'b0;
    defparam \ADC_VDC.i39_3_lut_4_lut_LC_10_4_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i39_3_lut_4_lut_LC_10_4_5 .LUT_INIT=16'b1110010000110011;
    LogicCell40 \ADC_VDC.i39_3_lut_4_lut_LC_10_4_5  (
            .in0(N__51153),
            .in1(N__51975),
            .in2(N__31662),
            .in3(N__51881),
            .lcout(\ADC_VDC.n18 ),
            .ltout(\ADC_VDC.n18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i19428_4_lut_LC_10_4_6 .C_ON=1'b0;
    defparam \ADC_VDC.i19428_4_lut_LC_10_4_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i19428_4_lut_LC_10_4_6 .LUT_INIT=16'b1010101111101111;
    LogicCell40 \ADC_VDC.i19428_4_lut_LC_10_4_6  (
            .in0(N__51327),
            .in1(N__51634),
            .in2(N__26538),
            .in3(N__29687),
            .lcout(\ADC_VDC.n16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i18466_2_lut_3_lut_LC_10_4_7 .C_ON=1'b0;
    defparam \ADC_VDC.i18466_2_lut_3_lut_LC_10_4_7 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i18466_2_lut_3_lut_LC_10_4_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \ADC_VDC.i18466_2_lut_3_lut_LC_10_4_7  (
            .in0(N__51152),
            .in1(N__51974),
            .in2(_gnd_net_),
            .in3(N__51880),
            .lcout(\ADC_VDC.n21193 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i7_LC_10_5_4.C_ON=1'b0;
    defparam buf_control_i7_LC_10_5_4.SEQ_MODE=4'b1000;
    defparam buf_control_i7_LC_10_5_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 buf_control_i7_LC_10_5_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26535),
            .lcout(buf_control_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55940),
            .ce(N__42069),
            .sr(N__42093));
    defparam \ADC_VDC.avg_cnt_i0_LC_10_6_0 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i0_LC_10_6_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i0_LC_10_6_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i0_LC_10_6_0  (
            .in0(_gnd_net_),
            .in1(N__26517),
            .in2(_gnd_net_),
            .in3(N__26505),
            .lcout(\ADC_VDC.avg_cnt_0 ),
            .ltout(),
            .carryin(bfn_10_6_0_),
            .carryout(\ADC_VDC.n19877 ),
            .clk(N__42362),
            .ce(N__26940),
            .sr(N__26864));
    defparam \ADC_VDC.avg_cnt_i1_LC_10_6_1 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i1_LC_10_6_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i1_LC_10_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i1_LC_10_6_1  (
            .in0(_gnd_net_),
            .in1(N__26690),
            .in2(_gnd_net_),
            .in3(N__26676),
            .lcout(\ADC_VDC.avg_cnt_1 ),
            .ltout(),
            .carryin(\ADC_VDC.n19877 ),
            .carryout(\ADC_VDC.n19878 ),
            .clk(N__42362),
            .ce(N__26940),
            .sr(N__26864));
    defparam \ADC_VDC.avg_cnt_i2_LC_10_6_2 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i2_LC_10_6_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i2_LC_10_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i2_LC_10_6_2  (
            .in0(_gnd_net_),
            .in1(N__26669),
            .in2(_gnd_net_),
            .in3(N__26655),
            .lcout(\ADC_VDC.avg_cnt_2 ),
            .ltout(),
            .carryin(\ADC_VDC.n19878 ),
            .carryout(\ADC_VDC.n19879 ),
            .clk(N__42362),
            .ce(N__26940),
            .sr(N__26864));
    defparam \ADC_VDC.avg_cnt_i3_LC_10_6_3 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i3_LC_10_6_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i3_LC_10_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i3_LC_10_6_3  (
            .in0(_gnd_net_),
            .in1(N__30171),
            .in2(_gnd_net_),
            .in3(N__26652),
            .lcout(\ADC_VDC.avg_cnt_3 ),
            .ltout(),
            .carryin(\ADC_VDC.n19879 ),
            .carryout(\ADC_VDC.n19880 ),
            .clk(N__42362),
            .ce(N__26940),
            .sr(N__26864));
    defparam \ADC_VDC.avg_cnt_i4_LC_10_6_4 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i4_LC_10_6_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i4_LC_10_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i4_LC_10_6_4  (
            .in0(_gnd_net_),
            .in1(N__26648),
            .in2(_gnd_net_),
            .in3(N__26634),
            .lcout(\ADC_VDC.avg_cnt_4 ),
            .ltout(),
            .carryin(\ADC_VDC.n19880 ),
            .carryout(\ADC_VDC.n19881 ),
            .clk(N__42362),
            .ce(N__26940),
            .sr(N__26864));
    defparam \ADC_VDC.avg_cnt_i5_LC_10_6_5 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i5_LC_10_6_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i5_LC_10_6_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i5_LC_10_6_5  (
            .in0(_gnd_net_),
            .in1(N__26630),
            .in2(_gnd_net_),
            .in3(N__26616),
            .lcout(\ADC_VDC.avg_cnt_5 ),
            .ltout(),
            .carryin(\ADC_VDC.n19881 ),
            .carryout(\ADC_VDC.n19882 ),
            .clk(N__42362),
            .ce(N__26940),
            .sr(N__26864));
    defparam \ADC_VDC.avg_cnt_i6_LC_10_6_6 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i6_LC_10_6_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i6_LC_10_6_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i6_LC_10_6_6  (
            .in0(_gnd_net_),
            .in1(N__30185),
            .in2(_gnd_net_),
            .in3(N__26613),
            .lcout(\ADC_VDC.avg_cnt_6 ),
            .ltout(),
            .carryin(\ADC_VDC.n19882 ),
            .carryout(\ADC_VDC.n19883 ),
            .clk(N__42362),
            .ce(N__26940),
            .sr(N__26864));
    defparam \ADC_VDC.avg_cnt_i7_LC_10_6_7 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i7_LC_10_6_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i7_LC_10_6_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i7_LC_10_6_7  (
            .in0(_gnd_net_),
            .in1(N__26609),
            .in2(_gnd_net_),
            .in3(N__26595),
            .lcout(\ADC_VDC.avg_cnt_7 ),
            .ltout(),
            .carryin(\ADC_VDC.n19883 ),
            .carryout(\ADC_VDC.n19884 ),
            .clk(N__42362),
            .ce(N__26940),
            .sr(N__26864));
    defparam \ADC_VDC.avg_cnt_i8_LC_10_7_0 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i8_LC_10_7_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i8_LC_10_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i8_LC_10_7_0  (
            .in0(_gnd_net_),
            .in1(N__30198),
            .in2(_gnd_net_),
            .in3(N__26592),
            .lcout(\ADC_VDC.avg_cnt_8 ),
            .ltout(),
            .carryin(bfn_10_7_0_),
            .carryout(\ADC_VDC.n19885 ),
            .clk(N__42409),
            .ce(N__26929),
            .sr(N__26863));
    defparam \ADC_VDC.avg_cnt_i9_LC_10_7_1 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i9_LC_10_7_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i9_LC_10_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i9_LC_10_7_1  (
            .in0(_gnd_net_),
            .in1(N__30210),
            .in2(_gnd_net_),
            .in3(N__26589),
            .lcout(\ADC_VDC.avg_cnt_9 ),
            .ltout(),
            .carryin(\ADC_VDC.n19885 ),
            .carryout(\ADC_VDC.n19886 ),
            .clk(N__42409),
            .ce(N__26929),
            .sr(N__26863));
    defparam \ADC_VDC.avg_cnt_i10_LC_10_7_2 .C_ON=1'b1;
    defparam \ADC_VDC.avg_cnt_i10_LC_10_7_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i10_LC_10_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i10_LC_10_7_2  (
            .in0(_gnd_net_),
            .in1(N__26976),
            .in2(_gnd_net_),
            .in3(N__26964),
            .lcout(\ADC_VDC.avg_cnt_10 ),
            .ltout(),
            .carryin(\ADC_VDC.n19886 ),
            .carryout(\ADC_VDC.n19887 ),
            .clk(N__42409),
            .ce(N__26929),
            .sr(N__26863));
    defparam \ADC_VDC.avg_cnt_i11_LC_10_7_3 .C_ON=1'b0;
    defparam \ADC_VDC.avg_cnt_i11_LC_10_7_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.avg_cnt_i11_LC_10_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.avg_cnt_i11_LC_10_7_3  (
            .in0(_gnd_net_),
            .in1(N__26958),
            .in2(_gnd_net_),
            .in3(N__26961),
            .lcout(\ADC_VDC.avg_cnt_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42409),
            .ce(N__26929),
            .sr(N__26863));
    defparam \ADC_VDC.ADC_DATA_i12_LC_10_8_0 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i12_LC_10_8_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i12_LC_10_8_0 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i12_LC_10_8_0  (
            .in0(N__31587),
            .in1(N__51483),
            .in2(N__28019),
            .in3(N__26796),
            .lcout(buf_adcdata_vdc_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42425),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i7_LC_10_8_1 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i7_LC_10_8_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i7_LC_10_8_1 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \ADC_VDC.ADC_DATA_i7_LC_10_8_1  (
            .in0(N__26781),
            .in1(N__26759),
            .in2(N__51501),
            .in3(N__31589),
            .lcout(buf_adcdata_vdc_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42425),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_5_i23_3_lut_LC_10_8_2.C_ON=1'b0;
    defparam mux_128_Mux_5_i23_3_lut_LC_10_8_2.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_5_i23_3_lut_LC_10_8_2.LUT_INIT=16'b1110111001000100;
    LogicCell40 mux_128_Mux_5_i23_3_lut_LC_10_8_2 (
            .in0(N__57185),
            .in1(N__35996),
            .in2(_gnd_net_),
            .in3(N__33048),
            .lcout(n23_adj_1668),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_3_lut_4_lut_adj_35_LC_10_8_3 .C_ON=1'b0;
    defparam \ADC_VDC.i1_3_lut_4_lut_adj_35_LC_10_8_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_3_lut_4_lut_adj_35_LC_10_8_3 .LUT_INIT=16'b1000100011001000;
    LogicCell40 \ADC_VDC.i1_3_lut_4_lut_adj_35_LC_10_8_3  (
            .in0(N__51480),
            .in1(N__51745),
            .in2(N__51915),
            .in3(N__51197),
            .lcout(n11891),
            .ltout(n11891_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i15_LC_10_8_4 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i15_LC_10_8_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i15_LC_10_8_4 .LUT_INIT=16'b0011101000001010;
    LogicCell40 \ADC_VDC.ADC_DATA_i15_LC_10_8_4  (
            .in0(N__28403),
            .in1(N__51484),
            .in2(N__26748),
            .in3(N__26745),
            .lcout(buf_adcdata_vdc_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42425),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i14_LC_10_8_5 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i14_LC_10_8_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i14_LC_10_8_5 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \ADC_VDC.ADC_DATA_i14_LC_10_8_5  (
            .in0(N__51481),
            .in1(N__31588),
            .in2(N__32489),
            .in3(N__26727),
            .lcout(buf_adcdata_vdc_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42425),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i11_LC_10_8_6 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i11_LC_10_8_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i11_LC_10_8_6 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \ADC_VDC.ADC_DATA_i11_LC_10_8_6  (
            .in0(N__31586),
            .in1(N__51482),
            .in2(N__35069),
            .in3(N__26709),
            .lcout(buf_adcdata_vdc_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42425),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_7_i23_3_lut_LC_10_9_0.C_ON=1'b0;
    defparam mux_128_Mux_7_i23_3_lut_LC_10_9_0.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_7_i23_3_lut_LC_10_9_0.LUT_INIT=16'b1110111000100010;
    LogicCell40 mux_128_Mux_7_i23_3_lut_LC_10_9_0 (
            .in0(N__27198),
            .in1(N__56957),
            .in2(_gnd_net_),
            .in3(N__31184),
            .lcout(n23_adj_1658),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.SCLK_27_LC_10_9_1 .C_ON=1'b0;
    defparam \CLK_DDS.SCLK_27_LC_10_9_1 .SEQ_MODE=4'b1000;
    defparam \CLK_DDS.SCLK_27_LC_10_9_1 .LUT_INIT=16'b0111001000110001;
    LogicCell40 \CLK_DDS.SCLK_27_LC_10_9_1  (
            .in0(N__29840),
            .in1(N__30093),
            .in2(N__27179),
            .in3(N__29951),
            .lcout(DDS_SCK1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55952),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19833_LC_10_9_2.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19833_LC_10_9_2.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19833_LC_10_9_2.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_cmd_0__bdd_4_lut_19833_LC_10_9_2 (
            .in0(N__27014),
            .in1(N__56958),
            .in2(N__27162),
            .in3(N__46308),
            .lcout(),
            .ltout(n22593_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22593_bdd_4_lut_LC_10_9_3.C_ON=1'b0;
    defparam n22593_bdd_4_lut_LC_10_9_3.SEQ_MODE=4'b0000;
    defparam n22593_bdd_4_lut_LC_10_9_3.LUT_INIT=16'b1110010111100000;
    LogicCell40 n22593_bdd_4_lut_LC_10_9_3 (
            .in0(N__46309),
            .in1(N__27137),
            .in2(N__27123),
            .in3(N__27113),
            .lcout(n21240),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i6_LC_10_9_5.C_ON=1'b0;
    defparam buf_cfgRTD_i6_LC_10_9_5.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i6_LC_10_9_5.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_cfgRTD_i6_LC_10_9_5 (
            .in0(N__49377),
            .in1(N__39641),
            .in2(N__49569),
            .in3(N__27053),
            .lcout(buf_cfgRTD_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55952),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i7_LC_10_9_6.C_ON=1'b0;
    defparam buf_cfgRTD_i7_LC_10_9_6.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i7_LC_10_9_6.LUT_INIT=16'b0011000010101010;
    LogicCell40 buf_cfgRTD_i7_LC_10_9_6 (
            .in0(N__27015),
            .in1(N__49378),
            .in2(N__42554),
            .in3(N__39642),
            .lcout(buf_cfgRTD_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55952),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_60_LC_10_9_7.C_ON=1'b0;
    defparam i1_4_lut_adj_60_LC_10_9_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_60_LC_10_9_7.LUT_INIT=16'b0011000000110001;
    LogicCell40 i1_4_lut_adj_60_LC_10_9_7 (
            .in0(N__46307),
            .in1(N__37589),
            .in2(N__26985),
            .in3(N__47702),
            .lcout(comm_state_3_N_460_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_59_LC_10_10_0.C_ON=1'b0;
    defparam i1_2_lut_adj_59_LC_10_10_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_59_LC_10_10_0.LUT_INIT=16'b0011001100000000;
    LogicCell40 i1_2_lut_adj_59_LC_10_10_0 (
            .in0(_gnd_net_),
            .in1(N__56867),
            .in2(_gnd_net_),
            .in3(N__46306),
            .lcout(n5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i13_LC_10_10_1 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i13_LC_10_10_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i13_LC_10_10_1 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_VAC.ADC_DATA_i13_LC_10_10_1  (
            .in0(N__27998),
            .in1(N__27842),
            .in2(N__28313),
            .in3(N__28088),
            .lcout(buf_adcdata_vac_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55956),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_307_LC_10_10_2.C_ON=1'b0;
    defparam i1_2_lut_adj_307_LC_10_10_2.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_307_LC_10_10_2.LUT_INIT=16'b1100110000000000;
    LogicCell40 i1_2_lut_adj_307_LC_10_10_2 (
            .in0(_gnd_net_),
            .in1(N__47164),
            .in2(_gnd_net_),
            .in3(N__32390),
            .lcout(n4_adj_1455),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i11_LC_10_10_4 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i11_LC_10_10_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i11_LC_10_10_4 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_VAC.ADC_DATA_i11_LC_10_10_4  (
            .in0(N__27841),
            .in1(N__27997),
            .in2(N__27465),
            .in3(N__35044),
            .lcout(buf_adcdata_vac_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55956),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i4_LC_10_10_5.C_ON=1'b0;
    defparam buf_cfgRTD_i4_LC_10_10_5.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i4_LC_10_10_5.LUT_INIT=16'b0111010000110000;
    LogicCell40 buf_cfgRTD_i4_LC_10_10_5 (
            .in0(N__49385),
            .in1(N__39640),
            .in2(N__34999),
            .in3(N__47799),
            .lcout(buf_cfgRTD_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55956),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_5_i19_3_lut_LC_10_10_6.C_ON=1'b0;
    defparam mux_128_Mux_5_i19_3_lut_LC_10_10_6.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_5_i19_3_lut_LC_10_10_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_128_Mux_5_i19_3_lut_LC_10_10_6 (
            .in0(N__29508),
            .in1(N__27425),
            .in2(_gnd_net_),
            .in3(N__56868),
            .lcout(n19_adj_1666),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_5_i17_3_lut_LC_10_10_7.C_ON=1'b0;
    defparam mux_128_Mux_5_i17_3_lut_LC_10_10_7.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_5_i17_3_lut_LC_10_10_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_128_Mux_5_i17_3_lut_LC_10_10_7 (
            .in0(N__56869),
            .in1(N__28940),
            .in2(_gnd_net_),
            .in3(N__27383),
            .lcout(n17_adj_1665),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_2_i19_3_lut_LC_10_11_0.C_ON=1'b0;
    defparam mux_129_Mux_2_i19_3_lut_LC_10_11_0.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_2_i19_3_lut_LC_10_11_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_129_Mux_2_i19_3_lut_LC_10_11_0 (
            .in0(N__27354),
            .in1(N__27329),
            .in2(_gnd_net_),
            .in3(N__57026),
            .lcout(n19_adj_1646),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_0_i19_3_lut_LC_10_11_1.C_ON=1'b0;
    defparam mux_130_Mux_0_i19_3_lut_LC_10_11_1.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_0_i19_3_lut_LC_10_11_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_130_Mux_0_i19_3_lut_LC_10_11_1 (
            .in0(N__57025),
            .in1(N__27294),
            .in2(_gnd_net_),
            .in3(N__27272),
            .lcout(),
            .ltout(n19_adj_1534_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_0_i22_3_lut_LC_10_11_2.C_ON=1'b0;
    defparam mux_130_Mux_0_i22_3_lut_LC_10_11_2.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_0_i22_3_lut_LC_10_11_2.LUT_INIT=16'b1111000011001100;
    LogicCell40 mux_130_Mux_0_i22_3_lut_LC_10_11_2 (
            .in0(_gnd_net_),
            .in1(N__27230),
            .in2(N__27201),
            .in3(N__47519),
            .lcout(n22_adj_1532),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i0_LC_10_11_3.C_ON=1'b0;
    defparam comm_cmd_i0_LC_10_11_3.SEQ_MODE=4'b1000;
    defparam comm_cmd_i0_LC_10_11_3.LUT_INIT=16'b1100000010101010;
    LogicCell40 comm_cmd_i0_LC_10_11_3 (
            .in0(N__57028),
            .in1(N__48696),
            .in2(N__50980),
            .in3(N__37531),
            .lcout(comm_cmd_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55965),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19701_LC_10_11_4.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19701_LC_10_11_4.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19701_LC_10_11_4.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_19701_LC_10_11_4 (
            .in0(N__28359),
            .in1(N__46310),
            .in2(N__28347),
            .in3(N__47518),
            .lcout(n22431),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_5_i19_3_lut_LC_10_11_5.C_ON=1'b0;
    defparam mux_129_Mux_5_i19_3_lut_LC_10_11_5.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_5_i19_3_lut_LC_10_11_5.LUT_INIT=16'b1110111001000100;
    LogicCell40 mux_129_Mux_5_i19_3_lut_LC_10_11_5 (
            .in0(N__57027),
            .in1(N__28312),
            .in2(_gnd_net_),
            .in3(N__29631),
            .lcout(),
            .ltout(n19_adj_1629_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19653_LC_10_11_6.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19653_LC_10_11_6.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19653_LC_10_11_6.LUT_INIT=16'b1011100011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_19653_LC_10_11_6 (
            .in0(N__28287),
            .in1(N__46311),
            .in2(N__28272),
            .in3(N__47520),
            .lcout(n22365),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_adj_261_LC_10_11_7.C_ON=1'b0;
    defparam i2_4_lut_adj_261_LC_10_11_7.SEQ_MODE=4'b0000;
    defparam i2_4_lut_adj_261_LC_10_11_7.LUT_INIT=16'b0000000000000100;
    LogicCell40 i2_4_lut_adj_261_LC_10_11_7 (
            .in0(N__31154),
            .in1(N__55418),
            .in2(N__28062),
            .in3(N__54008),
            .lcout(n10695),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.cmd_rdadctmp_i21_LC_10_12_0 .C_ON=1'b0;
    defparam \ADC_VAC.cmd_rdadctmp_i21_LC_10_12_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.cmd_rdadctmp_i21_LC_10_12_0 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_VAC.cmd_rdadctmp_i21_LC_10_12_0  (
            .in0(N__27843),
            .in1(N__28078),
            .in2(N__27513),
            .in3(N__28266),
            .lcout(cmd_rdadctmp_21_adj_1471),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55976),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_6__I_0_368_i8_2_lut_LC_10_12_1.C_ON=1'b0;
    defparam comm_cmd_6__I_0_368_i8_2_lut_LC_10_12_1.SEQ_MODE=4'b0000;
    defparam comm_cmd_6__I_0_368_i8_2_lut_LC_10_12_1.LUT_INIT=16'b1111111100110011;
    LogicCell40 comm_cmd_6__I_0_368_i8_2_lut_LC_10_12_1 (
            .in0(_gnd_net_),
            .in1(N__46291),
            .in2(_gnd_net_),
            .in3(N__47601),
            .lcout(n8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_stop_328_LC_10_12_2.C_ON=1'b0;
    defparam eis_stop_328_LC_10_12_2.SEQ_MODE=4'b1000;
    defparam eis_stop_328_LC_10_12_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 eis_stop_328_LC_10_12_2 (
            .in0(N__53448),
            .in1(N__28034),
            .in2(_gnd_net_),
            .in3(N__43028),
            .lcout(eis_stop),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55976),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_4_i19_3_lut_LC_10_12_3.C_ON=1'b0;
    defparam mux_129_Mux_4_i19_3_lut_LC_10_12_3.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_4_i19_3_lut_LC_10_12_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_129_Mux_4_i19_3_lut_LC_10_12_3 (
            .in0(N__28023),
            .in1(N__27481),
            .in2(_gnd_net_),
            .in3(N__56873),
            .lcout(n19_adj_1634),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VAC.ADC_DATA_i12_LC_10_12_5 .C_ON=1'b0;
    defparam \ADC_VAC.ADC_DATA_i12_LC_10_12_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VAC.ADC_DATA_i12_LC_10_12_5 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \ADC_VAC.ADC_DATA_i12_LC_10_12_5  (
            .in0(N__28000),
            .in1(N__27482),
            .in2(N__27857),
            .in3(N__27512),
            .lcout(buf_adcdata_vac_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55976),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i12_LC_10_12_6.C_ON=1'b0;
    defparam buf_dds1_i12_LC_10_12_6.SEQ_MODE=4'b1000;
    defparam buf_dds1_i12_LC_10_12_6.LUT_INIT=16'b1110001000000000;
    LogicCell40 buf_dds1_i12_LC_10_12_6 (
            .in0(N__36277),
            .in1(N__46898),
            .in2(N__47819),
            .in3(N__46746),
            .lcout(buf_dds1_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55976),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19658_LC_10_13_0.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19658_LC_10_13_0.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19658_LC_10_13_0.LUT_INIT=16'b1111010110001000;
    LogicCell40 comm_cmd_0__bdd_4_lut_19658_LC_10_13_0 (
            .in0(N__46369),
            .in1(N__28994),
            .in2(N__29202),
            .in3(N__56899),
            .lcout(n22371),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_4_lut_4_lut_LC_10_13_1.C_ON=1'b0;
    defparam i3_4_lut_4_lut_LC_10_13_1.SEQ_MODE=4'b0000;
    defparam i3_4_lut_4_lut_LC_10_13_1.LUT_INIT=16'b0010000000000000;
    LogicCell40 i3_4_lut_4_lut_LC_10_13_1 (
            .in0(N__30963),
            .in1(N__35709),
            .in2(N__28665),
            .in3(N__37771),
            .lcout(iac_raw_buf_N_774),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1564638_i1_3_lut_LC_10_13_2.C_ON=1'b0;
    defparam i1564638_i1_3_lut_LC_10_13_2.SEQ_MODE=4'b0000;
    defparam i1564638_i1_3_lut_LC_10_13_2.LUT_INIT=16'b1110111001000100;
    LogicCell40 i1564638_i1_3_lut_LC_10_13_2 (
            .in0(N__47245),
            .in1(N__28494),
            .in2(_gnd_net_),
            .in3(N__28488),
            .lcout(n30_adj_1679),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_7_i26_3_lut_LC_10_13_3.C_ON=1'b0;
    defparam mux_128_Mux_7_i26_3_lut_LC_10_13_3.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_7_i26_3_lut_LC_10_13_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_128_Mux_7_i26_3_lut_LC_10_13_3 (
            .in0(N__28482),
            .in1(N__57205),
            .in2(_gnd_net_),
            .in3(N__28643),
            .lcout(),
            .ltout(n26_adj_1659_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18597_4_lut_LC_10_13_4.C_ON=1'b0;
    defparam i18597_4_lut_LC_10_13_4.SEQ_MODE=4'b0000;
    defparam i18597_4_lut_LC_10_13_4.LUT_INIT=16'b0101000011011000;
    LogicCell40 i18597_4_lut_LC_10_13_4 (
            .in0(N__46371),
            .in1(N__28467),
            .in2(N__28446),
            .in3(N__56900),
            .lcout(),
            .ltout(n21324_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_2__bdd_4_lut_19799_LC_10_13_5.C_ON=1'b0;
    defparam comm_cmd_2__bdd_4_lut_19799_LC_10_13_5.SEQ_MODE=4'b0000;
    defparam comm_cmd_2__bdd_4_lut_19799_LC_10_13_5.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_2__bdd_4_lut_19799_LC_10_13_5 (
            .in0(N__28365),
            .in1(N__47244),
            .in2(N__28443),
            .in3(N__47703),
            .lcout(n22401),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_7_i19_3_lut_LC_10_13_6.C_ON=1'b0;
    defparam mux_129_Mux_7_i19_3_lut_LC_10_13_6.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_7_i19_3_lut_LC_10_13_6.LUT_INIT=16'b1100110010101010;
    LogicCell40 mux_129_Mux_7_i19_3_lut_LC_10_13_6 (
            .in0(N__28433),
            .in1(N__28407),
            .in2(_gnd_net_),
            .in3(N__56898),
            .lcout(n19_adj_1621),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18596_4_lut_LC_10_13_7.C_ON=1'b0;
    defparam i18596_4_lut_LC_10_13_7.SEQ_MODE=4'b0000;
    defparam i18596_4_lut_LC_10_13_7.LUT_INIT=16'b0010001011110000;
    LogicCell40 i18596_4_lut_LC_10_13_7 (
            .in0(N__34494),
            .in1(N__57204),
            .in2(N__28377),
            .in3(N__46370),
            .lcout(n21323),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22371_bdd_4_lut_LC_10_14_0.C_ON=1'b0;
    defparam n22371_bdd_4_lut_LC_10_14_0.SEQ_MODE=4'b0000;
    defparam n22371_bdd_4_lut_LC_10_14_0.LUT_INIT=16'b1100110010111000;
    LogicCell40 n22371_bdd_4_lut_LC_10_14_0 (
            .in0(N__30889),
            .in1(N__28722),
            .in2(N__31299),
            .in3(N__46318),
            .lcout(n22374),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18_3_lut_LC_10_14_1.C_ON=1'b0;
    defparam i18_3_lut_LC_10_14_1.SEQ_MODE=4'b0000;
    defparam i18_3_lut_LC_10_14_1.LUT_INIT=16'b1110111001000100;
    LogicCell40 i18_3_lut_LC_10_14_1 (
            .in0(N__35874),
            .in1(N__35776),
            .in2(_gnd_net_),
            .in3(N__30968),
            .lcout(),
            .ltout(n12_adj_1454_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_trig_300_LC_10_14_2.C_ON=1'b0;
    defparam acadc_trig_300_LC_10_14_2.SEQ_MODE=4'b1000;
    defparam acadc_trig_300_LC_10_14_2.LUT_INIT=16'b1111111000000100;
    LogicCell40 acadc_trig_300_LC_10_14_2 (
            .in0(N__35733),
            .in1(N__28664),
            .in2(N__28716),
            .in3(N__28697),
            .lcout(acadc_trig),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVacadc_trig_300C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_209_LC_10_14_3.C_ON=1'b0;
    defparam i1_2_lut_adj_209_LC_10_14_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_209_LC_10_14_3.LUT_INIT=16'b0000000011001100;
    LogicCell40 i1_2_lut_adj_209_LC_10_14_3 (
            .in0(_gnd_net_),
            .in1(N__35859),
            .in2(_gnd_net_),
            .in3(N__35775),
            .lcout(n21053),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15227_2_lut_3_lut_LC_10_14_4.C_ON=1'b0;
    defparam i15227_2_lut_3_lut_LC_10_14_4.SEQ_MODE=4'b0000;
    defparam i15227_2_lut_3_lut_LC_10_14_4.LUT_INIT=16'b0010001010101010;
    LogicCell40 i15227_2_lut_3_lut_LC_10_14_4 (
            .in0(N__30966),
            .in1(N__28848),
            .in2(_gnd_net_),
            .in3(N__28806),
            .lcout(eis_state_2_N_392_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_adj_269_LC_10_14_5.C_ON=1'b0;
    defparam i2_3_lut_adj_269_LC_10_14_5.SEQ_MODE=4'b0000;
    defparam i2_3_lut_adj_269_LC_10_14_5.LUT_INIT=16'b0010001000000000;
    LogicCell40 i2_3_lut_adj_269_LC_10_14_5 (
            .in0(N__35873),
            .in1(N__28862),
            .in2(_gnd_net_),
            .in3(N__30908),
            .lcout(),
            .ltout(n21042_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_4_lut_adj_286_LC_10_14_6.C_ON=1'b0;
    defparam i1_4_lut_4_lut_adj_286_LC_10_14_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_4_lut_adj_286_LC_10_14_6.LUT_INIT=16'b1101000111110011;
    LogicCell40 i1_4_lut_4_lut_adj_286_LC_10_14_6 (
            .in0(N__30967),
            .in1(N__35800),
            .in2(N__28650),
            .in3(N__35875),
            .lcout(),
            .ltout(n21030_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_end_299_LC_10_14_7.C_ON=1'b0;
    defparam eis_end_299_LC_10_14_7.SEQ_MODE=4'b1000;
    defparam eis_end_299_LC_10_14_7.LUT_INIT=16'b1011101010001010;
    LogicCell40 eis_end_299_LC_10_14_7 (
            .in0(N__28644),
            .in1(N__35734),
            .in2(N__28647),
            .in3(N__35777),
            .lcout(eis_end),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVacadc_trig_300C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_state_1__bdd_4_lut_19731_4_lut_LC_10_15_0.C_ON=1'b0;
    defparam eis_state_1__bdd_4_lut_19731_4_lut_LC_10_15_0.SEQ_MODE=4'b0000;
    defparam eis_state_1__bdd_4_lut_19731_4_lut_LC_10_15_0.LUT_INIT=16'b0110111000101010;
    LogicCell40 eis_state_1__bdd_4_lut_19731_4_lut_LC_10_15_0 (
            .in0(N__35866),
            .in1(N__35783),
            .in2(N__30981),
            .in3(N__28764),
            .lcout(n22437),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19465_3_lut_4_lut_LC_10_15_1.C_ON=1'b0;
    defparam i19465_3_lut_4_lut_LC_10_15_1.SEQ_MODE=4'b0000;
    defparam i19465_3_lut_4_lut_LC_10_15_1.LUT_INIT=16'b0000000000010101;
    LogicCell40 i19465_3_lut_4_lut_LC_10_15_1 (
            .in0(N__35860),
            .in1(N__30955),
            .in2(N__35794),
            .in3(N__35707),
            .lcout(n11989),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i24_4_lut_LC_10_15_2.C_ON=1'b0;
    defparam i24_4_lut_LC_10_15_2.SEQ_MODE=4'b0000;
    defparam i24_4_lut_LC_10_15_2.LUT_INIT=16'b1110111111100000;
    LogicCell40 i24_4_lut_LC_10_15_2 (
            .in0(N__31029),
            .in1(N__43043),
            .in2(N__30980),
            .in3(N__28863),
            .lcout(),
            .ltout(n11_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19423_3_lut_LC_10_15_3.C_ON=1'b0;
    defparam i19423_3_lut_LC_10_15_3.SEQ_MODE=4'b0000;
    defparam i19423_3_lut_LC_10_15_3.LUT_INIT=16'b0101111111111111;
    LogicCell40 i19423_3_lut_LC_10_15_3 (
            .in0(N__35782),
            .in1(_gnd_net_),
            .in2(N__28851),
            .in3(N__35865),
            .lcout(n11908),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_4_lut_adj_270_LC_10_15_4.C_ON=1'b0;
    defparam i2_4_lut_4_lut_adj_270_LC_10_15_4.SEQ_MODE=4'b0000;
    defparam i2_4_lut_4_lut_adj_270_LC_10_15_4.LUT_INIT=16'b0000000001000101;
    LogicCell40 i2_4_lut_4_lut_adj_270_LC_10_15_4 (
            .in0(N__35708),
            .in1(N__30964),
            .in2(N__35876),
            .in3(N__35781),
            .lcout(n11933),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15247_2_lut_3_lut_LC_10_15_5.C_ON=1'b0;
    defparam i15247_2_lut_3_lut_LC_10_15_5.SEQ_MODE=4'b0000;
    defparam i15247_2_lut_3_lut_LC_10_15_5.LUT_INIT=16'b1110111010101010;
    LogicCell40 i15247_2_lut_3_lut_LC_10_15_5 (
            .in0(N__35861),
            .in1(N__28847),
            .in2(_gnd_net_),
            .in3(N__28802),
            .lcout(eis_state_2_N_392_1),
            .ltout(eis_state_2_N_392_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_state_2__I_0_371_Mux_1_i2_4_lut_LC_10_15_6.C_ON=1'b0;
    defparam eis_state_2__I_0_371_Mux_1_i2_4_lut_LC_10_15_6.SEQ_MODE=4'b0000;
    defparam eis_state_2__I_0_371_Mux_1_i2_4_lut_LC_10_15_6.LUT_INIT=16'b1100000011100010;
    LogicCell40 eis_state_2__I_0_371_Mux_1_i2_4_lut_LC_10_15_6 (
            .in0(N__31030),
            .in1(N__30965),
            .in2(N__28758),
            .in3(N__32815),
            .lcout(),
            .ltout(n2_adj_1696_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_state_i1_LC_10_15_7.C_ON=1'b0;
    defparam eis_state_i1_LC_10_15_7.SEQ_MODE=4'b1010;
    defparam eis_state_i1_LC_10_15_7.LUT_INIT=16'b1111101001000100;
    LogicCell40 eis_state_i1_LC_10_15_7 (
            .in0(N__35784),
            .in1(N__30962),
            .in2(N__28755),
            .in3(N__28752),
            .lcout(eis_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVeis_state_i1C_net),
            .ce(N__30995),
            .sr(N__35735));
    defparam \ADC_IAC.ADC_DATA_i15_LC_10_16_1 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i15_LC_10_16_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i15_LC_10_16_1 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_IAC.ADC_DATA_i15_LC_10_16_1  (
            .in0(N__38737),
            .in1(N__38551),
            .in2(N__42046),
            .in3(N__28746),
            .lcout(buf_adcdata_iac_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56034),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i9_LC_10_16_2.C_ON=1'b0;
    defparam acadc_skipCount_i9_LC_10_16_2.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i9_LC_10_16_2.LUT_INIT=16'b0111001101000000;
    LogicCell40 acadc_skipCount_i9_LC_10_16_2 (
            .in0(N__49302),
            .in1(N__47863),
            .in2(N__53466),
            .in3(N__42977),
            .lcout(acadc_skipCount_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56034),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i12_LC_10_16_4.C_ON=1'b0;
    defparam buf_dds0_i12_LC_10_16_4.SEQ_MODE=4'b1000;
    defparam buf_dds0_i12_LC_10_16_4.LUT_INIT=16'b0101000011001100;
    LogicCell40 buf_dds0_i12_LC_10_16_4 (
            .in0(N__49303),
            .in1(N__36256),
            .in2(N__47820),
            .in3(N__41665),
            .lcout(buf_dds0_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56034),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i8_LC_10_16_5.C_ON=1'b0;
    defparam buf_device_acadc_i8_LC_10_16_5.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i8_LC_10_16_5.LUT_INIT=16'b0011101100001000;
    LogicCell40 buf_device_acadc_i8_LC_10_16_5 (
            .in0(N__42543),
            .in1(N__39516),
            .in2(N__49382),
            .in3(N__28990),
            .lcout(VAC_FLT1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56034),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i15_LC_10_16_6.C_ON=1'b0;
    defparam acadc_skipCount_i15_LC_10_16_6.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i15_LC_10_16_6.LUT_INIT=16'b0111010000110000;
    LogicCell40 acadc_skipCount_i15_LC_10_16_6 (
            .in0(N__49301),
            .in1(N__47862),
            .in2(N__31185),
            .in3(N__42542),
            .lcout(acadc_skipCount_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56034),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i21_LC_10_16_7 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i21_LC_10_16_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i21_LC_10_16_7 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i21_LC_10_16_7  (
            .in0(N__38738),
            .in1(N__38552),
            .in2(N__28971),
            .in3(N__28933),
            .lcout(buf_adcdata_iac_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56034),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i20_LC_10_17_0 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i20_LC_10_17_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i20_LC_10_17_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i20_LC_10_17_0  (
            .in0(N__38746),
            .in1(N__38504),
            .in2(N__28911),
            .in3(N__32128),
            .lcout(buf_adcdata_iac_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56050),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i3_LC_10_17_2.C_ON=1'b0;
    defparam buf_device_acadc_i3_LC_10_17_2.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i3_LC_10_17_2.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_device_acadc_i3_LC_10_17_2 (
            .in0(N__49337),
            .in1(N__39528),
            .in2(N__45878),
            .in3(N__30526),
            .lcout(IAC_FLT0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56050),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i12_LC_10_17_3 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i12_LC_10_17_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i12_LC_10_17_3 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i12_LC_10_17_3  (
            .in0(N__38503),
            .in1(N__38745),
            .in2(N__29430),
            .in3(N__30601),
            .lcout(buf_adcdata_iac_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56050),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i11_LC_10_17_5.C_ON=1'b0;
    defparam buf_dds0_i11_LC_10_17_5.SEQ_MODE=4'b1000;
    defparam buf_dds0_i11_LC_10_17_5.LUT_INIT=16'b0101000011001100;
    LogicCell40 buf_dds0_i11_LC_10_17_5 (
            .in0(N__49336),
            .in1(N__31367),
            .in2(N__45356),
            .in3(N__41667),
            .lcout(buf_dds0_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56050),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i8_LC_10_17_7.C_ON=1'b0;
    defparam acadc_skipCount_i8_LC_10_17_7.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i8_LC_10_17_7.LUT_INIT=16'b0111001101000000;
    LogicCell40 acadc_skipCount_i8_LC_10_17_7 (
            .in0(N__49335),
            .in1(N__47864),
            .in2(N__45646),
            .in3(N__32719),
            .lcout(acadc_skipCount_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56050),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i26_LC_10_18_3 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i26_LC_10_18_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i26_LC_10_18_3 .LUT_INIT=16'b1110010001000100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i26_LC_10_18_3  (
            .in0(N__29364),
            .in1(N__32779),
            .in2(N__28886),
            .in3(N__38597),
            .lcout(cmd_rdadctmp_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56064),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.cmd_rdadctmp_i21_LC_10_18_6 .C_ON=1'b0;
    defparam \ADC_IAC.cmd_rdadctmp_i21_LC_10_18_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.cmd_rdadctmp_i21_LC_10_18_6 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \ADC_IAC.cmd_rdadctmp_i21_LC_10_18_6  (
            .in0(N__38595),
            .in1(N__33097),
            .in2(N__29428),
            .in3(N__29365),
            .lcout(cmd_rdadctmp_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56064),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i23_LC_10_18_7 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i23_LC_10_18_7 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i23_LC_10_18_7 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i23_LC_10_18_7  (
            .in0(N__38744),
            .in1(N__38596),
            .in2(N__29217),
            .in3(N__29188),
            .lcout(buf_adcdata_iac_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56064),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.adc_state_i2_LC_11_3_0 .C_ON=1'b0;
    defparam \ADC_VDC.adc_state_i2_LC_11_3_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.adc_state_i2_LC_11_3_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ADC_VDC.adc_state_i2_LC_11_3_0  (
            .in0(N__51867),
            .in1(N__51344),
            .in2(_gnd_net_),
            .in3(N__51180),
            .lcout(adc_state_2_adj_1500),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42364),
            .ce(N__29166),
            .sr(N__31383));
    defparam \ADC_VDC.i19237_4_lut_LC_11_4_0 .C_ON=1'b0;
    defparam \ADC_VDC.i19237_4_lut_LC_11_4_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i19237_4_lut_LC_11_4_0 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \ADC_VDC.i19237_4_lut_LC_11_4_0  (
            .in0(N__34374),
            .in1(N__34338),
            .in2(N__34440),
            .in3(N__34401),
            .lcout(),
            .ltout(\ADC_VDC.n21593_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i19248_4_lut_LC_11_4_1 .C_ON=1'b0;
    defparam \ADC_VDC.i19248_4_lut_LC_11_4_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i19248_4_lut_LC_11_4_1 .LUT_INIT=16'b1010100010001000;
    LogicCell40 \ADC_VDC.i19248_4_lut_LC_11_4_1  (
            .in0(N__51892),
            .in1(N__31680),
            .in2(N__29154),
            .in3(N__34305),
            .lcout(),
            .ltout(\ADC_VDC.n21590_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.n22587_bdd_4_lut_4_lut_LC_11_4_2 .C_ON=1'b0;
    defparam \ADC_VDC.n22587_bdd_4_lut_4_lut_LC_11_4_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.n22587_bdd_4_lut_4_lut_LC_11_4_2 .LUT_INIT=16'b1011101101010000;
    LogicCell40 \ADC_VDC.n22587_bdd_4_lut_4_lut_LC_11_4_2  (
            .in0(N__51356),
            .in1(N__51893),
            .in2(N__29151),
            .in3(N__30291),
            .lcout(\ADC_VDC.n22590 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_3_lut_4_lut_adj_34_LC_11_4_3 .C_ON=1'b0;
    defparam \ADC_VDC.i1_3_lut_4_lut_adj_34_LC_11_4_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_3_lut_4_lut_adj_34_LC_11_4_3 .LUT_INIT=16'b1100110001000000;
    LogicCell40 \ADC_VDC.i1_3_lut_4_lut_adj_34_LC_11_4_3  (
            .in0(N__51151),
            .in1(N__51355),
            .in2(N__51909),
            .in3(N__51711),
            .lcout(n13324),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i24_3_lut_4_lut_LC_11_4_4 .C_ON=1'b0;
    defparam \ADC_VDC.i24_3_lut_4_lut_LC_11_4_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i24_3_lut_4_lut_LC_11_4_4 .LUT_INIT=16'b0011010100110000;
    LogicCell40 \ADC_VDC.i24_3_lut_4_lut_LC_11_4_4  (
            .in0(N__51710),
            .in1(N__51149),
            .in2(N__51414),
            .in3(N__51986),
            .lcout(\ADC_VDC.n11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_2_lut_LC_11_4_5 .C_ON=1'b0;
    defparam \ADC_VDC.i1_2_lut_LC_11_4_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_2_lut_LC_11_4_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ADC_VDC.i1_2_lut_LC_11_4_5  (
            .in0(_gnd_net_),
            .in1(N__51357),
            .in2(_gnd_net_),
            .in3(N__51713),
            .lcout(\ADC_VDC.n5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i16264_3_lut_LC_11_4_6 .C_ON=1'b0;
    defparam \ADC_VDC.i16264_3_lut_LC_11_4_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i16264_3_lut_LC_11_4_6 .LUT_INIT=16'b1110111001100110;
    LogicCell40 \ADC_VDC.i16264_3_lut_LC_11_4_6  (
            .in0(N__51856),
            .in1(N__51985),
            .in2(_gnd_net_),
            .in3(N__51150),
            .lcout(),
            .ltout(\ADC_VDC.n7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_4_lut_adj_32_LC_11_4_7 .C_ON=1'b0;
    defparam \ADC_VDC.i1_4_lut_adj_32_LC_11_4_7 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_4_lut_adj_32_LC_11_4_7 .LUT_INIT=16'b1011101011111110;
    LogicCell40 \ADC_VDC.i1_4_lut_adj_32_LC_11_4_7  (
            .in0(N__51442),
            .in1(N__51712),
            .in2(N__29691),
            .in3(N__29686),
            .lcout(\ADC_VDC.n65 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i8_LC_11_5_0 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i8_LC_11_5_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i8_LC_11_5_0 .LUT_INIT=16'b0010111000100010;
    LogicCell40 \ADC_VDC.ADC_DATA_i8_LC_11_5_0  (
            .in0(N__43769),
            .in1(N__31601),
            .in2(N__51491),
            .in3(N__29670),
            .lcout(buf_adcdata_vdc_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42305),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i13_LC_11_5_1 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i13_LC_11_5_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i13_LC_11_5_1 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \ADC_VDC.ADC_DATA_i13_LC_11_5_1  (
            .in0(N__51361),
            .in1(N__29621),
            .in2(N__31617),
            .in3(N__29649),
            .lcout(buf_adcdata_vdc_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42305),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i19_LC_11_5_2 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i19_LC_11_5_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i19_LC_11_5_2 .LUT_INIT=16'b0010111000100010;
    LogicCell40 \ADC_VDC.ADC_DATA_i19_LC_11_5_2  (
            .in0(N__29582),
            .in1(N__31600),
            .in2(N__51490),
            .in3(N__29610),
            .lcout(buf_adcdata_vdc_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42305),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i17_LC_11_5_3 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i17_LC_11_5_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i17_LC_11_5_3 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \ADC_VDC.ADC_DATA_i17_LC_11_5_3  (
            .in0(N__51362),
            .in1(N__29540),
            .in2(N__31618),
            .in3(N__29571),
            .lcout(buf_adcdata_vdc_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42305),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i21_LC_11_5_4 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i21_LC_11_5_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i21_LC_11_5_4 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \ADC_VDC.ADC_DATA_i21_LC_11_5_4  (
            .in0(N__29529),
            .in1(N__31590),
            .in2(N__29501),
            .in3(N__51364),
            .lcout(buf_adcdata_vdc_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42305),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i20_LC_11_5_5 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i20_LC_11_5_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i20_LC_11_5_5 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \ADC_VDC.ADC_DATA_i20_LC_11_5_5  (
            .in0(N__51363),
            .in1(N__31895),
            .in2(N__31619),
            .in3(N__29484),
            .lcout(buf_adcdata_vdc_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42305),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_4_i16_3_lut_LC_11_5_6.C_ON=1'b0;
    defparam mux_129_Mux_4_i16_3_lut_LC_11_5_6.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_4_i16_3_lut_LC_11_5_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_129_Mux_4_i16_3_lut_LC_11_5_6 (
            .in0(N__29463),
            .in1(N__32255),
            .in2(_gnd_net_),
            .in3(N__57208),
            .lcout(n16_adj_1633),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.adc_state_1__bdd_4_lut_4_lut_LC_11_5_7 .C_ON=1'b0;
    defparam \ADC_VDC.adc_state_1__bdd_4_lut_4_lut_LC_11_5_7 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.adc_state_1__bdd_4_lut_4_lut_LC_11_5_7 .LUT_INIT=16'b0010110001101100;
    LogicCell40 \ADC_VDC.adc_state_1__bdd_4_lut_4_lut_LC_11_5_7  (
            .in0(N__51860),
            .in1(N__51175),
            .in2(N__51415),
            .in3(N__30285),
            .lcout(\ADC_VDC.n22587 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i3_4_lut_adj_30_LC_11_6_1 .C_ON=1'b0;
    defparam \ADC_VDC.i3_4_lut_adj_30_LC_11_6_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i3_4_lut_adj_30_LC_11_6_1 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \ADC_VDC.i3_4_lut_adj_30_LC_11_6_1  (
            .in0(N__34369),
            .in1(N__31470),
            .in2(N__34436),
            .in3(N__31671),
            .lcout(\ADC_VDC.n10708 ),
            .ltout(\ADC_VDC.n10708_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.cmd_rdadctmp_i23_LC_11_6_2 .C_ON=1'b0;
    defparam \ADC_VDC.cmd_rdadctmp_i23_LC_11_6_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.cmd_rdadctmp_i23_LC_11_6_2 .LUT_INIT=16'b1010010111001100;
    LogicCell40 \ADC_VDC.cmd_rdadctmp_i23_LC_11_6_2  (
            .in0(N__30236),
            .in1(N__30278),
            .in2(N__30246),
            .in3(N__51203),
            .lcout(\ADC_VDC.cmd_rdadctmp_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42414),
            .ce(N__31941),
            .sr(N__30222));
    defparam \ADC_VDC.i8_4_lut_LC_11_6_3 .C_ON=1'b0;
    defparam \ADC_VDC.i8_4_lut_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i8_4_lut_LC_11_6_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.i8_4_lut_LC_11_6_3  (
            .in0(N__30209),
            .in1(N__30197),
            .in2(N__30186),
            .in3(N__30170),
            .lcout(\ADC_VDC.n20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.i19393_4_lut_LC_11_6_4 .C_ON=1'b0;
    defparam \CLK_DDS.i19393_4_lut_LC_11_6_4 .SEQ_MODE=4'b0000;
    defparam \CLK_DDS.i19393_4_lut_LC_11_6_4 .LUT_INIT=16'b1010101000100110;
    LogicCell40 \CLK_DDS.i19393_4_lut_LC_11_6_4  (
            .in0(N__30072),
            .in1(N__29947),
            .in2(N__38828),
            .in3(N__29792),
            .lcout(\CLK_DDS.n13005 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.i23_4_lut_LC_11_6_5 .C_ON=1'b0;
    defparam \CLK_DDS.i23_4_lut_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \CLK_DDS.i23_4_lut_LC_11_6_5 .LUT_INIT=16'b1111101000010101;
    LogicCell40 \CLK_DDS.i23_4_lut_LC_11_6_5  (
            .in0(N__29794),
            .in1(N__38824),
            .in2(N__29952),
            .in3(N__30074),
            .lcout(\CLK_DDS.n9_adj_1433 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \CLK_DDS.i19409_4_lut_LC_11_6_6 .C_ON=1'b0;
    defparam \CLK_DDS.i19409_4_lut_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \CLK_DDS.i19409_4_lut_LC_11_6_6 .LUT_INIT=16'b1111111110111110;
    LogicCell40 \CLK_DDS.i19409_4_lut_LC_11_6_6  (
            .in0(N__30073),
            .in1(N__29946),
            .in2(N__38829),
            .in3(N__29793),
            .lcout(\CLK_DDS.n9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam secclk_cnt_3765_3766__i1_LC_11_7_0.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i1_LC_11_7_0.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i1_LC_11_7_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i1_LC_11_7_0 (
            .in0(_gnd_net_),
            .in1(N__34554),
            .in2(_gnd_net_),
            .in3(N__29694),
            .lcout(secclk_cnt_0),
            .ltout(),
            .carryin(bfn_11_7_0_),
            .carryout(n19956),
            .clk(N__50782),
            .ce(),
            .sr(N__34714));
    defparam secclk_cnt_3765_3766__i2_LC_11_7_1.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i2_LC_11_7_1.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i2_LC_11_7_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i2_LC_11_7_1 (
            .in0(_gnd_net_),
            .in1(N__34610),
            .in2(_gnd_net_),
            .in3(N__30318),
            .lcout(secclk_cnt_1),
            .ltout(),
            .carryin(n19956),
            .carryout(n19957),
            .clk(N__50782),
            .ce(),
            .sr(N__34714));
    defparam secclk_cnt_3765_3766__i3_LC_11_7_2.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i3_LC_11_7_2.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i3_LC_11_7_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i3_LC_11_7_2 (
            .in0(_gnd_net_),
            .in1(N__31785),
            .in2(_gnd_net_),
            .in3(N__30315),
            .lcout(secclk_cnt_2),
            .ltout(),
            .carryin(n19957),
            .carryout(n19958),
            .clk(N__50782),
            .ce(),
            .sr(N__34714));
    defparam secclk_cnt_3765_3766__i4_LC_11_7_3.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i4_LC_11_7_3.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i4_LC_11_7_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i4_LC_11_7_3 (
            .in0(_gnd_net_),
            .in1(N__31803),
            .in2(_gnd_net_),
            .in3(N__30312),
            .lcout(secclk_cnt_3),
            .ltout(),
            .carryin(n19958),
            .carryout(n19959),
            .clk(N__50782),
            .ce(),
            .sr(N__34714));
    defparam secclk_cnt_3765_3766__i5_LC_11_7_4.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i5_LC_11_7_4.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i5_LC_11_7_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i5_LC_11_7_4 (
            .in0(_gnd_net_),
            .in1(N__34517),
            .in2(_gnd_net_),
            .in3(N__30309),
            .lcout(secclk_cnt_4),
            .ltout(),
            .carryin(n19959),
            .carryout(n19960),
            .clk(N__50782),
            .ce(),
            .sr(N__34714));
    defparam secclk_cnt_3765_3766__i6_LC_11_7_5.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i6_LC_11_7_5.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i6_LC_11_7_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i6_LC_11_7_5 (
            .in0(_gnd_net_),
            .in1(N__34592),
            .in2(_gnd_net_),
            .in3(N__30306),
            .lcout(secclk_cnt_5),
            .ltout(),
            .carryin(n19960),
            .carryout(n19961),
            .clk(N__50782),
            .ce(),
            .sr(N__34714));
    defparam secclk_cnt_3765_3766__i7_LC_11_7_6.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i7_LC_11_7_6.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i7_LC_11_7_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i7_LC_11_7_6 (
            .in0(_gnd_net_),
            .in1(N__31845),
            .in2(_gnd_net_),
            .in3(N__30303),
            .lcout(secclk_cnt_6),
            .ltout(),
            .carryin(n19961),
            .carryout(n19962),
            .clk(N__50782),
            .ce(),
            .sr(N__34714));
    defparam secclk_cnt_3765_3766__i8_LC_11_7_7.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i8_LC_11_7_7.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i8_LC_11_7_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i8_LC_11_7_7 (
            .in0(_gnd_net_),
            .in1(N__31760),
            .in2(_gnd_net_),
            .in3(N__30300),
            .lcout(secclk_cnt_7),
            .ltout(),
            .carryin(n19962),
            .carryout(n19963),
            .clk(N__50782),
            .ce(),
            .sr(N__34714));
    defparam secclk_cnt_3765_3766__i9_LC_11_8_0.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i9_LC_11_8_0.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i9_LC_11_8_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i9_LC_11_8_0 (
            .in0(_gnd_net_),
            .in1(N__34625),
            .in2(_gnd_net_),
            .in3(N__30297),
            .lcout(secclk_cnt_8),
            .ltout(),
            .carryin(bfn_11_8_0_),
            .carryout(n19964),
            .clk(N__50786),
            .ce(),
            .sr(N__34716));
    defparam secclk_cnt_3765_3766__i10_LC_11_8_1.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i10_LC_11_8_1.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i10_LC_11_8_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i10_LC_11_8_1 (
            .in0(_gnd_net_),
            .in1(N__35144),
            .in2(_gnd_net_),
            .in3(N__30294),
            .lcout(secclk_cnt_9),
            .ltout(),
            .carryin(n19964),
            .carryout(n19965),
            .clk(N__50786),
            .ce(),
            .sr(N__34716));
    defparam secclk_cnt_3765_3766__i11_LC_11_8_2.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i11_LC_11_8_2.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i11_LC_11_8_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i11_LC_11_8_2 (
            .in0(_gnd_net_),
            .in1(N__31817),
            .in2(_gnd_net_),
            .in3(N__30345),
            .lcout(secclk_cnt_10),
            .ltout(),
            .carryin(n19965),
            .carryout(n19966),
            .clk(N__50786),
            .ce(),
            .sr(N__34716));
    defparam secclk_cnt_3765_3766__i12_LC_11_8_3.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i12_LC_11_8_3.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i12_LC_11_8_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i12_LC_11_8_3 (
            .in0(_gnd_net_),
            .in1(N__34532),
            .in2(_gnd_net_),
            .in3(N__30342),
            .lcout(secclk_cnt_11),
            .ltout(),
            .carryin(n19966),
            .carryout(n19967),
            .clk(N__50786),
            .ce(),
            .sr(N__34716));
    defparam secclk_cnt_3765_3766__i13_LC_11_8_4.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i13_LC_11_8_4.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i13_LC_11_8_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i13_LC_11_8_4 (
            .in0(_gnd_net_),
            .in1(N__30392),
            .in2(_gnd_net_),
            .in3(N__30339),
            .lcout(secclk_cnt_12),
            .ltout(),
            .carryin(n19967),
            .carryout(n19968),
            .clk(N__50786),
            .ce(),
            .sr(N__34716));
    defparam secclk_cnt_3765_3766__i14_LC_11_8_5.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i14_LC_11_8_5.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i14_LC_11_8_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i14_LC_11_8_5 (
            .in0(_gnd_net_),
            .in1(N__31773),
            .in2(_gnd_net_),
            .in3(N__30336),
            .lcout(secclk_cnt_13),
            .ltout(),
            .carryin(n19968),
            .carryout(n19969),
            .clk(N__50786),
            .ce(),
            .sr(N__34716));
    defparam secclk_cnt_3765_3766__i15_LC_11_8_6.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i15_LC_11_8_6.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i15_LC_11_8_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i15_LC_11_8_6 (
            .in0(_gnd_net_),
            .in1(N__31833),
            .in2(_gnd_net_),
            .in3(N__30333),
            .lcout(secclk_cnt_14),
            .ltout(),
            .carryin(n19969),
            .carryout(n19970),
            .clk(N__50786),
            .ce(),
            .sr(N__34716));
    defparam secclk_cnt_3765_3766__i16_LC_11_8_7.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i16_LC_11_8_7.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i16_LC_11_8_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i16_LC_11_8_7 (
            .in0(_gnd_net_),
            .in1(N__34643),
            .in2(_gnd_net_),
            .in3(N__30330),
            .lcout(secclk_cnt_15),
            .ltout(),
            .carryin(n19970),
            .carryout(n19971),
            .clk(N__50786),
            .ce(),
            .sr(N__34716));
    defparam secclk_cnt_3765_3766__i17_LC_11_9_0.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i17_LC_11_9_0.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i17_LC_11_9_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i17_LC_11_9_0 (
            .in0(_gnd_net_),
            .in1(N__31746),
            .in2(_gnd_net_),
            .in3(N__30327),
            .lcout(secclk_cnt_16),
            .ltout(),
            .carryin(bfn_11_9_0_),
            .carryout(n19972),
            .clk(N__50788),
            .ce(),
            .sr(N__34715));
    defparam secclk_cnt_3765_3766__i18_LC_11_9_1.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i18_LC_11_9_1.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i18_LC_11_9_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i18_LC_11_9_1 (
            .in0(_gnd_net_),
            .in1(N__35129),
            .in2(_gnd_net_),
            .in3(N__30324),
            .lcout(secclk_cnt_17),
            .ltout(),
            .carryin(n19972),
            .carryout(n19973),
            .clk(N__50788),
            .ce(),
            .sr(N__34715));
    defparam secclk_cnt_3765_3766__i19_LC_11_9_2.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i19_LC_11_9_2.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i19_LC_11_9_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i19_LC_11_9_2 (
            .in0(_gnd_net_),
            .in1(N__34571),
            .in2(_gnd_net_),
            .in3(N__30321),
            .lcout(secclk_cnt_18),
            .ltout(),
            .carryin(n19973),
            .carryout(n19974),
            .clk(N__50788),
            .ce(),
            .sr(N__34715));
    defparam secclk_cnt_3765_3766__i20_LC_11_9_3.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i20_LC_11_9_3.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i20_LC_11_9_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i20_LC_11_9_3 (
            .in0(_gnd_net_),
            .in1(N__30408),
            .in2(_gnd_net_),
            .in3(N__30435),
            .lcout(secclk_cnt_19),
            .ltout(),
            .carryin(n19974),
            .carryout(n19975),
            .clk(N__50788),
            .ce(),
            .sr(N__34715));
    defparam secclk_cnt_3765_3766__i21_LC_11_9_4.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i21_LC_11_9_4.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i21_LC_11_9_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i21_LC_11_9_4 (
            .in0(_gnd_net_),
            .in1(N__31928),
            .in2(_gnd_net_),
            .in3(N__30432),
            .lcout(secclk_cnt_20),
            .ltout(),
            .carryin(n19975),
            .carryout(n19976),
            .clk(N__50788),
            .ce(),
            .sr(N__34715));
    defparam secclk_cnt_3765_3766__i22_LC_11_9_5.C_ON=1'b1;
    defparam secclk_cnt_3765_3766__i22_LC_11_9_5.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i22_LC_11_9_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i22_LC_11_9_5 (
            .in0(_gnd_net_),
            .in1(N__30422),
            .in2(_gnd_net_),
            .in3(N__30429),
            .lcout(secclk_cnt_21),
            .ltout(),
            .carryin(n19976),
            .carryout(n19977),
            .clk(N__50788),
            .ce(),
            .sr(N__34715));
    defparam secclk_cnt_3765_3766__i23_LC_11_9_6.C_ON=1'b0;
    defparam secclk_cnt_3765_3766__i23_LC_11_9_6.SEQ_MODE=4'b1000;
    defparam secclk_cnt_3765_3766__i23_LC_11_9_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 secclk_cnt_3765_3766__i23_LC_11_9_6 (
            .in0(_gnd_net_),
            .in1(N__30378),
            .in2(_gnd_net_),
            .in3(N__30426),
            .lcout(secclk_cnt_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50788),
            .ce(),
            .sr(N__34715));
    defparam i6_4_lut_adj_201_LC_11_10_0.C_ON=1'b0;
    defparam i6_4_lut_adj_201_LC_11_10_0.SEQ_MODE=4'b0000;
    defparam i6_4_lut_adj_201_LC_11_10_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 i6_4_lut_adj_201_LC_11_10_0 (
            .in0(N__30423),
            .in1(N__30407),
            .in2(N__30396),
            .in3(N__30377),
            .lcout(n14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6751_2_lut_LC_11_10_1.C_ON=1'b0;
    defparam i6751_2_lut_LC_11_10_1.SEQ_MODE=4'b0000;
    defparam i6751_2_lut_LC_11_10_1.LUT_INIT=16'b0011001100000000;
    LogicCell40 i6751_2_lut_LC_11_10_1 (
            .in0(_gnd_net_),
            .in1(N__54500),
            .in2(_gnd_net_),
            .in3(N__54001),
            .lcout(n9269),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i11_LC_11_10_2.C_ON=1'b0;
    defparam acadc_skipCount_i11_LC_11_10_2.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i11_LC_11_10_2.LUT_INIT=16'b0111010000110000;
    LogicCell40 acadc_skipCount_i11_LC_11_10_2 (
            .in0(N__49350),
            .in1(N__47923),
            .in2(N__32562),
            .in3(N__45335),
            .lcout(acadc_skipCount_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55953),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i14_LC_11_10_3.C_ON=1'b0;
    defparam acadc_skipCount_i14_LC_11_10_3.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i14_LC_11_10_3.LUT_INIT=16'b0111010100100000;
    LogicCell40 acadc_skipCount_i14_LC_11_10_3 (
            .in0(N__47924),
            .in1(N__49351),
            .in2(N__49586),
            .in3(N__32217),
            .lcout(acadc_skipCount_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55953),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i8_LC_11_10_4.C_ON=1'b0;
    defparam req_data_cnt_i8_LC_11_10_4.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i8_LC_11_10_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 req_data_cnt_i8_LC_11_10_4 (
            .in0(N__35561),
            .in1(N__40447),
            .in2(_gnd_net_),
            .in3(N__30841),
            .lcout(req_data_cnt_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55953),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i14_LC_11_10_5.C_ON=1'b0;
    defparam req_data_cnt_i14_LC_11_10_5.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i14_LC_11_10_5.LUT_INIT=16'b1100110010101010;
    LogicCell40 req_data_cnt_i14_LC_11_10_5 (
            .in0(N__31991),
            .in1(N__30366),
            .in2(_gnd_net_),
            .in3(N__35560),
            .lcout(req_data_cnt_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55953),
            .ce(),
            .sr(_gnd_net_));
    defparam i18602_4_lut_LC_11_10_6.C_ON=1'b0;
    defparam i18602_4_lut_LC_11_10_6.SEQ_MODE=4'b0000;
    defparam i18602_4_lut_LC_11_10_6.LUT_INIT=16'b0111001001010000;
    LogicCell40 i18602_4_lut_LC_11_10_6 (
            .in0(N__46455),
            .in1(N__56865),
            .in2(N__32226),
            .in3(N__31990),
            .lcout(n21329),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_2_i17_3_lut_LC_11_10_7.C_ON=1'b0;
    defparam mux_128_Mux_2_i17_3_lut_LC_11_10_7.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_2_i17_3_lut_LC_11_10_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_128_Mux_2_i17_3_lut_LC_11_10_7 (
            .in0(N__56866),
            .in1(N__32756),
            .in2(_gnd_net_),
            .in3(N__30542),
            .lcout(n17_adj_1682),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_310_LC_11_11_0.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_310_LC_11_11_0.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_310_LC_11_11_0.LUT_INIT=16'b1101110111111111;
    LogicCell40 i1_2_lut_3_lut_adj_310_LC_11_11_0 (
            .in0(N__56751),
            .in1(N__37572),
            .in2(_gnd_net_),
            .in3(N__47133),
            .lcout(n11570),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22401_bdd_4_lut_LC_11_11_1.C_ON=1'b0;
    defparam n22401_bdd_4_lut_LC_11_11_1.SEQ_MODE=4'b0000;
    defparam n22401_bdd_4_lut_LC_11_11_1.LUT_INIT=16'b1111101001000100;
    LogicCell40 n22401_bdd_4_lut_LC_11_11_1 (
            .in0(N__47136),
            .in1(N__30507),
            .in2(N__30498),
            .in3(N__30486),
            .lcout(n22404),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i15_LC_11_11_2.C_ON=1'b0;
    defparam buf_dds0_i15_LC_11_11_2.SEQ_MODE=4'b1000;
    defparam buf_dds0_i15_LC_11_11_2.LUT_INIT=16'b0010001011110000;
    LogicCell40 buf_dds0_i15_LC_11_11_2 (
            .in0(N__42535),
            .in1(N__49325),
            .in2(N__31294),
            .in3(N__41668),
            .lcout(buf_dds0_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55957),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_278_LC_11_11_3.C_ON=1'b0;
    defparam i1_3_lut_adj_278_LC_11_11_3.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_278_LC_11_11_3.LUT_INIT=16'b1111111111111010;
    LogicCell40 i1_3_lut_adj_278_LC_11_11_3 (
            .in0(N__47134),
            .in1(_gnd_net_),
            .in2(N__37582),
            .in3(N__54007),
            .lcout(n21122),
            .ltout(n21122_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_276_LC_11_11_4.C_ON=1'b0;
    defparam i1_4_lut_adj_276_LC_11_11_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_276_LC_11_11_4.LUT_INIT=16'b1100110100000000;
    LogicCell40 i1_4_lut_adj_276_LC_11_11_4 (
            .in0(N__32637),
            .in1(N__49323),
            .in2(N__30465),
            .in3(N__55296),
            .lcout(n12610),
            .ltout(n12610_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i5_LC_11_11_5.C_ON=1'b0;
    defparam buf_device_acadc_i5_LC_11_11_5.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i5_LC_11_11_5.LUT_INIT=16'b0100111101000000;
    LogicCell40 buf_device_acadc_i5_LC_11_11_5 (
            .in0(N__49324),
            .in1(N__47787),
            .in2(N__30462),
            .in3(N__32090),
            .lcout(VAC_OSR0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55957),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_5_i30_3_lut_LC_11_11_6.C_ON=1'b0;
    defparam mux_130_Mux_5_i30_3_lut_LC_11_11_6.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_5_i30_3_lut_LC_11_11_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_130_Mux_5_i30_3_lut_LC_11_11_6 (
            .in0(N__30459),
            .in1(N__30444),
            .in2(_gnd_net_),
            .in3(N__47135),
            .lcout(n30_adj_1605),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_53_LC_11_11_7.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_53_LC_11_11_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_53_LC_11_11_7.LUT_INIT=16'b1111111110111011;
    LogicCell40 i1_2_lut_3_lut_adj_53_LC_11_11_7 (
            .in0(N__37571),
            .in1(N__56752),
            .in2(_gnd_net_),
            .in3(N__54006),
            .lcout(n28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_4_i26_3_lut_LC_11_12_0.C_ON=1'b0;
    defparam mux_129_Mux_4_i26_3_lut_LC_11_12_0.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_4_i26_3_lut_LC_11_12_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_129_Mux_4_i26_3_lut_LC_11_12_0 (
            .in0(N__30678),
            .in1(N__56874),
            .in2(_gnd_net_),
            .in3(N__37695),
            .lcout(),
            .ltout(n26_adj_1635_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19706_LC_11_12_1.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19706_LC_11_12_1.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19706_LC_11_12_1.LUT_INIT=16'b1011100011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_19706_LC_11_12_1 (
            .in0(N__57318),
            .in1(N__46296),
            .in2(N__30651),
            .in3(N__47706),
            .lcout(),
            .ltout(n22443_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22443_bdd_4_lut_LC_11_12_2.C_ON=1'b0;
    defparam n22443_bdd_4_lut_LC_11_12_2.SEQ_MODE=4'b0000;
    defparam n22443_bdd_4_lut_LC_11_12_2.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22443_bdd_4_lut_LC_11_12_2 (
            .in0(N__47707),
            .in1(N__32667),
            .in2(N__30648),
            .in3(N__35335),
            .lcout(),
            .ltout(n22446_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1569462_i1_3_lut_LC_11_12_3.C_ON=1'b0;
    defparam i1569462_i1_3_lut_LC_11_12_3.SEQ_MODE=4'b0000;
    defparam i1569462_i1_3_lut_LC_11_12_3.LUT_INIT=16'b1111000011001100;
    LogicCell40 i1569462_i1_3_lut_LC_11_12_3 (
            .in0(_gnd_net_),
            .in1(N__30564),
            .in2(N__30645),
            .in3(N__47269),
            .lcout(),
            .ltout(n30_adj_1636_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i4_LC_11_12_4.C_ON=1'b0;
    defparam comm_buf_1__i4_LC_11_12_4.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i4_LC_11_12_4.LUT_INIT=16'b1111101001010000;
    LogicCell40 comm_buf_1__i4_LC_11_12_4 (
            .in0(N__54571),
            .in1(_gnd_net_),
            .in2(N__30642),
            .in3(N__53644),
            .lcout(comm_buf_1_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55966),
            .ce(N__45213),
            .sr(N__44015));
    defparam comm_cmd_1__bdd_4_lut_19736_LC_11_12_5.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19736_LC_11_12_5.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19736_LC_11_12_5.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_19736_LC_11_12_5 (
            .in0(N__30639),
            .in1(N__46295),
            .in2(N__30633),
            .in3(N__47704),
            .lcout(),
            .ltout(n22467_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22467_bdd_4_lut_LC_11_12_6.C_ON=1'b0;
    defparam n22467_bdd_4_lut_LC_11_12_6.SEQ_MODE=4'b0000;
    defparam n22467_bdd_4_lut_LC_11_12_6.LUT_INIT=16'b1110010111100000;
    LogicCell40 n22467_bdd_4_lut_LC_11_12_6 (
            .in0(N__47705),
            .in1(N__30608),
            .in2(N__30579),
            .in3(N__30576),
            .lcout(n22470),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19726_LC_11_13_0.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19726_LC_11_13_0.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19726_LC_11_13_0.LUT_INIT=16'b1110011010100010;
    LogicCell40 comm_cmd_0__bdd_4_lut_19726_LC_11_13_0 (
            .in0(N__57203),
            .in1(N__46458),
            .in2(N__31045),
            .in3(N__30845),
            .lcout(),
            .ltout(n22395_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22395_bdd_4_lut_LC_11_13_1.C_ON=1'b0;
    defparam n22395_bdd_4_lut_LC_11_13_1.SEQ_MODE=4'b0000;
    defparam n22395_bdd_4_lut_LC_11_13_1.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22395_bdd_4_lut_LC_11_13_1 (
            .in0(N__46459),
            .in1(N__44791),
            .in2(N__30849),
            .in3(N__32727),
            .lcout(n22398),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_4_lut_adj_155_LC_11_13_2.C_ON=1'b0;
    defparam i3_4_lut_adj_155_LC_11_13_2.SEQ_MODE=4'b0000;
    defparam i3_4_lut_adj_155_LC_11_13_2.LUT_INIT=16'b0111101111011110;
    LogicCell40 i3_4_lut_adj_155_LC_11_13_2 (
            .in0(N__40905),
            .in1(N__37908),
            .in2(N__30846),
            .in3(N__34768),
            .lcout(n19_adj_1526),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_LC_11_13_3.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_LC_11_13_3.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_LC_11_13_3.LUT_INIT=16'b1111010110001000;
    LogicCell40 comm_cmd_0__bdd_4_lut_LC_11_13_3 (
            .in0(N__46456),
            .in1(N__30805),
            .in2(N__30780),
            .in3(N__57202),
            .lcout(),
            .ltout(n22635_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22635_bdd_4_lut_LC_11_13_4.C_ON=1'b0;
    defparam n22635_bdd_4_lut_LC_11_13_4.SEQ_MODE=4'b0000;
    defparam n22635_bdd_4_lut_LC_11_13_4.LUT_INIT=16'b1111000011001010;
    LogicCell40 n22635_bdd_4_lut_LC_11_13_4 (
            .in0(N__31323),
            .in1(N__35630),
            .in2(N__30738),
            .in3(N__46457),
            .lcout(n21236),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i13_LC_11_13_5.C_ON=1'b0;
    defparam req_data_cnt_i13_LC_11_13_5.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i13_LC_11_13_5.LUT_INIT=16'b1111000010101010;
    LogicCell40 req_data_cnt_i13_LC_11_13_5 (
            .in0(N__34769),
            .in1(_gnd_net_),
            .in2(N__30722),
            .in3(N__35570),
            .lcout(req_data_cnt_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55977),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i6_LC_11_13_6.C_ON=1'b0;
    defparam req_data_cnt_i6_LC_11_13_6.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i6_LC_11_13_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 req_data_cnt_i6_LC_11_13_6 (
            .in0(N__35571),
            .in1(N__31728),
            .in2(_gnd_net_),
            .in3(N__43517),
            .lcout(req_data_cnt_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55977),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i0_LC_11_13_7.C_ON=1'b0;
    defparam req_data_cnt_i0_LC_11_13_7.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i0_LC_11_13_7.LUT_INIT=16'b1011101110001000;
    LogicCell40 req_data_cnt_i0_LC_11_13_7 (
            .in0(N__43199),
            .in1(N__35569),
            .in2(_gnd_net_),
            .in3(N__43648),
            .lcout(req_data_cnt_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55977),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_state_2__I_0_371_Mux_0_i2_4_lut_4_lut_LC_11_14_0.C_ON=1'b0;
    defparam eis_state_2__I_0_371_Mux_0_i2_4_lut_4_lut_LC_11_14_0.SEQ_MODE=4'b0000;
    defparam eis_state_2__I_0_371_Mux_0_i2_4_lut_4_lut_LC_11_14_0.LUT_INIT=16'b0000011111110111;
    LogicCell40 eis_state_2__I_0_371_Mux_0_i2_4_lut_4_lut_LC_11_14_0 (
            .in0(N__31047),
            .in1(N__32816),
            .in2(N__30984),
            .in3(N__37780),
            .lcout(),
            .ltout(n2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_state_i0_LC_11_14_1.C_ON=1'b0;
    defparam eis_state_i0_LC_11_14_1.SEQ_MODE=4'b1010;
    defparam eis_state_i0_LC_11_14_1.LUT_INIT=16'b1111101000010001;
    LogicCell40 eis_state_i0_LC_11_14_1 (
            .in0(N__35792),
            .in1(N__30979),
            .in2(N__30681),
            .in3(N__31053),
            .lcout(eis_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVeis_state_i0C_net),
            .ce(N__30996),
            .sr(N__35732));
    defparam i19138_2_lut_4_lut_LC_11_14_2.C_ON=1'b0;
    defparam i19138_2_lut_4_lut_LC_11_14_2.SEQ_MODE=4'b0000;
    defparam i19138_2_lut_4_lut_LC_11_14_2.LUT_INIT=16'b1111101011111011;
    LogicCell40 i19138_2_lut_4_lut_LC_11_14_2 (
            .in0(N__43042),
            .in1(N__32421),
            .in2(N__30982),
            .in3(N__32069),
            .lcout(),
            .ltout(n21501_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_state_1__bdd_4_lut_LC_11_14_3.C_ON=1'b0;
    defparam eis_state_1__bdd_4_lut_LC_11_14_3.SEQ_MODE=4'b0000;
    defparam eis_state_1__bdd_4_lut_LC_11_14_3.LUT_INIT=16'b1110011011000100;
    LogicCell40 eis_state_1__bdd_4_lut_LC_11_14_3 (
            .in0(N__35791),
            .in1(N__35871),
            .in2(N__31062),
            .in3(N__31059),
            .lcout(n22479),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i29_4_lut_LC_11_14_4.C_ON=1'b0;
    defparam i29_4_lut_LC_11_14_4.SEQ_MODE=4'b0000;
    defparam i29_4_lut_LC_11_14_4.LUT_INIT=16'b1111110100001101;
    LogicCell40 i29_4_lut_LC_11_14_4 (
            .in0(N__31046),
            .in1(N__32817),
            .in2(N__30983),
            .in3(N__37779),
            .lcout(),
            .ltout(n11_adj_1632_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam eis_state_i2_LC_11_14_5.C_ON=1'b0;
    defparam eis_state_i2_LC_11_14_5.SEQ_MODE=4'b1010;
    defparam eis_state_i2_LC_11_14_5.LUT_INIT=16'b1110101001100010;
    LogicCell40 eis_state_i2_LC_11_14_5 (
            .in0(N__35793),
            .in1(N__35872),
            .in2(N__30999),
            .in3(N__30909),
            .lcout(eis_state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVeis_state_i0C_net),
            .ce(N__30996),
            .sr(N__35732));
    defparam i1_2_lut_4_lut_4_lut_LC_11_14_6.C_ON=1'b0;
    defparam i1_2_lut_4_lut_4_lut_LC_11_14_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_4_lut_4_lut_LC_11_14_6.LUT_INIT=16'b0100010001000101;
    LogicCell40 i1_2_lut_4_lut_4_lut_LC_11_14_6 (
            .in0(N__30969),
            .in1(N__43041),
            .in2(N__32073),
            .in3(N__32420),
            .lcout(n21041),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_1_i16_3_lut_LC_11_15_0.C_ON=1'b0;
    defparam mux_129_Mux_1_i16_3_lut_LC_11_15_0.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_1_i16_3_lut_LC_11_15_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_129_Mux_1_i16_3_lut_LC_11_15_0 (
            .in0(N__57207),
            .in1(N__35603),
            .in2(_gnd_net_),
            .in3(N__31198),
            .lcout(n16_adj_1651),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_2_i16_3_lut_LC_11_15_1.C_ON=1'b0;
    defparam mux_128_Mux_2_i16_3_lut_LC_11_15_1.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_2_i16_3_lut_LC_11_15_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_128_Mux_2_i16_3_lut_LC_11_15_1 (
            .in0(N__30862),
            .in1(N__31091),
            .in2(_gnd_net_),
            .in3(N__57206),
            .lcout(n16_adj_1681),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i15_LC_11_15_3.C_ON=1'b0;
    defparam buf_dds1_i15_LC_11_15_3.SEQ_MODE=4'b1000;
    defparam buf_dds1_i15_LC_11_15_3.LUT_INIT=16'b1000101010000000;
    LogicCell40 buf_dds1_i15_LC_11_15_3 (
            .in0(N__46755),
            .in1(N__42555),
            .in2(N__46899),
            .in3(N__30893),
            .lcout(buf_dds1_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56004),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i10_LC_11_15_4.C_ON=1'b0;
    defparam buf_dds1_i10_LC_11_15_4.SEQ_MODE=4'b1000;
    defparam buf_dds1_i10_LC_11_15_4.LUT_INIT=16'b1110001000000000;
    LogicCell40 buf_dds1_i10_LC_11_15_4 (
            .in0(N__30872),
            .in1(N__46874),
            .in2(N__45874),
            .in3(N__46756),
            .lcout(buf_dds1_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56004),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_4_lut_adj_161_LC_11_15_5.C_ON=1'b0;
    defparam i1_2_lut_4_lut_adj_161_LC_11_15_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_4_lut_adj_161_LC_11_15_5.LUT_INIT=16'b0000000000000100;
    LogicCell40 i1_2_lut_4_lut_adj_161_LC_11_15_5 (
            .in0(N__46453),
            .in1(N__47192),
            .in2(N__57261),
            .in3(N__47666),
            .lcout(n5_adj_1536),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i6_LC_11_15_6.C_ON=1'b0;
    defparam data_index_i6_LC_11_15_6.SEQ_MODE=4'b1000;
    defparam data_index_i6_LC_11_15_6.LUT_INIT=16'b0011101100001000;
    LogicCell40 data_index_i6_LC_11_15_6 (
            .in0(N__36129),
            .in1(N__55433),
            .in2(N__49341),
            .in3(N__38033),
            .lcout(data_index_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56004),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i1_LC_11_15_7.C_ON=1'b0;
    defparam buf_dds0_i1_LC_11_15_7.SEQ_MODE=4'b1000;
    defparam buf_dds0_i1_LC_11_15_7.LUT_INIT=16'b1100110010101010;
    LogicCell40 buf_dds0_i1_LC_11_15_7 (
            .in0(N__31199),
            .in1(N__36171),
            .in2(_gnd_net_),
            .in3(N__41662),
            .lcout(buf_dds0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56004),
            .ce(),
            .sr(_gnd_net_));
    defparam i8_4_lut_LC_11_16_0.C_ON=1'b0;
    defparam i8_4_lut_LC_11_16_0.SEQ_MODE=4'b0000;
    defparam i8_4_lut_LC_11_16_0.LUT_INIT=16'b0111110110111110;
    LogicCell40 i8_4_lut_LC_11_16_0 (
            .in0(N__36780),
            .in1(N__31171),
            .in2(N__37065),
            .in3(N__42973),
            .lcout(n24_adj_1593),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12382_2_lut_LC_11_16_2.C_ON=1'b0;
    defparam i12382_2_lut_LC_11_16_2.SEQ_MODE=4'b0000;
    defparam i12382_2_lut_LC_11_16_2.LUT_INIT=16'b0000000010101010;
    LogicCell40 i12382_2_lut_LC_11_16_2 (
            .in0(N__37808),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35870),
            .lcout(n14907),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_4_lut_LC_11_16_4.C_ON=1'b0;
    defparam i3_4_lut_LC_11_16_4.SEQ_MODE=4'b0000;
    defparam i3_4_lut_LC_11_16_4.LUT_INIT=16'b1111111111111011;
    LogicCell40 i3_4_lut_LC_11_16_4 (
            .in0(N__46460),
            .in1(N__47665),
            .in2(N__31158),
            .in3(N__54009),
            .lcout(n8841),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam EIS_SYNCCLK_I_0_1_lut_LC_11_16_6.C_ON=1'b0;
    defparam EIS_SYNCCLK_I_0_1_lut_LC_11_16_6.SEQ_MODE=4'b0000;
    defparam EIS_SYNCCLK_I_0_1_lut_LC_11_16_6.LUT_INIT=16'b0101010101010101;
    LogicCell40 EIS_SYNCCLK_I_0_1_lut_LC_11_16_6 (
            .in0(N__31140),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(IAC_CLK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i14_LC_11_16_7.C_ON=1'b0;
    defparam buf_dds0_i14_LC_11_16_7.SEQ_MODE=4'b1000;
    defparam buf_dds0_i14_LC_11_16_7.LUT_INIT=16'b0101000011001100;
    LogicCell40 buf_dds0_i14_LC_11_16_7 (
            .in0(N__49297),
            .in1(N__31318),
            .in2(N__49587),
            .in3(N__41658),
            .lcout(buf_dds0_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56021),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i10_LC_11_17_0 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i10_LC_11_17_0 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i10_LC_11_17_0 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \SIG_DDS.tmp_buf_i10_LC_11_17_0  (
            .in0(N__44638),
            .in1(N__44492),
            .in2(N__31233),
            .in3(N__31092),
            .lcout(\SIG_DDS.tmp_buf_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56035),
            .ce(N__43910),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i11_LC_11_17_1 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i11_LC_11_17_1 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i11_LC_11_17_1 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \SIG_DDS.tmp_buf_i11_LC_11_17_1  (
            .in0(N__44493),
            .in1(N__44642),
            .in2(N__31377),
            .in3(N__31368),
            .lcout(\SIG_DDS.tmp_buf_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56035),
            .ce(N__43910),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i12_LC_11_17_2 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i12_LC_11_17_2 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i12_LC_11_17_2 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \SIG_DDS.tmp_buf_i12_LC_11_17_2  (
            .in0(N__44639),
            .in1(N__44494),
            .in2(N__31350),
            .in3(N__36257),
            .lcout(\SIG_DDS.tmp_buf_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56035),
            .ce(N__43910),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i13_LC_11_17_3 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i13_LC_11_17_3 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i13_LC_11_17_3 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \SIG_DDS.tmp_buf_i13_LC_11_17_3  (
            .in0(N__44495),
            .in1(N__44643),
            .in2(N__31341),
            .in3(N__35310),
            .lcout(\SIG_DDS.tmp_buf_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56035),
            .ce(N__43910),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i14_LC_11_17_4 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i14_LC_11_17_4 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i14_LC_11_17_4 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \SIG_DDS.tmp_buf_i14_LC_11_17_4  (
            .in0(N__44640),
            .in1(N__44496),
            .in2(N__31332),
            .in3(N__31319),
            .lcout(\SIG_DDS.tmp_buf_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56035),
            .ce(N__43910),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i15_LC_11_17_5 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i15_LC_11_17_5 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i15_LC_11_17_5 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \SIG_DDS.tmp_buf_i15_LC_11_17_5  (
            .in0(N__44497),
            .in1(N__44644),
            .in2(N__31298),
            .in3(N__31263),
            .lcout(tmp_buf_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56035),
            .ce(N__43910),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i9_LC_11_17_6 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i9_LC_11_17_6 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i9_LC_11_17_6 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \SIG_DDS.tmp_buf_i9_LC_11_17_6  (
            .in0(N__44641),
            .in1(N__44499),
            .in2(N__31224),
            .in3(N__31257),
            .lcout(\SIG_DDS.tmp_buf_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56035),
            .ce(N__43910),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i8_LC_11_17_7 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i8_LC_11_17_7 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i8_LC_11_17_7 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \SIG_DDS.tmp_buf_i8_LC_11_17_7  (
            .in0(N__44498),
            .in1(N__36621),
            .in2(N__39081),
            .in3(N__44645),
            .lcout(\SIG_DDS.tmp_buf_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56035),
            .ce(N__43910),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i0_LC_11_18_0 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i0_LC_11_18_0 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i0_LC_11_18_0 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \SIG_DDS.tmp_buf_i0_LC_11_18_0  (
            .in0(N__44646),
            .in1(N__44449),
            .in2(N__39005),
            .in3(N__41538),
            .lcout(\SIG_DDS.tmp_buf_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56051),
            .ce(N__43911),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i1_LC_11_18_1 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i1_LC_11_18_1 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i1_LC_11_18_1 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \SIG_DDS.tmp_buf_i1_LC_11_18_1  (
            .in0(N__44450),
            .in1(N__44650),
            .in2(N__31212),
            .in3(N__31203),
            .lcout(\SIG_DDS.tmp_buf_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56051),
            .ce(N__43911),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i2_LC_11_18_2 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i2_LC_11_18_2 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i2_LC_11_18_2 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \SIG_DDS.tmp_buf_i2_LC_11_18_2  (
            .in0(N__44647),
            .in1(N__44451),
            .in2(N__31464),
            .in3(N__31455),
            .lcout(\SIG_DDS.tmp_buf_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56051),
            .ce(N__43911),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i3_LC_11_18_4 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i3_LC_11_18_4 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i3_LC_11_18_4 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \SIG_DDS.tmp_buf_i3_LC_11_18_4  (
            .in0(N__44648),
            .in1(N__32996),
            .in2(N__31434),
            .in3(N__44452),
            .lcout(\SIG_DDS.tmp_buf_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56051),
            .ce(N__43911),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i4_LC_11_18_5 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i4_LC_11_18_5 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i4_LC_11_18_5 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \SIG_DDS.tmp_buf_i4_LC_11_18_5  (
            .in0(N__44453),
            .in1(N__44651),
            .in2(N__31425),
            .in3(N__32256),
            .lcout(\SIG_DDS.tmp_buf_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56051),
            .ce(N__43911),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i5_LC_11_18_6 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i5_LC_11_18_6 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i5_LC_11_18_6 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \SIG_DDS.tmp_buf_i5_LC_11_18_6  (
            .in0(N__44649),
            .in1(N__44454),
            .in2(N__31416),
            .in3(N__33023),
            .lcout(\SIG_DDS.tmp_buf_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56051),
            .ce(N__43911),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i6_LC_11_18_7 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i6_LC_11_18_7 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i6_LC_11_18_7 .LUT_INIT=16'b0111001101000000;
    LogicCell40 \SIG_DDS.tmp_buf_i6_LC_11_18_7  (
            .in0(N__44455),
            .in1(N__44652),
            .in2(N__31407),
            .in3(N__41463),
            .lcout(\SIG_DDS.tmp_buf_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56051),
            .ce(N__43911),
            .sr(_gnd_net_));
    defparam \comm_spi.data_rx_i0_12301_12302_set_LC_12_3_1 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i0_12301_12302_set_LC_12_3_1 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_rx_i0_12301_12302_set_LC_12_3_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.data_rx_i0_12301_12302_set_LC_12_3_1  (
            .in0(N__36912),
            .in1(N__36887),
            .in2(_gnd_net_),
            .in3(N__45033),
            .lcout(\comm_spi.n14822 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__58358),
            .ce(),
            .sr(N__37170));
    defparam \ADC_VDC.adc_state_i0_LC_12_4_2 .C_ON=1'b0;
    defparam \ADC_VDC.adc_state_i0_LC_12_4_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.adc_state_i0_LC_12_4_2 .LUT_INIT=16'b0001000101010100;
    LogicCell40 \ADC_VDC.adc_state_i0_LC_12_4_2  (
            .in0(N__51859),
            .in1(N__51722),
            .in2(N__52000),
            .in3(N__51345),
            .lcout(\ADC_VDC.adc_state_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42372),
            .ce(N__31686),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i2_3_lut_adj_28_LC_12_4_3 .C_ON=1'b0;
    defparam \ADC_VDC.i2_3_lut_adj_28_LC_12_4_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i2_3_lut_adj_28_LC_12_4_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \ADC_VDC.i2_3_lut_adj_28_LC_12_4_3  (
            .in0(N__51993),
            .in1(N__51858),
            .in2(_gnd_net_),
            .in3(N__51184),
            .lcout(\ADC_VDC.n21007 ),
            .ltout(\ADC_VDC.n21007_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i19461_3_lut_LC_12_4_4 .C_ON=1'b0;
    defparam \ADC_VDC.i19461_3_lut_LC_12_4_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i19461_3_lut_LC_12_4_4 .LUT_INIT=16'b1010111100000000;
    LogicCell40 \ADC_VDC.i19461_3_lut_LC_12_4_4  (
            .in0(N__51331),
            .in1(_gnd_net_),
            .in2(N__31386),
            .in3(N__51721),
            .lcout(\ADC_VDC.n4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_2_lut_adj_27_LC_12_4_7 .C_ON=1'b0;
    defparam \ADC_VDC.i1_2_lut_adj_27_LC_12_4_7 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_2_lut_adj_27_LC_12_4_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ADC_VDC.i1_2_lut_adj_27_LC_12_4_7  (
            .in0(_gnd_net_),
            .in1(N__51720),
            .in2(_gnd_net_),
            .in3(N__51330),
            .lcout(\ADC_VDC.n21133 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_3_lut_3_lut_4_lut_LC_12_5_0 .C_ON=1'b0;
    defparam \ADC_VDC.i1_3_lut_3_lut_4_lut_LC_12_5_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_3_lut_3_lut_4_lut_LC_12_5_0 .LUT_INIT=16'b1100000011101010;
    LogicCell40 \ADC_VDC.i1_3_lut_3_lut_4_lut_LC_12_5_0  (
            .in0(N__31707),
            .in1(N__51385),
            .in2(N__51754),
            .in3(N__51857),
            .lcout(\ADC_VDC.n15273 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_4_lut_adj_33_LC_12_5_2 .C_ON=1'b0;
    defparam \ADC_VDC.i1_4_lut_adj_33_LC_12_5_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_4_lut_adj_33_LC_12_5_2 .LUT_INIT=16'b1010001010101010;
    LogicCell40 \ADC_VDC.i1_4_lut_adj_33_LC_12_5_2  (
            .in0(N__31701),
            .in1(N__51210),
            .in2(N__31695),
            .in3(N__31632),
            .lcout(\ADC_VDC.n42_adj_1452 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i2_3_lut_LC_12_6_0 .C_ON=1'b0;
    defparam \ADC_VDC.i2_3_lut_LC_12_6_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i2_3_lut_LC_12_6_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \ADC_VDC.i2_3_lut_LC_12_6_0  (
            .in0(N__34253),
            .in1(N__34273),
            .in2(_gnd_net_),
            .in3(N__34751),
            .lcout(\ADC_VDC.n20998 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_2_lut_4_lut_LC_12_6_1 .C_ON=1'b0;
    defparam \ADC_VDC.i1_2_lut_4_lut_LC_12_6_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_2_lut_4_lut_LC_12_6_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.i1_2_lut_4_lut_LC_12_6_1  (
            .in0(N__34750),
            .in1(N__34252),
            .in2(N__34275),
            .in3(N__34393),
            .lcout(\ADC_VDC.n11494 ),
            .ltout(\ADC_VDC.n11494_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i3_4_lut_LC_12_6_2 .C_ON=1'b0;
    defparam \ADC_VDC.i3_4_lut_LC_12_6_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i3_4_lut_LC_12_6_2 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \ADC_VDC.i3_4_lut_LC_12_6_2  (
            .in0(N__34297),
            .in1(N__31947),
            .in2(N__31665),
            .in3(N__34333),
            .lcout(\ADC_VDC.n15 ),
            .ltout(\ADC_VDC.n15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i18458_2_lut_LC_12_6_3 .C_ON=1'b0;
    defparam \ADC_VDC.i18458_2_lut_LC_12_6_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i18458_2_lut_LC_12_6_3 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \ADC_VDC.i18458_2_lut_LC_12_6_3  (
            .in0(N__51904),
            .in1(_gnd_net_),
            .in2(N__31635),
            .in3(_gnd_net_),
            .lcout(\ADC_VDC.n21185 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.ADC_DATA_i1_LC_12_6_4 .C_ON=1'b0;
    defparam \ADC_VDC.ADC_DATA_i1_LC_12_6_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.ADC_DATA_i1_LC_12_6_4 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \ADC_VDC.ADC_DATA_i1_LC_12_6_4  (
            .in0(N__31608),
            .in1(N__51456),
            .in2(N__31497),
            .in3(N__32195),
            .lcout(buf_adcdata_vdc_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42334),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i18476_2_lut_LC_12_6_5 .C_ON=1'b0;
    defparam \ADC_VDC.i18476_2_lut_LC_12_6_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i18476_2_lut_LC_12_6_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ADC_VDC.i18476_2_lut_LC_12_6_5  (
            .in0(_gnd_net_),
            .in1(N__34326),
            .in2(_gnd_net_),
            .in3(N__34296),
            .lcout(\ADC_VDC.n21203 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i18484_2_lut_LC_12_6_6 .C_ON=1'b0;
    defparam \ADC_VDC.i18484_2_lut_LC_12_6_6 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i18484_2_lut_LC_12_6_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \ADC_VDC.i18484_2_lut_LC_12_6_6  (
            .in0(_gnd_net_),
            .in1(N__34422),
            .in2(_gnd_net_),
            .in3(N__34359),
            .lcout(\ADC_VDC.n21211 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_4_lut_LC_12_6_7 .C_ON=1'b0;
    defparam \ADC_VDC.i1_4_lut_LC_12_6_7 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_4_lut_LC_12_6_7 .LUT_INIT=16'b1010001010101000;
    LogicCell40 \ADC_VDC.i1_4_lut_LC_12_6_7  (
            .in0(N__51455),
            .in1(N__51896),
            .in2(N__51762),
            .in3(N__51209),
            .lcout(\ADC_VDC.n13368 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i6_12325_12326_reset_LC_12_7_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i6_12325_12326_reset_LC_12_7_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i6_12325_12326_reset_LC_12_7_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i6_12325_12326_reset_LC_12_7_0  (
            .in0(N__34806),
            .in1(N__52632),
            .in2(_gnd_net_),
            .in3(N__57474),
            .lcout(\comm_spi.n14847 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__58400),
            .ce(),
            .sr(N__35226));
    defparam i15_4_lut_adj_203_LC_12_8_0.C_ON=1'b0;
    defparam i15_4_lut_adj_203_LC_12_8_0.SEQ_MODE=4'b0000;
    defparam i15_4_lut_adj_203_LC_12_8_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i15_4_lut_adj_203_LC_12_8_0 (
            .in0(N__31734),
            .in1(N__31791),
            .in2(N__34503),
            .in3(N__34578),
            .lcout(),
            .ltout(n20048_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7_4_lut_adj_204_LC_12_8_1.C_ON=1'b0;
    defparam i7_4_lut_adj_204_LC_12_8_1.SEQ_MODE=4'b0000;
    defparam i7_4_lut_adj_204_LC_12_8_1.LUT_INIT=16'b0000100000000000;
    LogicCell40 i7_4_lut_adj_204_LC_12_8_1 (
            .in0(N__31932),
            .in1(N__35115),
            .in2(N__31914),
            .in3(N__31911),
            .lcout(n14899),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_4_i19_3_lut_LC_12_8_2.C_ON=1'b0;
    defparam mux_128_Mux_4_i19_3_lut_LC_12_8_2.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_4_i19_3_lut_LC_12_8_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_128_Mux_4_i19_3_lut_LC_12_8_2 (
            .in0(N__31902),
            .in1(N__31871),
            .in2(_gnd_net_),
            .in3(N__57184),
            .lcout(n19_adj_1673),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i11_4_lut_adj_200_LC_12_8_3.C_ON=1'b0;
    defparam i11_4_lut_adj_200_LC_12_8_3.SEQ_MODE=4'b0000;
    defparam i11_4_lut_adj_200_LC_12_8_3.LUT_INIT=16'b1111111111111110;
    LogicCell40 i11_4_lut_adj_200_LC_12_8_3 (
            .in0(N__31844),
            .in1(N__31832),
            .in2(N__31821),
            .in3(N__31802),
            .lcout(n27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10_4_lut_adj_199_LC_12_8_4.C_ON=1'b0;
    defparam i10_4_lut_adj_199_LC_12_8_4.SEQ_MODE=4'b0000;
    defparam i10_4_lut_adj_199_LC_12_8_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i10_4_lut_adj_199_LC_12_8_4 (
            .in0(N__31784),
            .in1(N__31772),
            .in2(N__31761),
            .in3(N__31745),
            .lcout(n26_adj_1656),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15472_2_lut_3_lut_LC_12_8_6.C_ON=1'b0;
    defparam i15472_2_lut_3_lut_LC_12_8_6.SEQ_MODE=4'b0000;
    defparam i15472_2_lut_3_lut_LC_12_8_6.LUT_INIT=16'b0000000000100010;
    LogicCell40 i15472_2_lut_3_lut_LC_12_8_6 (
            .in0(N__49496),
            .in1(N__54851),
            .in2(_gnd_net_),
            .in3(N__54341),
            .lcout(n14_adj_1552),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i14_4_lut_adj_158_LC_12_9_0.C_ON=1'b0;
    defparam i14_4_lut_adj_158_LC_12_9_0.SEQ_MODE=4'b0000;
    defparam i14_4_lut_adj_158_LC_12_9_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i14_4_lut_adj_158_LC_12_9_0 (
            .in0(N__31953),
            .in1(N__34866),
            .in2(N__34728),
            .in3(N__34461),
            .lcout(n30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i10_LC_12_9_1.C_ON=1'b0;
    defparam req_data_cnt_i10_LC_12_9_1.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i10_LC_12_9_1.LUT_INIT=16'b1011101110001000;
    LogicCell40 req_data_cnt_i10_LC_12_9_1 (
            .in0(N__32046),
            .in1(N__35533),
            .in2(_gnd_net_),
            .in3(N__35206),
            .lcout(req_data_cnt_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55942),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i11_LC_12_9_2.C_ON=1'b0;
    defparam req_data_cnt_i11_LC_12_9_2.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i11_LC_12_9_2.LUT_INIT=16'b1111101000001010;
    LogicCell40 req_data_cnt_i11_LC_12_9_2 (
            .in0(N__31967),
            .in1(_gnd_net_),
            .in2(N__35556),
            .in3(N__35246),
            .lcout(req_data_cnt_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55942),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i15_LC_12_9_3.C_ON=1'b0;
    defparam req_data_cnt_i15_LC_12_9_3.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i15_LC_12_9_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 req_data_cnt_i15_LC_12_9_3 (
            .in0(N__37476),
            .in1(N__35537),
            .in2(_gnd_net_),
            .in3(N__34480),
            .lcout(req_data_cnt_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55942),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i7_LC_12_9_4.C_ON=1'b0;
    defparam req_data_cnt_i7_LC_12_9_4.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i7_LC_12_9_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 req_data_cnt_i7_LC_12_9_4 (
            .in0(N__35538),
            .in1(N__32270),
            .in2(_gnd_net_),
            .in3(N__46571),
            .lcout(req_data_cnt_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55942),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_3_i30_3_lut_LC_12_9_5.C_ON=1'b0;
    defparam mux_130_Mux_3_i30_3_lut_LC_12_9_5.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_3_i30_3_lut_LC_12_9_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_130_Mux_3_i30_3_lut_LC_12_9_5 (
            .in0(N__32019),
            .in1(N__32001),
            .in2(_gnd_net_),
            .in3(N__47258),
            .lcout(n30_adj_1611),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7_4_lut_adj_149_LC_12_9_7.C_ON=1'b0;
    defparam i7_4_lut_adj_149_LC_12_9_7.SEQ_MODE=4'b0000;
    defparam i7_4_lut_adj_149_LC_12_9_7.LUT_INIT=16'b0111101111011110;
    LogicCell40 i7_4_lut_adj_149_LC_12_9_7 (
            .in0(N__37887),
            .in1(N__37962),
            .in2(N__31992),
            .in3(N__31966),
            .lcout(n23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i5_LC_12_10_0.C_ON=1'b0;
    defparam buf_cfgRTD_i5_LC_12_10_0.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i5_LC_12_10_0.LUT_INIT=16'b0111010100100000;
    LogicCell40 buf_cfgRTD_i5_LC_12_10_0 (
            .in0(N__39649),
            .in1(N__49388),
            .in2(N__52275),
            .in3(N__34919),
            .lcout(buf_cfgRTD_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55944),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i5_LC_12_10_1.C_ON=1'b0;
    defparam req_data_cnt_i5_LC_12_10_1.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i5_LC_12_10_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 req_data_cnt_i5_LC_12_10_1 (
            .in0(N__35558),
            .in1(N__37250),
            .in2(_gnd_net_),
            .in3(N__32305),
            .lcout(req_data_cnt_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55944),
            .ce(),
            .sr(_gnd_net_));
    defparam i15471_2_lut_3_lut_LC_12_10_3.C_ON=1'b0;
    defparam i15471_2_lut_3_lut_LC_12_10_3.SEQ_MODE=4'b0000;
    defparam i15471_2_lut_3_lut_LC_12_10_3.LUT_INIT=16'b0000000000100010;
    LogicCell40 i15471_2_lut_3_lut_LC_12_10_3 (
            .in0(N__44061),
            .in1(N__54825),
            .in2(_gnd_net_),
            .in3(N__54501),
            .lcout(n14_adj_1551),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i3_LC_12_10_4.C_ON=1'b0;
    defparam req_data_cnt_i3_LC_12_10_4.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i3_LC_12_10_4.LUT_INIT=16'b1011101110001000;
    LogicCell40 req_data_cnt_i3_LC_12_10_4 (
            .in0(N__36481),
            .in1(N__35557),
            .in2(_gnd_net_),
            .in3(N__41192),
            .lcout(req_data_cnt_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55944),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i4_LC_12_10_5.C_ON=1'b0;
    defparam buf_dds0_i4_LC_12_10_5.SEQ_MODE=4'b1000;
    defparam buf_dds0_i4_LC_12_10_5.LUT_INIT=16'b0101000011001100;
    LogicCell40 buf_dds0_i4_LC_12_10_5 (
            .in0(N__49387),
            .in1(N__32245),
            .in2(N__42707),
            .in3(N__41669),
            .lcout(buf_dds0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55944),
            .ce(),
            .sr(_gnd_net_));
    defparam i14639_3_lut_LC_12_10_6.C_ON=1'b0;
    defparam i14639_3_lut_LC_12_10_6.SEQ_MODE=4'b0000;
    defparam i14639_3_lut_LC_12_10_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 i14639_3_lut_LC_12_10_6 (
            .in0(N__32216),
            .in1(N__50720),
            .in2(_gnd_net_),
            .in3(N__57093),
            .lcout(n23_adj_1661),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i7_4_lut_LC_12_10_7.C_ON=1'b0;
    defparam i7_4_lut_LC_12_10_7.SEQ_MODE=4'b0000;
    defparam i7_4_lut_LC_12_10_7.LUT_INIT=16'b0110111111110110;
    LogicCell40 i7_4_lut_LC_12_10_7 (
            .in0(N__37092),
            .in1(N__32215),
            .in2(N__36756),
            .in3(N__32554),
            .lcout(n23_adj_1591),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i4_LC_12_11_0.C_ON=1'b0;
    defparam req_data_cnt_i4_LC_12_11_0.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i4_LC_12_11_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 req_data_cnt_i4_LC_12_11_0 (
            .in0(N__35559),
            .in1(N__36197),
            .in2(_gnd_net_),
            .in3(N__35336),
            .lcout(req_data_cnt_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55950),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_1_i19_3_lut_LC_12_11_1.C_ON=1'b0;
    defparam mux_130_Mux_1_i19_3_lut_LC_12_11_1.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_1_i19_3_lut_LC_12_11_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_130_Mux_1_i19_3_lut_LC_12_11_1 (
            .in0(N__32202),
            .in1(N__32174),
            .in2(_gnd_net_),
            .in3(N__57023),
            .lcout(n19_adj_1616),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_4_i17_3_lut_LC_12_11_2.C_ON=1'b0;
    defparam mux_128_Mux_4_i17_3_lut_LC_12_11_2.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_4_i17_3_lut_LC_12_11_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_128_Mux_4_i17_3_lut_LC_12_11_2 (
            .in0(N__57024),
            .in1(N__32141),
            .in2(_gnd_net_),
            .in3(N__32089),
            .lcout(n17_adj_1672),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i4_LC_12_11_3.C_ON=1'b0;
    defparam comm_cmd_i4_LC_12_11_3.SEQ_MODE=4'b1000;
    defparam comm_cmd_i4_LC_12_11_3.LUT_INIT=16'b1011100000110000;
    LogicCell40 comm_cmd_i4_LC_12_11_3 (
            .in0(N__50983),
            .in1(N__37523),
            .in2(N__32391),
            .in3(N__53640),
            .lcout(comm_cmd_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55950),
            .ce(),
            .sr(_gnd_net_));
    defparam i4_4_lut_adj_153_LC_12_11_4.C_ON=1'b0;
    defparam i4_4_lut_adj_153_LC_12_11_4.SEQ_MODE=4'b0000;
    defparam i4_4_lut_adj_153_LC_12_11_4.LUT_INIT=16'b0111101111011110;
    LogicCell40 i4_4_lut_adj_153_LC_12_11_4 (
            .in0(N__37668),
            .in1(N__41223),
            .in2(N__32306),
            .in3(N__41188),
            .lcout(n20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i5_LC_12_11_5.C_ON=1'b0;
    defparam comm_cmd_i5_LC_12_11_5.SEQ_MODE=4'b1000;
    defparam comm_cmd_i5_LC_12_11_5.LUT_INIT=16'b1100000010101010;
    LogicCell40 comm_cmd_i5_LC_12_11_5 (
            .in0(N__48821),
            .in1(N__53342),
            .in2(N__50990),
            .in3(N__37524),
            .lcout(comm_cmd_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55950),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_LC_12_11_6.C_ON=1'b0;
    defparam i2_3_lut_LC_12_11_6.SEQ_MODE=4'b0000;
    defparam i2_3_lut_LC_12_11_6.LUT_INIT=16'b1111111111011101;
    LogicCell40 i2_3_lut_LC_12_11_6 (
            .in0(N__32377),
            .in1(N__48847),
            .in2(_gnd_net_),
            .in3(N__48820),
            .lcout(n16818),
            .ltout(n16818_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_LC_12_11_7.C_ON=1'b0;
    defparam i1_2_lut_LC_12_11_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_LC_12_11_7.LUT_INIT=16'b1111000011111111;
    LogicCell40 i1_2_lut_LC_12_11_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32364),
            .in3(N__47132),
            .lcout(n12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22365_bdd_4_lut_LC_12_12_1.C_ON=1'b0;
    defparam n22365_bdd_4_lut_LC_12_12_1.SEQ_MODE=4'b0000;
    defparam n22365_bdd_4_lut_LC_12_12_1.LUT_INIT=16'b1100110011100010;
    LogicCell40 n22365_bdd_4_lut_LC_12_12_1 (
            .in0(N__32361),
            .in1(N__32346),
            .in2(N__33084),
            .in3(N__47671),
            .lcout(n22368),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_5_i26_3_lut_LC_12_12_2.C_ON=1'b0;
    defparam mux_129_Mux_5_i26_3_lut_LC_12_12_2.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_5_i26_3_lut_LC_12_12_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_129_Mux_5_i26_3_lut_LC_12_12_2 (
            .in0(N__32334),
            .in1(N__57194),
            .in2(_gnd_net_),
            .in3(N__37667),
            .lcout(),
            .ltout(n26_adj_1630_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19711_LC_12_12_3.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19711_LC_12_12_3.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19711_LC_12_12_3.LUT_INIT=16'b1011100011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_19711_LC_12_12_3 (
            .in0(N__57336),
            .in1(N__46297),
            .in2(N__32313),
            .in3(N__47672),
            .lcout(),
            .ltout(n22449_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22449_bdd_4_lut_LC_12_12_4.C_ON=1'b0;
    defparam n22449_bdd_4_lut_LC_12_12_4.SEQ_MODE=4'b0000;
    defparam n22449_bdd_4_lut_LC_12_12_4.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22449_bdd_4_lut_LC_12_12_4 (
            .in0(N__47673),
            .in1(N__32976),
            .in2(N__32310),
            .in3(N__32307),
            .lcout(),
            .ltout(n22452_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1570065_i1_3_lut_LC_12_12_5.C_ON=1'b0;
    defparam i1570065_i1_3_lut_LC_12_12_5.SEQ_MODE=4'b0000;
    defparam i1570065_i1_3_lut_LC_12_12_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 i1570065_i1_3_lut_LC_12_12_5 (
            .in0(_gnd_net_),
            .in1(N__32283),
            .in2(N__32277),
            .in3(N__47243),
            .lcout(),
            .ltout(n30_adj_1631_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i5_LC_12_12_6.C_ON=1'b0;
    defparam comm_buf_1__i5_LC_12_12_6.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i5_LC_12_12_6.LUT_INIT=16'b1010101011110000;
    LogicCell40 comm_buf_1__i5_LC_12_12_6 (
            .in0(N__53343),
            .in1(_gnd_net_),
            .in2(N__32640),
            .in3(N__54572),
            .lcout(comm_buf_1_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55954),
            .ce(N__45212),
            .sr(N__44016));
    defparam equal_188_i9_2_lut_3_lut_LC_12_13_0.C_ON=1'b0;
    defparam equal_188_i9_2_lut_3_lut_LC_12_13_0.SEQ_MODE=4'b0000;
    defparam equal_188_i9_2_lut_3_lut_LC_12_13_0.LUT_INIT=16'b1111111111011101;
    LogicCell40 equal_188_i9_2_lut_3_lut_LC_12_13_0 (
            .in0(N__46410),
            .in1(N__47667),
            .in2(_gnd_net_),
            .in3(N__57132),
            .lcout(n9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18603_4_lut_LC_12_13_1.C_ON=1'b0;
    defparam i18603_4_lut_LC_12_13_1.SEQ_MODE=4'b0000;
    defparam i18603_4_lut_LC_12_13_1.LUT_INIT=16'b0100010010100000;
    LogicCell40 i18603_4_lut_LC_12_13_1 (
            .in0(N__57133),
            .in1(N__32625),
            .in2(N__32604),
            .in3(N__46411),
            .lcout(n21330),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_3_i23_3_lut_LC_12_13_2.C_ON=1'b0;
    defparam mux_128_Mux_3_i23_3_lut_LC_12_13_2.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_3_i23_3_lut_LC_12_13_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_128_Mux_3_i23_3_lut_LC_12_13_2 (
            .in0(N__32561),
            .in1(N__36214),
            .in2(_gnd_net_),
            .in3(N__57134),
            .lcout(n23_adj_1677),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i9_LC_12_13_3.C_ON=1'b0;
    defparam buf_dds1_i9_LC_12_13_3.SEQ_MODE=4'b1000;
    defparam buf_dds1_i9_LC_12_13_3.LUT_INIT=16'b1100000010100000;
    LogicCell40 buf_dds1_i9_LC_12_13_3 (
            .in0(N__32518),
            .in1(N__53435),
            .in2(N__46767),
            .in3(N__46873),
            .lcout(buf_dds1_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55963),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_6_i19_3_lut_LC_12_13_4.C_ON=1'b0;
    defparam mux_129_Mux_6_i19_3_lut_LC_12_13_4.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_6_i19_3_lut_LC_12_13_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_129_Mux_6_i19_3_lut_LC_12_13_4 (
            .in0(N__32499),
            .in1(N__32468),
            .in2(_gnd_net_),
            .in3(N__57135),
            .lcout(n19_adj_1625),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_157_LC_12_13_5.C_ON=1'b0;
    defparam i1_4_lut_adj_157_LC_12_13_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_157_LC_12_13_5.LUT_INIT=16'b0111101111011110;
    LogicCell40 i1_4_lut_adj_157_LC_12_13_5 (
            .in0(N__43844),
            .in1(N__43437),
            .in2(N__43649),
            .in3(N__43513),
            .lcout(),
            .ltout(n17_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i13_4_lut_adj_160_LC_12_13_6.C_ON=1'b0;
    defparam i13_4_lut_adj_160_LC_12_13_6.SEQ_MODE=4'b0000;
    defparam i13_4_lut_adj_160_LC_12_13_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i13_4_lut_adj_160_LC_12_13_6 (
            .in0(N__35316),
            .in1(N__32439),
            .in2(N__32430),
            .in3(N__32427),
            .lcout(n29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19285_2_lut_LC_12_13_7.C_ON=1'b0;
    defparam i19285_2_lut_LC_12_13_7.SEQ_MODE=4'b0000;
    defparam i19285_2_lut_LC_12_13_7.LUT_INIT=16'b1010101000000000;
    LogicCell40 i19285_2_lut_LC_12_13_7 (
            .in0(N__57136),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32412),
            .lcout(n21671),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_3_i16_3_lut_LC_12_14_0.C_ON=1'b0;
    defparam mux_129_Mux_3_i16_3_lut_LC_12_14_0.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_3_i16_3_lut_LC_12_14_0.LUT_INIT=16'b1100110010101010;
    LogicCell40 mux_129_Mux_3_i16_3_lut_LC_12_14_0 (
            .in0(N__32997),
            .in1(N__32683),
            .in2(_gnd_net_),
            .in3(N__57147),
            .lcout(n16_adj_1640),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i0_LC_12_14_1.C_ON=1'b0;
    defparam buf_control_i0_LC_12_14_1.SEQ_MODE=4'b1000;
    defparam buf_control_i0_LC_12_14_1.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_control_i0_LC_12_14_1 (
            .in0(N__49280),
            .in1(N__42001),
            .in2(N__45645),
            .in3(N__44792),
            .lcout(buf_control_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55974),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i3_LC_12_14_2.C_ON=1'b0;
    defparam buf_dds1_i3_LC_12_14_2.SEQ_MODE=4'b1000;
    defparam buf_dds1_i3_LC_12_14_2.LUT_INIT=16'b1110111000101110;
    LogicCell40 buf_dds1_i3_LC_12_14_2 (
            .in0(N__32687),
            .in1(N__46872),
            .in2(N__55434),
            .in3(N__36485),
            .lcout(buf_dds1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55974),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i0_LC_12_14_3.C_ON=1'b0;
    defparam acadc_skipCount_i0_LC_12_14_3.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i0_LC_12_14_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 acadc_skipCount_i0_LC_12_14_3 (
            .in0(N__43198),
            .in1(N__47905),
            .in2(_gnd_net_),
            .in3(N__43676),
            .lcout(acadc_skipCount_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55974),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i4_LC_12_14_4.C_ON=1'b0;
    defparam acadc_skipCount_i4_LC_12_14_4.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i4_LC_12_14_4.LUT_INIT=16'b1111010110100000;
    LogicCell40 acadc_skipCount_i4_LC_12_14_4 (
            .in0(N__47907),
            .in1(_gnd_net_),
            .in2(N__36196),
            .in3(N__32660),
            .lcout(acadc_skipCount_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55974),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i1_LC_12_14_5.C_ON=1'b0;
    defparam acadc_skipCount_i1_LC_12_14_5.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i1_LC_12_14_5.LUT_INIT=16'b1100110010101010;
    LogicCell40 acadc_skipCount_i1_LC_12_14_5 (
            .in0(N__44165),
            .in1(N__36165),
            .in2(_gnd_net_),
            .in3(N__47906),
            .lcout(acadc_skipCount_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55974),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_LC_12_14_6.C_ON=1'b0;
    defparam i2_4_lut_LC_12_14_6.SEQ_MODE=4'b0000;
    defparam i2_4_lut_LC_12_14_6.LUT_INIT=16'b0111110110111110;
    LogicCell40 i2_4_lut_LC_12_14_6 (
            .in0(N__36726),
            .in1(N__32659),
            .in2(N__36660),
            .in3(N__44164),
            .lcout(n18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i6_LC_12_14_7.C_ON=1'b0;
    defparam acadc_skipCount_i6_LC_12_14_7.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i6_LC_12_14_7.LUT_INIT=16'b0111001101000000;
    LogicCell40 acadc_skipCount_i6_LC_12_14_7 (
            .in0(N__49279),
            .in1(N__47908),
            .in2(N__49497),
            .in3(N__43538),
            .lcout(acadc_skipCount_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55974),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i7_LC_12_15_0.C_ON=1'b0;
    defparam data_index_i7_LC_12_15_0.SEQ_MODE=4'b1000;
    defparam data_index_i7_LC_12_15_0.LUT_INIT=16'b0011101100001000;
    LogicCell40 data_index_i7_LC_12_15_0 (
            .in0(N__32646),
            .in1(N__55432),
            .in2(N__49316),
            .in3(N__37989),
            .lcout(data_index_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55986),
            .ce(),
            .sr(_gnd_net_));
    defparam i6314_3_lut_LC_12_15_1.C_ON=1'b0;
    defparam i6314_3_lut_LC_12_15_1.SEQ_MODE=4'b0000;
    defparam i6314_3_lut_LC_12_15_1.LUT_INIT=16'b1100110010101010;
    LogicCell40 i6314_3_lut_LC_12_15_1 (
            .in0(N__44059),
            .in1(N__38008),
            .in2(_gnd_net_),
            .in3(N__41096),
            .lcout(n8_adj_1560),
            .ltout(n8_adj_1560_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_354_Mux_7_i15_4_lut_LC_12_15_2.C_ON=1'b0;
    defparam comm_state_3__I_0_354_Mux_7_i15_4_lut_LC_12_15_2.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_354_Mux_7_i15_4_lut_LC_12_15_2.LUT_INIT=16'b0111001101000000;
    LogicCell40 comm_state_3__I_0_354_Mux_7_i15_4_lut_LC_12_15_2 (
            .in0(N__49203),
            .in1(N__55431),
            .in2(N__32949),
            .in3(N__37988),
            .lcout(data_index_9_N_212_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i7_LC_12_15_3.C_ON=1'b0;
    defparam acadc_skipCount_i7_LC_12_15_3.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i7_LC_12_15_3.LUT_INIT=16'b0000110010101100;
    LogicCell40 acadc_skipCount_i7_LC_12_15_3 (
            .in0(N__44060),
            .in1(N__46598),
            .in2(N__47922),
            .in3(N__49207),
            .lcout(acadc_skipCount_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55986),
            .ce(),
            .sr(_gnd_net_));
    defparam i6_4_lut_adj_63_LC_12_15_4.C_ON=1'b0;
    defparam i6_4_lut_adj_63_LC_12_15_4.SEQ_MODE=4'b0000;
    defparam i6_4_lut_adj_63_LC_12_15_4.LUT_INIT=16'b0111110110111110;
    LogicCell40 i6_4_lut_adj_63_LC_12_15_4 (
            .in0(N__36702),
            .in1(N__46594),
            .in2(N__36825),
            .in3(N__35392),
            .lcout(),
            .ltout(n22_adj_1590_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i14_4_lut_adj_75_LC_12_15_5.C_ON=1'b0;
    defparam i14_4_lut_adj_75_LC_12_15_5.SEQ_MODE=4'b0000;
    defparam i14_4_lut_adj_75_LC_12_15_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i14_4_lut_adj_75_LC_12_15_5 (
            .in0(N__32844),
            .in1(N__32838),
            .in2(N__32829),
            .in3(N__50592),
            .lcout(),
            .ltout(n30_adj_1543_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15_4_lut_adj_79_LC_12_15_6.C_ON=1'b0;
    defparam i15_4_lut_adj_79_LC_12_15_6.SEQ_MODE=4'b0000;
    defparam i15_4_lut_adj_79_LC_12_15_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i15_4_lut_adj_79_LC_12_15_6 (
            .in0(N__32826),
            .in1(N__36021),
            .in2(N__32820),
            .in3(N__32694),
            .lcout(n31_adj_1537),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i2_LC_12_15_7.C_ON=1'b0;
    defparam acadc_skipCount_i2_LC_12_15_7.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i2_LC_12_15_7.LUT_INIT=16'b1111101000001010;
    LogicCell40 acadc_skipCount_i2_LC_12_15_7 (
            .in0(N__35393),
            .in1(_gnd_net_),
            .in2(N__47921),
            .in3(N__34860),
            .lcout(acadc_skipCount_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55986),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i18_LC_12_16_0 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i18_LC_12_16_0 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i18_LC_12_16_0 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i18_LC_12_16_0  (
            .in0(N__38599),
            .in1(N__38748),
            .in2(N__32796),
            .in3(N__32749),
            .lcout(buf_adcdata_iac_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55999),
            .ce(),
            .sr(_gnd_net_));
    defparam equal_61_i14_2_lut_LC_12_16_1.C_ON=1'b0;
    defparam equal_61_i14_2_lut_LC_12_16_1.SEQ_MODE=4'b0000;
    defparam equal_61_i14_2_lut_LC_12_16_1.LUT_INIT=16'b0011001111001100;
    LogicCell40 equal_61_i14_2_lut_LC_12_16_1 (
            .in0(_gnd_net_),
            .in1(N__37113),
            .in2(_gnd_net_),
            .in3(N__33040),
            .lcout(),
            .ltout(n14_adj_1538_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i10_4_lut_LC_12_16_2.C_ON=1'b0;
    defparam i10_4_lut_LC_12_16_2.SEQ_MODE=4'b0000;
    defparam i10_4_lut_LC_12_16_2.LUT_INIT=16'b1111111111110110;
    LogicCell40 i10_4_lut_LC_12_16_2 (
            .in0(N__36801),
            .in1(N__32726),
            .in2(N__32697),
            .in3(N__32955),
            .lcout(n26_adj_1525),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i13_LC_12_16_3 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i13_LC_12_16_3 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i13_LC_12_16_3 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_IAC.ADC_DATA_i13_LC_12_16_3  (
            .in0(N__38747),
            .in1(N__38600),
            .in2(N__33083),
            .in3(N__33113),
            .lcout(buf_adcdata_iac_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55999),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i13_LC_12_16_4.C_ON=1'b0;
    defparam acadc_skipCount_i13_LC_12_16_4.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i13_LC_12_16_4.LUT_INIT=16'b0011000010101010;
    LogicCell40 acadc_skipCount_i13_LC_12_16_4 (
            .in0(N__33041),
            .in1(N__49318),
            .in2(N__52286),
            .in3(N__47909),
            .lcout(acadc_skipCount_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55999),
            .ce(),
            .sr(_gnd_net_));
    defparam i6324_3_lut_LC_12_16_5.C_ON=1'b0;
    defparam i6324_3_lut_LC_12_16_5.SEQ_MODE=4'b0000;
    defparam i6324_3_lut_LC_12_16_5.LUT_INIT=16'b1110111001000100;
    LogicCell40 i6324_3_lut_LC_12_16_5 (
            .in0(N__41079),
            .in1(N__49494),
            .in2(_gnd_net_),
            .in3(N__38050),
            .lcout(n8_adj_1562),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i5_LC_12_16_6.C_ON=1'b0;
    defparam buf_dds0_i5_LC_12_16_6.SEQ_MODE=4'b1000;
    defparam buf_dds0_i5_LC_12_16_6.LUT_INIT=16'b0101000011001100;
    LogicCell40 buf_dds0_i5_LC_12_16_6 (
            .in0(N__49134),
            .in1(N__33016),
            .in2(N__50424),
            .in3(N__41613),
            .lcout(buf_dds0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55999),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i5_LC_12_16_7.C_ON=1'b0;
    defparam acadc_skipCount_i5_LC_12_16_7.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i5_LC_12_16_7.LUT_INIT=16'b0101110100001000;
    LogicCell40 acadc_skipCount_i5_LC_12_16_7 (
            .in0(N__47910),
            .in1(N__50418),
            .in2(N__49376),
            .in3(N__32975),
            .lcout(acadc_skipCount_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55999),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.dds_state_i2_LC_12_17_0 .C_ON=1'b0;
    defparam \SIG_DDS.dds_state_i2_LC_12_17_0 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.dds_state_i2_LC_12_17_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \SIG_DDS.dds_state_i2_LC_12_17_0  (
            .in0(N__44515),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44653),
            .lcout(dds_state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56015),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i3_LC_12_17_1.C_ON=1'b0;
    defparam buf_dds0_i3_LC_12_17_1.SEQ_MODE=4'b1000;
    defparam buf_dds0_i3_LC_12_17_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 buf_dds0_i3_LC_12_17_1 (
            .in0(N__36465),
            .in1(N__32995),
            .in2(_gnd_net_),
            .in3(N__41657),
            .lcout(buf_dds0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56015),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i3_LC_12_17_2.C_ON=1'b0;
    defparam acadc_skipCount_i3_LC_12_17_2.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i3_LC_12_17_2.LUT_INIT=16'b1100110010101010;
    LogicCell40 acadc_skipCount_i3_LC_12_17_2 (
            .in0(N__41162),
            .in1(N__36466),
            .in2(_gnd_net_),
            .in3(N__47916),
            .lcout(acadc_skipCount_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56015),
            .ce(),
            .sr(_gnd_net_));
    defparam i4_4_lut_LC_12_17_3.C_ON=1'b0;
    defparam i4_4_lut_LC_12_17_3.SEQ_MODE=4'b0000;
    defparam i4_4_lut_LC_12_17_3.LUT_INIT=16'b0111110110111110;
    LogicCell40 i4_4_lut_LC_12_17_3 (
            .in0(N__36681),
            .in1(N__32971),
            .in2(N__36867),
            .in3(N__41161),
            .lcout(n20_adj_1670),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i8_LC_12_17_4 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i8_LC_12_17_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i8_LC_12_17_4 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_IAC.ADC_DATA_i8_LC_12_17_4  (
            .in0(N__38505),
            .in1(N__38771),
            .in2(N__41701),
            .in3(N__33810),
            .lcout(buf_adcdata_iac_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56015),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i9_LC_12_17_6 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i9_LC_12_17_6 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i9_LC_12_17_6 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \ADC_IAC.ADC_DATA_i9_LC_12_17_6  (
            .in0(N__38506),
            .in1(N__38772),
            .in2(N__33783),
            .in3(N__43601),
            .lcout(buf_adcdata_iac_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56015),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i8_LC_12_17_7.C_ON=1'b0;
    defparam buf_dds0_i8_LC_12_17_7.SEQ_MODE=4'b1000;
    defparam buf_dds0_i8_LC_12_17_7.LUT_INIT=16'b0011101000001010;
    LogicCell40 buf_dds0_i8_LC_12_17_7 (
            .in0(N__39076),
            .in1(N__49322),
            .in2(N__41670),
            .in3(N__45634),
            .lcout(buf_dds0_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56015),
            .ce(),
            .sr(_gnd_net_));
    defparam data_count_i0_i0_LC_12_18_0.C_ON=1'b1;
    defparam data_count_i0_i0_LC_12_18_0.SEQ_MODE=4'b1000;
    defparam data_count_i0_i0_LC_12_18_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i0_LC_12_18_0 (
            .in0(_gnd_net_),
            .in1(N__33673),
            .in2(N__37785),
            .in3(_gnd_net_),
            .lcout(data_count_0),
            .ltout(),
            .carryin(bfn_12_18_0_),
            .carryout(n19765),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__37843),
            .sr(N__38139));
    defparam data_count_i0_i1_LC_12_18_1.C_ON=1'b1;
    defparam data_count_i0_i1_LC_12_18_1.SEQ_MODE=4'b1000;
    defparam data_count_i0_i1_LC_12_18_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i1_LC_12_18_1 (
            .in0(_gnd_net_),
            .in1(N__33571),
            .in2(_gnd_net_),
            .in3(N__33549),
            .lcout(data_count_1),
            .ltout(),
            .carryin(n19765),
            .carryout(n19766),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__37843),
            .sr(N__38139));
    defparam data_count_i0_i2_LC_12_18_2.C_ON=1'b1;
    defparam data_count_i0_i2_LC_12_18_2.SEQ_MODE=4'b1000;
    defparam data_count_i0_i2_LC_12_18_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i2_LC_12_18_2 (
            .in0(_gnd_net_),
            .in1(N__33460),
            .in2(_gnd_net_),
            .in3(N__33438),
            .lcout(data_count_2),
            .ltout(),
            .carryin(n19766),
            .carryout(n19767),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__37843),
            .sr(N__38139));
    defparam data_count_i0_i3_LC_12_18_3.C_ON=1'b1;
    defparam data_count_i0_i3_LC_12_18_3.SEQ_MODE=4'b1000;
    defparam data_count_i0_i3_LC_12_18_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i3_LC_12_18_3 (
            .in0(_gnd_net_),
            .in1(N__33349),
            .in2(_gnd_net_),
            .in3(N__33327),
            .lcout(data_count_3),
            .ltout(),
            .carryin(n19767),
            .carryout(n19768),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__37843),
            .sr(N__38139));
    defparam data_count_i0_i4_LC_12_18_4.C_ON=1'b1;
    defparam data_count_i0_i4_LC_12_18_4.SEQ_MODE=4'b1000;
    defparam data_count_i0_i4_LC_12_18_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i4_LC_12_18_4 (
            .in0(_gnd_net_),
            .in1(N__33247),
            .in2(_gnd_net_),
            .in3(N__33225),
            .lcout(data_count_4),
            .ltout(),
            .carryin(n19768),
            .carryout(n19769),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__37843),
            .sr(N__38139));
    defparam data_count_i0_i5_LC_12_18_5.C_ON=1'b1;
    defparam data_count_i0_i5_LC_12_18_5.SEQ_MODE=4'b1000;
    defparam data_count_i0_i5_LC_12_18_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i5_LC_12_18_5 (
            .in0(_gnd_net_),
            .in1(N__33142),
            .in2(_gnd_net_),
            .in3(N__33117),
            .lcout(data_count_5),
            .ltout(),
            .carryin(n19769),
            .carryout(n19770),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__37843),
            .sr(N__38139));
    defparam data_count_i0_i6_LC_12_18_6.C_ON=1'b1;
    defparam data_count_i0_i6_LC_12_18_6.SEQ_MODE=4'b1000;
    defparam data_count_i0_i6_LC_12_18_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i6_LC_12_18_6 (
            .in0(_gnd_net_),
            .in1(N__34153),
            .in2(_gnd_net_),
            .in3(N__34131),
            .lcout(data_count_6),
            .ltout(),
            .carryin(n19770),
            .carryout(n19771),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__37843),
            .sr(N__38139));
    defparam data_count_i0_i7_LC_12_18_7.C_ON=1'b1;
    defparam data_count_i0_i7_LC_12_18_7.SEQ_MODE=4'b1000;
    defparam data_count_i0_i7_LC_12_18_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i7_LC_12_18_7 (
            .in0(_gnd_net_),
            .in1(N__34045),
            .in2(_gnd_net_),
            .in3(N__34023),
            .lcout(data_count_7),
            .ltout(),
            .carryin(n19771),
            .carryout(n19772),
            .clk(INVdata_count_i0_i0C_net),
            .ce(N__37843),
            .sr(N__38139));
    defparam data_count_i0_i8_LC_12_19_0.C_ON=1'b1;
    defparam data_count_i0_i8_LC_12_19_0.SEQ_MODE=4'b1000;
    defparam data_count_i0_i8_LC_12_19_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i8_LC_12_19_0 (
            .in0(_gnd_net_),
            .in1(N__33937),
            .in2(_gnd_net_),
            .in3(N__33915),
            .lcout(data_count_8),
            .ltout(),
            .carryin(bfn_12_19_0_),
            .carryout(n19773),
            .clk(INVdata_count_i0_i8C_net),
            .ce(N__37845),
            .sr(N__38149));
    defparam data_count_i0_i9_LC_12_19_1.C_ON=1'b0;
    defparam data_count_i0_i9_LC_12_19_1.SEQ_MODE=4'b1000;
    defparam data_count_i0_i9_LC_12_19_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_count_i0_i9_LC_12_19_1 (
            .in0(_gnd_net_),
            .in1(N__33835),
            .in2(_gnd_net_),
            .in3(N__33912),
            .lcout(data_count_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVdata_count_i0_i8C_net),
            .ce(N__37845),
            .sr(N__38149));
    defparam \comm_spi.imosi_44_12287_12288_reset_LC_13_2_0 .C_ON=1'b0;
    defparam \comm_spi.imosi_44_12287_12288_reset_LC_13_2_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.imosi_44_12287_12288_reset_LC_13_2_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \comm_spi.imosi_44_12287_12288_reset_LC_13_2_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50884),
            .lcout(\comm_spi.n14809 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55937),
            .ce(),
            .sr(N__50832));
    defparam \comm_spi.data_rx_i0_12301_12302_reset_LC_13_3_0 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i0_12301_12302_reset_LC_13_3_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i0_12301_12302_reset_LC_13_3_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.data_rx_i0_12301_12302_reset_LC_13_3_0  (
            .in0(N__36911),
            .in1(N__36886),
            .in2(_gnd_net_),
            .in3(N__45032),
            .lcout(\comm_spi.n14823 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__58352),
            .ce(),
            .sr(N__39774));
    defparam \comm_spi.i19525_4_lut_3_lut_LC_13_4_0 .C_ON=1'b0;
    defparam \comm_spi.i19525_4_lut_3_lut_LC_13_4_0 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19525_4_lut_3_lut_LC_13_4_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \comm_spi.i19525_4_lut_3_lut_LC_13_4_0  (
            .in0(N__36970),
            .in1(N__50466),
            .in2(_gnd_net_),
            .in3(N__58121),
            .lcout(\comm_spi.n23083 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i19500_4_lut_3_lut_LC_13_4_5 .C_ON=1'b0;
    defparam \comm_spi.i19500_4_lut_3_lut_LC_13_4_5 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19500_4_lut_3_lut_LC_13_4_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \comm_spi.i19500_4_lut_3_lut_LC_13_4_5  (
            .in0(N__58120),
            .in1(N__33816),
            .in2(_gnd_net_),
            .in3(N__39785),
            .lcout(\comm_spi.n23089 ),
            .ltout(\comm_spi.n23089_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i12303_3_lut_LC_13_4_6 .C_ON=1'b0;
    defparam \comm_spi.i12303_3_lut_LC_13_4_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i12303_3_lut_LC_13_4_6 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \comm_spi.i12303_3_lut_LC_13_4_6  (
            .in0(_gnd_net_),
            .in1(N__34455),
            .in2(N__34449),
            .in3(N__34446),
            .lcout(comm_rx_buf_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.imosi_44_12287_12288_set_LC_13_5_0 .C_ON=1'b0;
    defparam \comm_spi.imosi_44_12287_12288_set_LC_13_5_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.imosi_44_12287_12288_set_LC_13_5_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \comm_spi.imosi_44_12287_12288_set_LC_13_5_0  (
            .in0(_gnd_net_),
            .in1(N__50892),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\comm_spi.n14808 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55938),
            .ce(),
            .sr(N__37158));
    defparam \ADC_VDC.bit_cnt_3771__i0_LC_13_6_0 .C_ON=1'b1;
    defparam \ADC_VDC.bit_cnt_3771__i0_LC_13_6_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3771__i0_LC_13_6_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3771__i0_LC_13_6_0  (
            .in0(_gnd_net_),
            .in1(N__34429),
            .in2(_gnd_net_),
            .in3(N__34404),
            .lcout(\ADC_VDC.bit_cnt_0 ),
            .ltout(),
            .carryin(bfn_13_6_0_),
            .carryout(\ADC_VDC.n19918 ),
            .clk(N__42221),
            .ce(N__51075),
            .sr(N__34737));
    defparam \ADC_VDC.bit_cnt_3771__i1_LC_13_6_1 .C_ON=1'b1;
    defparam \ADC_VDC.bit_cnt_3771__i1_LC_13_6_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3771__i1_LC_13_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3771__i1_LC_13_6_1  (
            .in0(_gnd_net_),
            .in1(N__34397),
            .in2(_gnd_net_),
            .in3(N__34377),
            .lcout(\ADC_VDC.bit_cnt_1 ),
            .ltout(),
            .carryin(\ADC_VDC.n19918 ),
            .carryout(\ADC_VDC.n19919 ),
            .clk(N__42221),
            .ce(N__51075),
            .sr(N__34737));
    defparam \ADC_VDC.bit_cnt_3771__i2_LC_13_6_2 .C_ON=1'b1;
    defparam \ADC_VDC.bit_cnt_3771__i2_LC_13_6_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3771__i2_LC_13_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3771__i2_LC_13_6_2  (
            .in0(_gnd_net_),
            .in1(N__34373),
            .in2(_gnd_net_),
            .in3(N__34341),
            .lcout(\ADC_VDC.bit_cnt_2 ),
            .ltout(),
            .carryin(\ADC_VDC.n19919 ),
            .carryout(\ADC_VDC.n19920 ),
            .clk(N__42221),
            .ce(N__51075),
            .sr(N__34737));
    defparam \ADC_VDC.bit_cnt_3771__i3_LC_13_6_3 .C_ON=1'b1;
    defparam \ADC_VDC.bit_cnt_3771__i3_LC_13_6_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3771__i3_LC_13_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3771__i3_LC_13_6_3  (
            .in0(_gnd_net_),
            .in1(N__34337),
            .in2(_gnd_net_),
            .in3(N__34308),
            .lcout(\ADC_VDC.bit_cnt_3 ),
            .ltout(),
            .carryin(\ADC_VDC.n19920 ),
            .carryout(\ADC_VDC.n19921 ),
            .clk(N__42221),
            .ce(N__51075),
            .sr(N__34737));
    defparam \ADC_VDC.bit_cnt_3771__i4_LC_13_6_4 .C_ON=1'b1;
    defparam \ADC_VDC.bit_cnt_3771__i4_LC_13_6_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3771__i4_LC_13_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3771__i4_LC_13_6_4  (
            .in0(_gnd_net_),
            .in1(N__34301),
            .in2(_gnd_net_),
            .in3(N__34278),
            .lcout(\ADC_VDC.bit_cnt_4 ),
            .ltout(),
            .carryin(\ADC_VDC.n19921 ),
            .carryout(\ADC_VDC.n19922 ),
            .clk(N__42221),
            .ce(N__51075),
            .sr(N__34737));
    defparam \ADC_VDC.bit_cnt_3771__i5_LC_13_6_5 .C_ON=1'b1;
    defparam \ADC_VDC.bit_cnt_3771__i5_LC_13_6_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3771__i5_LC_13_6_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3771__i5_LC_13_6_5  (
            .in0(_gnd_net_),
            .in1(N__34274),
            .in2(_gnd_net_),
            .in3(N__34257),
            .lcout(\ADC_VDC.bit_cnt_5 ),
            .ltout(),
            .carryin(\ADC_VDC.n19922 ),
            .carryout(\ADC_VDC.n19923 ),
            .clk(N__42221),
            .ce(N__51075),
            .sr(N__34737));
    defparam \ADC_VDC.bit_cnt_3771__i6_LC_13_6_6 .C_ON=1'b1;
    defparam \ADC_VDC.bit_cnt_3771__i6_LC_13_6_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3771__i6_LC_13_6_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3771__i6_LC_13_6_6  (
            .in0(_gnd_net_),
            .in1(N__34254),
            .in2(_gnd_net_),
            .in3(N__34239),
            .lcout(\ADC_VDC.bit_cnt_6 ),
            .ltout(),
            .carryin(\ADC_VDC.n19923 ),
            .carryout(\ADC_VDC.n19924 ),
            .clk(N__42221),
            .ce(N__51075),
            .sr(N__34737));
    defparam \ADC_VDC.bit_cnt_3771__i7_LC_13_6_7 .C_ON=1'b0;
    defparam \ADC_VDC.bit_cnt_3771__i7_LC_13_6_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.bit_cnt_3771__i7_LC_13_6_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.bit_cnt_3771__i7_LC_13_6_7  (
            .in0(_gnd_net_),
            .in1(N__34752),
            .in2(_gnd_net_),
            .in3(N__34755),
            .lcout(\ADC_VDC.bit_cnt_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42221),
            .ce(N__51075),
            .sr(N__34737));
    defparam i1_4_lut_adj_311_LC_13_7_0.C_ON=1'b0;
    defparam i1_4_lut_adj_311_LC_13_7_0.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_311_LC_13_7_0.LUT_INIT=16'b1010000010100010;
    LogicCell40 i1_4_lut_adj_311_LC_13_7_0 (
            .in0(N__55346),
            .in1(N__37182),
            .in2(N__49392),
            .in3(N__35460),
            .lcout(n12662),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i5_4_lut_adj_150_LC_13_7_1.C_ON=1'b0;
    defparam i5_4_lut_adj_150_LC_13_7_1.SEQ_MODE=4'b0000;
    defparam i5_4_lut_adj_150_LC_13_7_1.LUT_INIT=16'b0111110110111110;
    LogicCell40 i5_4_lut_adj_150_LC_13_7_1 (
            .in0(N__37929),
            .in1(N__40683),
            .in2(N__35214),
            .in3(N__34879),
            .lcout(n21_adj_1594),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12_4_lut_adj_58_LC_13_7_2.C_ON=1'b0;
    defparam i12_4_lut_adj_58_LC_13_7_2.SEQ_MODE=4'b0000;
    defparam i12_4_lut_adj_58_LC_13_7_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i12_4_lut_adj_58_LC_13_7_2 (
            .in0(N__39744),
            .in1(N__40002),
            .in2(N__40080),
            .in3(N__39966),
            .lcout(n31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam SecClk_292_LC_13_7_3.C_ON=1'b0;
    defparam SecClk_292_LC_13_7_3.SEQ_MODE=4'b1000;
    defparam SecClk_292_LC_13_7_3.LUT_INIT=16'b0101010110101010;
    LogicCell40 SecClk_292_LC_13_7_3 (
            .in0(N__34693),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34664),
            .lcout(TEST_LED),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50783),
            .ce(),
            .sr(_gnd_net_));
    defparam i9_4_lut_LC_13_7_4.C_ON=1'b0;
    defparam i9_4_lut_LC_13_7_4.SEQ_MODE=4'b0000;
    defparam i9_4_lut_LC_13_7_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i9_4_lut_LC_13_7_4 (
            .in0(N__34647),
            .in1(N__34629),
            .in2(N__34611),
            .in3(N__34593),
            .lcout(n25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12_4_lut_adj_198_LC_13_7_5.C_ON=1'b0;
    defparam i12_4_lut_adj_198_LC_13_7_5.SEQ_MODE=4'b0000;
    defparam i12_4_lut_adj_198_LC_13_7_5.LUT_INIT=16'b1111111111111110;
    LogicCell40 i12_4_lut_adj_198_LC_13_7_5 (
            .in0(N__34572),
            .in1(N__34553),
            .in2(N__34539),
            .in3(N__34518),
            .lcout(n28_adj_1554),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i8_4_lut_adj_146_LC_13_8_0.C_ON=1'b0;
    defparam i8_4_lut_adj_146_LC_13_8_0.SEQ_MODE=4'b0000;
    defparam i8_4_lut_adj_146_LC_13_8_0.LUT_INIT=16'b0111101111011110;
    LogicCell40 i8_4_lut_adj_146_LC_13_8_0 (
            .in0(N__37863),
            .in1(N__43086),
            .in2(N__34487),
            .in3(N__42994),
            .lcout(n24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19343_2_lut_LC_13_8_1.C_ON=1'b0;
    defparam i19343_2_lut_LC_13_8_1.SEQ_MODE=4'b0000;
    defparam i19343_2_lut_LC_13_8_1.LUT_INIT=16'b0011001100000000;
    LogicCell40 i19343_2_lut_LC_13_8_1 (
            .in0(_gnd_net_),
            .in1(N__57186),
            .in2(_gnd_net_),
            .in3(N__34880),
            .lcout(n21703),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_93_2_lut_LC_13_8_2 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_93_2_lut_LC_13_8_2 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_93_2_lut_LC_13_8_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \comm_spi.RESET_I_0_93_2_lut_LC_13_8_2  (
            .in0(N__50462),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58066),
            .lcout(\comm_spi.data_tx_7__N_807 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i12_LC_13_8_3.C_ON=1'b0;
    defparam req_data_cnt_i12_LC_13_8_3.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i12_LC_13_8_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 req_data_cnt_i12_LC_13_8_3 (
            .in0(N__37196),
            .in1(N__35508),
            .in2(_gnd_net_),
            .in3(N__34881),
            .lcout(req_data_cnt_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55943),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i9_LC_13_8_4.C_ON=1'b0;
    defparam req_data_cnt_i9_LC_13_8_4.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i9_LC_13_8_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 req_data_cnt_i9_LC_13_8_4 (
            .in0(N__35510),
            .in1(N__37445),
            .in2(_gnd_net_),
            .in3(N__42995),
            .lcout(req_data_cnt_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55943),
            .ce(),
            .sr(_gnd_net_));
    defparam i6_4_lut_adj_148_LC_13_8_5.C_ON=1'b0;
    defparam i6_4_lut_adj_148_LC_13_8_5.SEQ_MODE=4'b0000;
    defparam i6_4_lut_adj_148_LC_13_8_5.LUT_INIT=16'b0111101111011110;
    LogicCell40 i6_4_lut_adj_148_LC_13_8_5 (
            .in0(N__37725),
            .in1(N__46527),
            .in2(N__35374),
            .in3(N__46567),
            .lcout(n22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i19520_4_lut_3_lut_LC_13_8_6 .C_ON=1'b0;
    defparam \comm_spi.i19520_4_lut_3_lut_LC_13_8_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19520_4_lut_3_lut_LC_13_8_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \comm_spi.i19520_4_lut_3_lut_LC_13_8_6  (
            .in0(N__34804),
            .in1(N__53685),
            .in2(_gnd_net_),
            .in3(N__58067),
            .lcout(\comm_spi.n23095 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i2_LC_13_8_7.C_ON=1'b0;
    defparam req_data_cnt_i2_LC_13_8_7.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i2_LC_13_8_7.LUT_INIT=16'b1011100010111000;
    LogicCell40 req_data_cnt_i2_LC_13_8_7 (
            .in0(N__34851),
            .in1(N__35509),
            .in2(N__35375),
            .in3(_gnd_net_),
            .lcout(req_data_cnt_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55943),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i6_12325_12326_set_LC_13_9_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i6_12325_12326_set_LC_13_9_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i6_12325_12326_set_LC_13_9_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i6_12325_12326_set_LC_13_9_0  (
            .in0(N__34805),
            .in1(N__52631),
            .in2(_gnd_net_),
            .in3(N__57470),
            .lcout(\comm_spi.n14846 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__58401),
            .ce(),
            .sr(N__34788));
    defparam i19332_2_lut_LC_13_9_1.C_ON=1'b0;
    defparam i19332_2_lut_LC_13_9_1.SEQ_MODE=4'b0000;
    defparam i19332_2_lut_LC_13_9_1.LUT_INIT=16'b0011001100000000;
    LogicCell40 i19332_2_lut_LC_13_9_1 (
            .in0(_gnd_net_),
            .in1(N__57213),
            .in2(_gnd_net_),
            .in3(N__34776),
            .lcout(n21702),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19431_2_lut_LC_13_9_3.C_ON=1'b0;
    defparam i19431_2_lut_LC_13_9_3.SEQ_MODE=4'b0000;
    defparam i19431_2_lut_LC_13_9_3.LUT_INIT=16'b0011001100000000;
    LogicCell40 i19431_2_lut_LC_13_9_3 (
            .in0(_gnd_net_),
            .in1(N__35811),
            .in2(_gnd_net_),
            .in3(N__37035),
            .lcout(n14915),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_LC_13_9_4.C_ON=1'b0;
    defparam i2_2_lut_LC_13_9_4.SEQ_MODE=4'b0000;
    defparam i2_2_lut_LC_13_9_4.LUT_INIT=16'b1100110000000000;
    LogicCell40 i2_2_lut_LC_13_9_4 (
            .in0(_gnd_net_),
            .in1(N__35148),
            .in2(_gnd_net_),
            .in3(N__35130),
            .lcout(n10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_13_9_6.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_13_9_6.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_13_9_6.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_13_9_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19746_LC_13_10_0.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19746_LC_13_10_0.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19746_LC_13_10_0.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_19746_LC_13_10_0 (
            .in0(N__35109),
            .in1(N__46402),
            .in2(N__35094),
            .in3(N__47729),
            .lcout(n22485),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18442_2_lut_LC_13_10_1.C_ON=1'b0;
    defparam i18442_2_lut_LC_13_10_1.SEQ_MODE=4'b0000;
    defparam i18442_2_lut_LC_13_10_1.LUT_INIT=16'b1111111111001100;
    LogicCell40 i18442_2_lut_LC_13_10_1 (
            .in0(_gnd_net_),
            .in1(N__37570),
            .in2(_gnd_net_),
            .in3(N__53997),
            .lcout(n11652),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_3_i19_3_lut_LC_13_10_3.C_ON=1'b0;
    defparam mux_129_Mux_3_i19_3_lut_LC_13_10_3.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_3_i19_3_lut_LC_13_10_3.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_129_Mux_3_i19_3_lut_LC_13_10_3 (
            .in0(N__35076),
            .in1(N__35045),
            .in2(_gnd_net_),
            .in3(N__57099),
            .lcout(n19_adj_1641),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_4_i20_3_lut_LC_13_10_4.C_ON=1'b0;
    defparam mux_128_Mux_4_i20_3_lut_LC_13_10_4.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_4_i20_3_lut_LC_13_10_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_128_Mux_4_i20_3_lut_LC_13_10_4 (
            .in0(N__57098),
            .in1(N__35025),
            .in2(_gnd_net_),
            .in3(N__34998),
            .lcout(n20_adj_1674),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_287_LC_13_10_5.C_ON=1'b0;
    defparam i1_4_lut_adj_287_LC_13_10_5.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_287_LC_13_10_5.LUT_INIT=16'b1000100011001000;
    LogicCell40 i1_4_lut_adj_287_LC_13_10_5 (
            .in0(N__55207),
            .in1(N__55544),
            .in2(N__35280),
            .in3(N__54803),
            .lcout(n16821),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_5_i16_3_lut_LC_13_10_6.C_ON=1'b0;
    defparam mux_128_Mux_5_i16_3_lut_LC_13_10_6.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_5_i16_3_lut_LC_13_10_6.LUT_INIT=16'b1111101001010000;
    LogicCell40 mux_128_Mux_5_i16_3_lut_LC_13_10_6 (
            .in0(N__57101),
            .in1(_gnd_net_),
            .in2(N__35309),
            .in3(N__34971),
            .lcout(n16_adj_1664),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_5_i20_3_lut_LC_13_10_7.C_ON=1'b0;
    defparam mux_128_Mux_5_i20_3_lut_LC_13_10_7.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_5_i20_3_lut_LC_13_10_7.LUT_INIT=16'b1100110010101010;
    LogicCell40 mux_128_Mux_5_i20_3_lut_LC_13_10_7 (
            .in0(N__34918),
            .in1(N__34902),
            .in2(_gnd_net_),
            .in3(N__57100),
            .lcout(n20_adj_1667),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_4_lut_adj_263_LC_13_11_0.C_ON=1'b0;
    defparam i1_3_lut_4_lut_adj_263_LC_13_11_0.SEQ_MODE=4'b0000;
    defparam i1_3_lut_4_lut_adj_263_LC_13_11_0.LUT_INIT=16'b1111111100011111;
    LogicCell40 i1_3_lut_4_lut_adj_263_LC_13_11_0 (
            .in0(N__54517),
            .in1(N__48237),
            .in2(N__54788),
            .in3(N__55298),
            .lcout(),
            .ltout(n12082_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_189_LC_13_11_1.C_ON=1'b0;
    defparam i1_4_lut_adj_189_LC_13_11_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_189_LC_13_11_1.LUT_INIT=16'b1110000000000000;
    LogicCell40 i1_4_lut_adj_189_LC_13_11_1 (
            .in0(N__35279),
            .in1(N__48341),
            .in2(N__35256),
            .in3(N__55562),
            .lcout(n12089),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i6_LC_13_11_2.C_ON=1'b0;
    defparam comm_cmd_i6_LC_13_11_2.SEQ_MODE=4'b1000;
    defparam comm_cmd_i6_LC_13_11_2.LUT_INIT=16'b1011001110000000;
    LogicCell40 comm_cmd_i6_LC_13_11_2 (
            .in0(N__50952),
            .in1(N__37496),
            .in2(N__53235),
            .in3(N__48851),
            .lcout(comm_cmd_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55958),
            .ce(),
            .sr(_gnd_net_));
    defparam i15463_2_lut_3_lut_LC_13_11_3.C_ON=1'b0;
    defparam i15463_2_lut_3_lut_LC_13_11_3.SEQ_MODE=4'b0000;
    defparam i15463_2_lut_3_lut_LC_13_11_3.LUT_INIT=16'b0000000000100010;
    LogicCell40 i15463_2_lut_3_lut_LC_13_11_3 (
            .in0(N__45302),
            .in1(N__54710),
            .in2(_gnd_net_),
            .in3(N__54518),
            .lcout(n14_adj_1573),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_101_2_lut_LC_13_11_4 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_101_2_lut_LC_13_11_4 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_101_2_lut_LC_13_11_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \comm_spi.RESET_I_0_101_2_lut_LC_13_11_4  (
            .in0(N__50455),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58065),
            .lcout(\comm_spi.data_tx_7__N_817 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_2_i24_3_lut_LC_13_11_5.C_ON=1'b0;
    defparam mux_128_Mux_2_i24_3_lut_LC_13_11_5.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_2_i24_3_lut_LC_13_11_5.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_128_Mux_2_i24_3_lut_LC_13_11_5 (
            .in0(N__35736),
            .in1(N__57163),
            .in2(_gnd_net_),
            .in3(N__35210),
            .lcout(n24_adj_1686),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_300_LC_13_11_6.C_ON=1'b0;
    defparam i1_2_lut_adj_300_LC_13_11_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_300_LC_13_11_6.LUT_INIT=16'b1111111110101010;
    LogicCell40 i1_2_lut_adj_300_LC_13_11_6 (
            .in0(N__54706),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55297),
            .lcout(n12442),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_i7_LC_13_11_7.C_ON=1'b0;
    defparam comm_cmd_i7_LC_13_11_7.SEQ_MODE=4'b1000;
    defparam comm_cmd_i7_LC_13_11_7.LUT_INIT=16'b1101010110000000;
    LogicCell40 comm_cmd_i7_LC_13_11_7 (
            .in0(N__37497),
            .in1(N__50953),
            .in2(N__48598),
            .in3(N__49993),
            .lcout(comm_cmd_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55958),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_LC_13_12_0.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_LC_13_12_0.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_LC_13_12_0.LUT_INIT=16'b1111010110001000;
    LogicCell40 comm_cmd_1__bdd_4_lut_LC_13_12_0 (
            .in0(N__47675),
            .in1(N__35187),
            .in2(N__35175),
            .in3(N__46465),
            .lcout(),
            .ltout(n22641_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22641_bdd_4_lut_LC_13_12_1.C_ON=1'b0;
    defparam n22641_bdd_4_lut_LC_13_12_1.SEQ_MODE=4'b0000;
    defparam n22641_bdd_4_lut_LC_13_12_1.LUT_INIT=16'b1111000010101100;
    LogicCell40 n22641_bdd_4_lut_LC_13_12_1 (
            .in0(N__38238),
            .in1(N__35442),
            .in2(N__35430),
            .in3(N__47676),
            .lcout(n22644),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_2_i26_3_lut_LC_13_12_2.C_ON=1'b0;
    defparam mux_129_Mux_2_i26_3_lut_LC_13_12_2.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_2_i26_3_lut_LC_13_12_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_129_Mux_2_i26_3_lut_LC_13_12_2 (
            .in0(N__35427),
            .in1(N__57195),
            .in2(_gnd_net_),
            .in3(N__37717),
            .lcout(),
            .ltout(n26_adj_1647_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19673_LC_13_12_3.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19673_LC_13_12_3.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19673_LC_13_12_3.LUT_INIT=16'b1101100010101010;
    LogicCell40 comm_cmd_1__bdd_4_lut_19673_LC_13_12_3 (
            .in0(N__46466),
            .in1(N__42570),
            .in2(N__35403),
            .in3(N__47677),
            .lcout(),
            .ltout(n22383_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22383_bdd_4_lut_LC_13_12_4.C_ON=1'b0;
    defparam n22383_bdd_4_lut_LC_13_12_4.SEQ_MODE=4'b0000;
    defparam n22383_bdd_4_lut_LC_13_12_4.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22383_bdd_4_lut_LC_13_12_4 (
            .in0(N__47678),
            .in1(N__35400),
            .in2(N__35379),
            .in3(N__35376),
            .lcout(),
            .ltout(n22386_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1568256_i1_3_lut_LC_13_12_5.C_ON=1'b0;
    defparam i1568256_i1_3_lut_LC_13_12_5.SEQ_MODE=4'b0000;
    defparam i1568256_i1_3_lut_LC_13_12_5.LUT_INIT=16'b1110010011100100;
    LogicCell40 i1568256_i1_3_lut_LC_13_12_5 (
            .in0(N__47233),
            .in1(N__35352),
            .in2(N__35346),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(n30_adj_1648_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i2_LC_13_12_6.C_ON=1'b0;
    defparam comm_buf_1__i2_LC_13_12_6.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i2_LC_13_12_6.LUT_INIT=16'b1010101011110000;
    LogicCell40 comm_buf_1__i2_LC_13_12_6 (
            .in0(N__50158),
            .in1(_gnd_net_),
            .in2(N__35343),
            .in3(N__54499),
            .lcout(comm_buf_1_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55967),
            .ce(N__45195),
            .sr(N__44002));
    defparam i2_3_lut_adj_266_LC_13_12_7.C_ON=1'b0;
    defparam i2_3_lut_adj_266_LC_13_12_7.SEQ_MODE=4'b0000;
    defparam i2_3_lut_adj_266_LC_13_12_7.LUT_INIT=16'b1111111111101110;
    LogicCell40 i2_3_lut_adj_266_LC_13_12_7 (
            .in0(N__47232),
            .in1(N__46290),
            .in2(_gnd_net_),
            .in3(N__47674),
            .lcout(n66),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_adj_154_LC_13_13_0.C_ON=1'b0;
    defparam i2_4_lut_adj_154_LC_13_13_0.SEQ_MODE=4'b0000;
    defparam i2_4_lut_adj_154_LC_13_13_0.LUT_INIT=16'b0111110110111110;
    LogicCell40 i2_4_lut_adj_154_LC_13_13_0 (
            .in0(N__44194),
            .in1(N__37690),
            .in2(N__35340),
            .in3(N__44140),
            .lcout(n18_adj_1644),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i13_LC_13_13_1.C_ON=1'b0;
    defparam buf_dds0_i13_LC_13_13_1.SEQ_MODE=4'b1000;
    defparam buf_dds0_i13_LC_13_13_1.LUT_INIT=16'b0011000010101010;
    LogicCell40 buf_dds0_i13_LC_13_13_1 (
            .in0(N__35299),
            .in1(N__49311),
            .in2(N__52276),
            .in3(N__41644),
            .lcout(buf_dds0_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55978),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_adj_267_LC_13_13_2.C_ON=1'b0;
    defparam i2_3_lut_adj_267_LC_13_13_2.SEQ_MODE=4'b0000;
    defparam i2_3_lut_adj_267_LC_13_13_2.LUT_INIT=16'b1111111111101110;
    LogicCell40 i2_3_lut_adj_267_LC_13_13_2 (
            .in0(N__35643),
            .in1(N__48259),
            .in2(_gnd_net_),
            .in3(N__57146),
            .lcout(n20011),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i14_LC_13_13_3.C_ON=1'b0;
    defparam buf_dds1_i14_LC_13_13_3.SEQ_MODE=4'b1000;
    defparam buf_dds1_i14_LC_13_13_3.LUT_INIT=16'b1100101000000000;
    LogicCell40 buf_dds1_i14_LC_13_13_3 (
            .in0(N__35629),
            .in1(N__49537),
            .in2(N__46910),
            .in3(N__46764),
            .lcout(buf_dds1_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55978),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i7_LC_13_13_5.C_ON=1'b0;
    defparam buf_dds1_i7_LC_13_13_5.SEQ_MODE=4'b1000;
    defparam buf_dds1_i7_LC_13_13_5.LUT_INIT=16'b1110010000000000;
    LogicCell40 buf_dds1_i7_LC_13_13_5 (
            .in0(N__46890),
            .in1(N__36568),
            .in2(N__44078),
            .in3(N__46765),
            .lcout(buf_dds1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55978),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i1_LC_13_13_6.C_ON=1'b0;
    defparam buf_dds1_i1_LC_13_13_6.SEQ_MODE=4'b1000;
    defparam buf_dds1_i1_LC_13_13_6.LUT_INIT=16'b1000100010100000;
    LogicCell40 buf_dds1_i1_LC_13_13_6 (
            .in0(N__46763),
            .in1(N__53510),
            .in2(N__35602),
            .in3(N__46894),
            .lcout(buf_dds1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55978),
            .ce(),
            .sr(_gnd_net_));
    defparam req_data_cnt_i1_LC_13_13_7.C_ON=1'b0;
    defparam req_data_cnt_i1_LC_13_13_7.SEQ_MODE=4'b1000;
    defparam req_data_cnt_i1_LC_13_13_7.LUT_INIT=16'b1111000010101010;
    LogicCell40 req_data_cnt_i1_LC_13_13_7 (
            .in0(N__44141),
            .in1(_gnd_net_),
            .in2(N__36166),
            .in3(N__35555),
            .lcout(req_data_cnt_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55978),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i1_LC_13_14_0.C_ON=1'b0;
    defparam buf_control_i1_LC_13_14_0.SEQ_MODE=4'b1000;
    defparam buf_control_i1_LC_13_14_0.LUT_INIT=16'b0011101100001000;
    LogicCell40 buf_control_i1_LC_13_14_0 (
            .in0(N__53436),
            .in1(N__41989),
            .in2(N__49361),
            .in3(N__42937),
            .lcout(DDS_RNG_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55991),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_271_LC_13_14_2.C_ON=1'b0;
    defparam i1_4_lut_adj_271_LC_13_14_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_271_LC_13_14_2.LUT_INIT=16'b1101110000000000;
    LogicCell40 i1_4_lut_adj_271_LC_13_14_2 (
            .in0(N__48266),
            .in1(N__49272),
            .in2(N__35478),
            .in3(N__55455),
            .lcout(n12144),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_4_lut_LC_13_14_3.C_ON=1'b0;
    defparam i2_2_lut_4_lut_LC_13_14_3.SEQ_MODE=4'b0000;
    defparam i2_2_lut_4_lut_LC_13_14_3.LUT_INIT=16'b1111111111110111;
    LogicCell40 i2_2_lut_4_lut_LC_13_14_3 (
            .in0(N__46377),
            .in1(N__47643),
            .in2(N__57209),
            .in3(N__53988),
            .lcout(n7_adj_1650),
            .ltout(n7_adj_1650_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_4_lut_adj_283_LC_13_14_4.C_ON=1'b0;
    defparam i3_4_lut_adj_283_LC_13_14_4.SEQ_MODE=4'b0000;
    defparam i3_4_lut_adj_283_LC_13_14_4.LUT_INIT=16'b1111111111111101;
    LogicCell40 i3_4_lut_adj_283_LC_13_14_4 (
            .in0(N__54738),
            .in1(N__54487),
            .in2(N__35463),
            .in3(N__35456),
            .lcout(n10756),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i3_LC_13_14_5.C_ON=1'b0;
    defparam buf_control_i3_LC_13_14_5.SEQ_MODE=4'b1000;
    defparam buf_control_i3_LC_13_14_5.LUT_INIT=16'b0101110100001000;
    LogicCell40 buf_control_i3_LC_13_14_5 (
            .in0(N__41988),
            .in1(N__45326),
            .in2(N__49355),
            .in3(N__36215),
            .lcout(SELIRNG1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55991),
            .ce(),
            .sr(_gnd_net_));
    defparam i15465_2_lut_3_lut_LC_13_14_6.C_ON=1'b0;
    defparam i15465_2_lut_3_lut_LC_13_14_6.SEQ_MODE=4'b0000;
    defparam i15465_2_lut_3_lut_LC_13_14_6.LUT_INIT=16'b0000000001000100;
    LogicCell40 i15465_2_lut_3_lut_LC_13_14_6 (
            .in0(N__54740),
            .in1(N__42710),
            .in2(_gnd_net_),
            .in3(N__54489),
            .lcout(n14_adj_1546),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15468_2_lut_3_lut_LC_13_14_7.C_ON=1'b0;
    defparam i15468_2_lut_3_lut_LC_13_14_7.SEQ_MODE=4'b0000;
    defparam i15468_2_lut_3_lut_LC_13_14_7.LUT_INIT=16'b0000000001000100;
    LogicCell40 i15468_2_lut_3_lut_LC_13_14_7 (
            .in0(N__54488),
            .in1(N__53511),
            .in2(_gnd_net_),
            .in3(N__54739),
            .lcout(n14_adj_1549),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_354_Mux_6_i15_4_lut_LC_13_15_0.C_ON=1'b0;
    defparam comm_state_3__I_0_354_Mux_6_i15_4_lut_LC_13_15_0.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_354_Mux_6_i15_4_lut_LC_13_15_0.LUT_INIT=16'b0111001001010000;
    LogicCell40 comm_state_3__I_0_354_Mux_6_i15_4_lut_LC_13_15_0 (
            .in0(N__55436),
            .in1(N__49209),
            .in2(N__38034),
            .in3(N__36128),
            .lcout(data_index_9_N_212_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_78_LC_13_15_1.C_ON=1'b0;
    defparam i1_4_lut_adj_78_LC_13_15_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_78_LC_13_15_1.LUT_INIT=16'b0111110110111110;
    LogicCell40 i1_4_lut_adj_78_LC_13_15_1 (
            .in0(N__36546),
            .in1(N__43534),
            .in2(N__36846),
            .in3(N__43672),
            .lcout(n17_adj_1553),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i5_LC_13_15_2.C_ON=1'b0;
    defparam buf_control_i5_LC_13_15_2.SEQ_MODE=4'b1000;
    defparam buf_control_i5_LC_13_15_2.LUT_INIT=16'b0010001011110000;
    LogicCell40 buf_control_i5_LC_13_15_2 (
            .in0(N__52277),
            .in1(N__49215),
            .in2(N__35989),
            .in3(N__41990),
            .lcout(AMPV_POW),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56005),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_256_LC_13_15_3.C_ON=1'b0;
    defparam i1_4_lut_adj_256_LC_13_15_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_256_LC_13_15_3.LUT_INIT=16'b1011101100001011;
    LogicCell40 i1_4_lut_adj_256_LC_13_15_3 (
            .in0(N__55563),
            .in1(N__36513),
            .in2(N__49317),
            .in3(N__55438),
            .lcout(n11611),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_354_Mux_3_i15_4_lut_LC_13_15_4.C_ON=1'b0;
    defparam comm_state_3__I_0_354_Mux_3_i15_4_lut_LC_13_15_4.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_354_Mux_3_i15_4_lut_LC_13_15_4.LUT_INIT=16'b0111010100100000;
    LogicCell40 comm_state_3__I_0_354_Mux_3_i15_4_lut_LC_13_15_4 (
            .in0(N__55435),
            .in1(N__49208),
            .in2(N__36237),
            .in3(N__38078),
            .lcout(data_index_9_N_212_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19459_2_lut_3_lut_LC_13_15_5.C_ON=1'b0;
    defparam i19459_2_lut_3_lut_LC_13_15_5.SEQ_MODE=4'b0000;
    defparam i19459_2_lut_3_lut_LC_13_15_5.LUT_INIT=16'b0000000000010001;
    LogicCell40 i19459_2_lut_3_lut_LC_13_15_5 (
            .in0(N__35880),
            .in1(N__35807),
            .in2(_gnd_net_),
            .in3(N__35710),
            .lcout(n21226),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i2_LC_13_15_6.C_ON=1'b0;
    defparam buf_control_i2_LC_13_15_6.SEQ_MODE=4'b1000;
    defparam buf_control_i2_LC_13_15_6.LUT_INIT=16'b0011000010101010;
    LogicCell40 buf_control_i2_LC_13_15_6 (
            .in0(N__45718),
            .in1(N__49214),
            .in2(N__45869),
            .in3(N__41991),
            .lcout(SELIRNG0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56005),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_268_LC_13_15_7.C_ON=1'b0;
    defparam i1_3_lut_adj_268_LC_13_15_7.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_268_LC_13_15_7.LUT_INIT=16'b1011101100000000;
    LogicCell40 i1_3_lut_adj_268_LC_13_15_7 (
            .in0(N__49210),
            .in1(N__36512),
            .in2(_gnd_net_),
            .in3(N__55437),
            .lcout(n12596),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_1_i22_3_lut_LC_13_16_0.C_ON=1'b0;
    defparam mux_130_Mux_1_i22_3_lut_LC_13_16_0.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_1_i22_3_lut_LC_13_16_0.LUT_INIT=16'b1100110010101010;
    LogicCell40 mux_130_Mux_1_i22_3_lut_LC_13_16_0 (
            .in0(N__36301),
            .in1(N__36501),
            .in2(_gnd_net_),
            .in3(N__47733),
            .lcout(n22_adj_1617),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15466_2_lut_3_lut_LC_13_16_1.C_ON=1'b0;
    defparam i15466_2_lut_3_lut_LC_13_16_1.SEQ_MODE=4'b0000;
    defparam i15466_2_lut_3_lut_LC_13_16_1.LUT_INIT=16'b0000000001000100;
    LogicCell40 i15466_2_lut_3_lut_LC_13_16_1 (
            .in0(N__54553),
            .in1(N__45282),
            .in2(_gnd_net_),
            .in3(N__54826),
            .lcout(n14_adj_1547),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6344_3_lut_LC_13_16_2.C_ON=1'b0;
    defparam i6344_3_lut_LC_13_16_2.SEQ_MODE=4'b0000;
    defparam i6344_3_lut_LC_13_16_2.LUT_INIT=16'b1100110010101010;
    LogicCell40 i6344_3_lut_LC_13_16_2 (
            .in0(N__42708),
            .in1(N__38182),
            .in2(_gnd_net_),
            .in3(N__41101),
            .lcout(n8_adj_1564),
            .ltout(n8_adj_1564_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_354_Mux_4_i15_4_lut_LC_13_16_3.C_ON=1'b0;
    defparam comm_state_3__I_0_354_Mux_4_i15_4_lut_LC_13_16_3.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_354_Mux_4_i15_4_lut_LC_13_16_3.LUT_INIT=16'b0111001101000000;
    LogicCell40 comm_state_3__I_0_354_Mux_4_i15_4_lut_LC_13_16_3 (
            .in0(N__49132),
            .in1(N__55439),
            .in2(N__36441),
            .in3(N__38195),
            .lcout(data_index_9_N_212_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i1_LC_13_16_4 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i1_LC_13_16_4 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i1_LC_13_16_4 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \ADC_IAC.ADC_DATA_i1_LC_13_16_4  (
            .in0(N__36302),
            .in1(N__38749),
            .in2(N__36351),
            .in3(N__38601),
            .lcout(buf_adcdata_iac_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56022),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_4_i16_3_lut_LC_13_16_5.C_ON=1'b0;
    defparam mux_128_Mux_4_i16_3_lut_LC_13_16_5.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_4_i16_3_lut_LC_13_16_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_128_Mux_4_i16_3_lut_LC_13_16_5 (
            .in0(N__36288),
            .in1(N__36258),
            .in2(_gnd_net_),
            .in3(N__57239),
            .lcout(n16_adj_1671),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6354_3_lut_LC_13_16_6.C_ON=1'b0;
    defparam i6354_3_lut_LC_13_16_6.SEQ_MODE=4'b0000;
    defparam i6354_3_lut_LC_13_16_6.LUT_INIT=16'b1100110010101010;
    LogicCell40 i6354_3_lut_LC_13_16_6 (
            .in0(N__45281),
            .in1(N__38096),
            .in2(_gnd_net_),
            .in3(N__41100),
            .lcout(n8_adj_1566),
            .ltout(n8_adj_1566_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i3_LC_13_16_7.C_ON=1'b0;
    defparam data_index_i3_LC_13_16_7.SEQ_MODE=4'b1000;
    defparam data_index_i3_LC_13_16_7.LUT_INIT=16'b0111001101000000;
    LogicCell40 data_index_i3_LC_13_16_7 (
            .in0(N__49133),
            .in1(N__55440),
            .in2(N__36636),
            .in3(N__38079),
            .lcout(data_index_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56022),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.tmp_buf_i7_LC_13_17_0 .C_ON=1'b0;
    defparam \SIG_DDS.tmp_buf_i7_LC_13_17_0 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.tmp_buf_i7_LC_13_17_0 .LUT_INIT=16'b0000110010101010;
    LogicCell40 \SIG_DDS.tmp_buf_i7_LC_13_17_0  (
            .in0(N__38789),
            .in1(N__36633),
            .in2(N__44491),
            .in3(N__44629),
            .lcout(\SIG_DDS.tmp_buf_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56036),
            .ce(N__43903),
            .sr(_gnd_net_));
    defparam \SIG_DDS.i23_4_lut_LC_13_17_2 .C_ON=1'b0;
    defparam \SIG_DDS.i23_4_lut_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \SIG_DDS.i23_4_lut_LC_13_17_2 .LUT_INIT=16'b1111101000010101;
    LogicCell40 \SIG_DDS.i23_4_lut_LC_13_17_2  (
            .in0(N__44445),
            .in1(N__43926),
            .in2(N__44753),
            .in3(N__44628),
            .lcout(\SIG_DDS.n9_adj_1434 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.i19478_4_lut_LC_13_17_3 .C_ON=1'b0;
    defparam \SIG_DDS.i19478_4_lut_LC_13_17_3 .SEQ_MODE=4'b0000;
    defparam \SIG_DDS.i19478_4_lut_LC_13_17_3 .LUT_INIT=16'b1111111110111110;
    LogicCell40 \SIG_DDS.i19478_4_lut_LC_13_17_3  (
            .in0(N__44626),
            .in1(N__44744),
            .in2(N__43936),
            .in3(N__44444),
            .lcout(\SIG_DDS.n9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.i19199_2_lut_LC_13_17_4 .C_ON=1'b0;
    defparam \SIG_DDS.i19199_2_lut_LC_13_17_4 .SEQ_MODE=4'b0000;
    defparam \SIG_DDS.i19199_2_lut_LC_13_17_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \SIG_DDS.i19199_2_lut_LC_13_17_4  (
            .in0(_gnd_net_),
            .in1(N__36612),
            .in2(_gnd_net_),
            .in3(N__44627),
            .lcout(\SIG_DDS.n21744 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_7_i16_3_lut_LC_13_17_5.C_ON=1'b0;
    defparam mux_129_Mux_7_i16_3_lut_LC_13_17_5.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_7_i16_3_lut_LC_13_17_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_129_Mux_7_i16_3_lut_LC_13_17_5 (
            .in0(N__36569),
            .in1(N__38788),
            .in2(_gnd_net_),
            .in3(N__57238),
            .lcout(n16_adj_1620),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipcnt_i0_i0_LC_13_18_0.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i0_LC_13_18_0.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i0_LC_13_18_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i0_LC_13_18_0 (
            .in0(_gnd_net_),
            .in1(N__37772),
            .in2(N__36545),
            .in3(_gnd_net_),
            .lcout(acadc_skipcnt_0),
            .ltout(),
            .carryin(bfn_13_18_0_),
            .carryout(n19789),
            .clk(INVacadc_skipcnt_i0_i0C_net),
            .ce(N__37043),
            .sr(N__36525));
    defparam add_73_2_THRU_CRY_0_LC_13_18_1.C_ON=1'b1;
    defparam add_73_2_THRU_CRY_0_LC_13_18_1.SEQ_MODE=4'b0000;
    defparam add_73_2_THRU_CRY_0_LC_13_18_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_73_2_THRU_CRY_0_LC_13_18_1 (
            .in0(_gnd_net_),
            .in1(N__58702),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n19789),
            .carryout(n19789_THRU_CRY_0_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_73_2_THRU_CRY_1_LC_13_18_2.C_ON=1'b1;
    defparam add_73_2_THRU_CRY_1_LC_13_18_2.SEQ_MODE=4'b0000;
    defparam add_73_2_THRU_CRY_1_LC_13_18_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_73_2_THRU_CRY_1_LC_13_18_2 (
            .in0(_gnd_net_),
            .in1(N__58706),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n19789_THRU_CRY_0_THRU_CO),
            .carryout(n19789_THRU_CRY_1_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_73_2_THRU_CRY_2_LC_13_18_3.C_ON=1'b1;
    defparam add_73_2_THRU_CRY_2_LC_13_18_3.SEQ_MODE=4'b0000;
    defparam add_73_2_THRU_CRY_2_LC_13_18_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_73_2_THRU_CRY_2_LC_13_18_3 (
            .in0(_gnd_net_),
            .in1(N__58703),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n19789_THRU_CRY_1_THRU_CO),
            .carryout(n19789_THRU_CRY_2_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_73_2_THRU_CRY_3_LC_13_18_4.C_ON=1'b1;
    defparam add_73_2_THRU_CRY_3_LC_13_18_4.SEQ_MODE=4'b0000;
    defparam add_73_2_THRU_CRY_3_LC_13_18_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_73_2_THRU_CRY_3_LC_13_18_4 (
            .in0(_gnd_net_),
            .in1(N__58707),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n19789_THRU_CRY_2_THRU_CO),
            .carryout(n19789_THRU_CRY_3_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_73_2_THRU_CRY_4_LC_13_18_5.C_ON=1'b1;
    defparam add_73_2_THRU_CRY_4_LC_13_18_5.SEQ_MODE=4'b0000;
    defparam add_73_2_THRU_CRY_4_LC_13_18_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_73_2_THRU_CRY_4_LC_13_18_5 (
            .in0(_gnd_net_),
            .in1(N__58704),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n19789_THRU_CRY_3_THRU_CO),
            .carryout(n19789_THRU_CRY_4_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_73_2_THRU_CRY_5_LC_13_18_6.C_ON=1'b1;
    defparam add_73_2_THRU_CRY_5_LC_13_18_6.SEQ_MODE=4'b0000;
    defparam add_73_2_THRU_CRY_5_LC_13_18_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_73_2_THRU_CRY_5_LC_13_18_6 (
            .in0(_gnd_net_),
            .in1(N__58708),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n19789_THRU_CRY_4_THRU_CO),
            .carryout(n19789_THRU_CRY_5_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_73_2_THRU_CRY_6_LC_13_18_7.C_ON=1'b1;
    defparam add_73_2_THRU_CRY_6_LC_13_18_7.SEQ_MODE=4'b0000;
    defparam add_73_2_THRU_CRY_6_LC_13_18_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 add_73_2_THRU_CRY_6_LC_13_18_7 (
            .in0(_gnd_net_),
            .in1(N__58705),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(n19789_THRU_CRY_5_THRU_CO),
            .carryout(n19789_THRU_CRY_6_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipcnt_i0_i1_LC_13_19_0.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i1_LC_13_19_0.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i1_LC_13_19_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i1_LC_13_19_0 (
            .in0(_gnd_net_),
            .in1(N__36719),
            .in2(_gnd_net_),
            .in3(N__36705),
            .lcout(acadc_skipcnt_1),
            .ltout(),
            .carryin(bfn_13_19_0_),
            .carryout(n19790),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__37042),
            .sr(N__36999));
    defparam acadc_skipcnt_i0_i2_LC_13_19_1.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i2_LC_13_19_1.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i2_LC_13_19_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i2_LC_13_19_1 (
            .in0(_gnd_net_),
            .in1(N__36698),
            .in2(_gnd_net_),
            .in3(N__36684),
            .lcout(acadc_skipcnt_2),
            .ltout(),
            .carryin(n19790),
            .carryout(n19791),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__37042),
            .sr(N__36999));
    defparam acadc_skipcnt_i0_i3_LC_13_19_2.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i3_LC_13_19_2.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i3_LC_13_19_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i3_LC_13_19_2 (
            .in0(_gnd_net_),
            .in1(N__36680),
            .in2(_gnd_net_),
            .in3(N__36663),
            .lcout(acadc_skipcnt_3),
            .ltout(),
            .carryin(n19791),
            .carryout(n19792),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__37042),
            .sr(N__36999));
    defparam acadc_skipcnt_i0_i4_LC_13_19_3.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i4_LC_13_19_3.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i4_LC_13_19_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i4_LC_13_19_3 (
            .in0(_gnd_net_),
            .in1(N__36653),
            .in2(_gnd_net_),
            .in3(N__36639),
            .lcout(acadc_skipcnt_4),
            .ltout(),
            .carryin(n19792),
            .carryout(n19793),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__37042),
            .sr(N__36999));
    defparam acadc_skipcnt_i0_i5_LC_13_19_4.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i5_LC_13_19_4.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i5_LC_13_19_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i5_LC_13_19_4 (
            .in0(_gnd_net_),
            .in1(N__36863),
            .in2(_gnd_net_),
            .in3(N__36849),
            .lcout(acadc_skipcnt_5),
            .ltout(),
            .carryin(n19793),
            .carryout(n19794),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__37042),
            .sr(N__36999));
    defparam acadc_skipcnt_i0_i6_LC_13_19_5.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i6_LC_13_19_5.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i6_LC_13_19_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i6_LC_13_19_5 (
            .in0(_gnd_net_),
            .in1(N__36842),
            .in2(_gnd_net_),
            .in3(N__36828),
            .lcout(acadc_skipcnt_6),
            .ltout(),
            .carryin(n19794),
            .carryout(n19795),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__37042),
            .sr(N__36999));
    defparam acadc_skipcnt_i0_i7_LC_13_19_6.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i7_LC_13_19_6.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i7_LC_13_19_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i7_LC_13_19_6 (
            .in0(_gnd_net_),
            .in1(N__36818),
            .in2(_gnd_net_),
            .in3(N__36804),
            .lcout(acadc_skipcnt_7),
            .ltout(),
            .carryin(n19795),
            .carryout(n19796),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__37042),
            .sr(N__36999));
    defparam acadc_skipcnt_i0_i8_LC_13_19_7.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i8_LC_13_19_7.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i8_LC_13_19_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i8_LC_13_19_7 (
            .in0(_gnd_net_),
            .in1(N__36797),
            .in2(_gnd_net_),
            .in3(N__36783),
            .lcout(acadc_skipcnt_8),
            .ltout(),
            .carryin(n19796),
            .carryout(n19797),
            .clk(INVacadc_skipcnt_i0_i1C_net),
            .ce(N__37042),
            .sr(N__36999));
    defparam acadc_skipcnt_i0_i9_LC_13_20_0.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i9_LC_13_20_0.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i9_LC_13_20_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i9_LC_13_20_0 (
            .in0(_gnd_net_),
            .in1(N__36776),
            .in2(_gnd_net_),
            .in3(N__36762),
            .lcout(acadc_skipcnt_9),
            .ltout(),
            .carryin(bfn_13_20_0_),
            .carryout(n19798),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__37044),
            .sr(N__36998));
    defparam acadc_skipcnt_i0_i10_LC_13_20_1.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i10_LC_13_20_1.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i10_LC_13_20_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i10_LC_13_20_1 (
            .in0(_gnd_net_),
            .in1(N__50663),
            .in2(_gnd_net_),
            .in3(N__36759),
            .lcout(acadc_skipcnt_10),
            .ltout(),
            .carryin(n19798),
            .carryout(n19799),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__37044),
            .sr(N__36998));
    defparam acadc_skipcnt_i0_i11_LC_13_20_2.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i11_LC_13_20_2.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i11_LC_13_20_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i11_LC_13_20_2 (
            .in0(_gnd_net_),
            .in1(N__36746),
            .in2(_gnd_net_),
            .in3(N__36732),
            .lcout(acadc_skipcnt_11),
            .ltout(),
            .carryin(n19799),
            .carryout(n19800),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__37044),
            .sr(N__36998));
    defparam acadc_skipcnt_i0_i12_LC_13_20_3.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i12_LC_13_20_3.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i12_LC_13_20_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i12_LC_13_20_3 (
            .in0(_gnd_net_),
            .in1(N__50621),
            .in2(_gnd_net_),
            .in3(N__36729),
            .lcout(acadc_skipcnt_12),
            .ltout(),
            .carryin(n19800),
            .carryout(n19801),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__37044),
            .sr(N__36998));
    defparam acadc_skipcnt_i0_i13_LC_13_20_4.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i13_LC_13_20_4.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i13_LC_13_20_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i13_LC_13_20_4 (
            .in0(_gnd_net_),
            .in1(N__37109),
            .in2(_gnd_net_),
            .in3(N__37095),
            .lcout(acadc_skipcnt_13),
            .ltout(),
            .carryin(n19801),
            .carryout(n19802),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__37044),
            .sr(N__36998));
    defparam acadc_skipcnt_i0_i14_LC_13_20_5.C_ON=1'b1;
    defparam acadc_skipcnt_i0_i14_LC_13_20_5.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i14_LC_13_20_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i14_LC_13_20_5 (
            .in0(_gnd_net_),
            .in1(N__37085),
            .in2(_gnd_net_),
            .in3(N__37071),
            .lcout(acadc_skipcnt_14),
            .ltout(),
            .carryin(n19802),
            .carryout(n19803),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__37044),
            .sr(N__36998));
    defparam acadc_skipcnt_i0_i15_LC_13_20_6.C_ON=1'b0;
    defparam acadc_skipcnt_i0_i15_LC_13_20_6.SEQ_MODE=4'b1000;
    defparam acadc_skipcnt_i0_i15_LC_13_20_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 acadc_skipcnt_i0_i15_LC_13_20_6 (
            .in0(_gnd_net_),
            .in1(N__37058),
            .in2(_gnd_net_),
            .in3(N__37068),
            .lcout(acadc_skipcnt_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVacadc_skipcnt_i0_i9C_net),
            .ce(N__37044),
            .sr(N__36998));
    defparam \comm_spi.imiso_83_12297_12298_reset_LC_14_2_0 .C_ON=1'b0;
    defparam \comm_spi.imiso_83_12297_12298_reset_LC_14_2_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.imiso_83_12297_12298_reset_LC_14_2_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.imiso_83_12297_12298_reset_LC_14_2_0  (
            .in0(N__39813),
            .in1(N__39797),
            .in2(_gnd_net_),
            .in3(N__44331),
            .lcout(\comm_spi.n14819 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.imiso_83_12297_12298_resetC_net ),
            .ce(),
            .sr(N__42888));
    defparam \comm_spi.data_tx_i7_12294_12295_reset_LC_14_3_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i7_12294_12295_reset_LC_14_3_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i7_12294_12295_reset_LC_14_3_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i7_12294_12295_reset_LC_14_3_0  (
            .in0(N__36972),
            .in1(N__36954),
            .in2(_gnd_net_),
            .in3(N__36933),
            .lcout(\comm_spi.n14816 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__58356),
            .ce(),
            .sr(N__42887));
    defparam \comm_spi.data_tx_i7_12294_12295_set_LC_14_4_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i7_12294_12295_set_LC_14_4_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i7_12294_12295_set_LC_14_4_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i7_12294_12295_set_LC_14_4_0  (
            .in0(N__36971),
            .in1(N__36950),
            .in2(_gnd_net_),
            .in3(N__36929),
            .lcout(\comm_spi.n14815 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__58257),
            .ce(),
            .sr(N__42836));
    defparam \ADC_VDC.genclk.t_clk_24_LC_14_5_1 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.t_clk_24_LC_14_5_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t_clk_24_LC_14_5_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ADC_VDC.genclk.t_clk_24_LC_14_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56586),
            .lcout(VDC_CLK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVADC_VDC.genclk.t_clk_24C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam i14_4_lut_LC_14_5_2.C_ON=1'b0;
    defparam i14_4_lut_LC_14_5_2.SEQ_MODE=4'b0000;
    defparam i14_4_lut_LC_14_5_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i14_4_lut_LC_14_5_2 (
            .in0(N__39758),
            .in1(N__39692),
            .in2(N__40038),
            .in3(N__39707),
            .lcout(n33),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i12289_3_lut_LC_14_5_4 .C_ON=1'b0;
    defparam \comm_spi.i12289_3_lut_LC_14_5_4 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i12289_3_lut_LC_14_5_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.i12289_3_lut_LC_14_5_4  (
            .in0(N__36904),
            .in1(N__36891),
            .in2(_gnd_net_),
            .in3(N__45025),
            .lcout(\comm_spi.imosi ),
            .ltout(\comm_spi.imosi_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_86_2_lut_LC_14_5_5 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_86_2_lut_LC_14_5_5 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_86_2_lut_LC_14_5_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \comm_spi.RESET_I_0_86_2_lut_LC_14_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__37173),
            .in3(N__58059),
            .lcout(\comm_spi.DOUT_7__N_786 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_88_2_lut_LC_14_5_7 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_88_2_lut_LC_14_5_7 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_88_2_lut_LC_14_5_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \comm_spi.RESET_I_0_88_2_lut_LC_14_5_7  (
            .in0(_gnd_net_),
            .in1(N__50891),
            .in2(_gnd_net_),
            .in3(N__58058),
            .lcout(\comm_spi.imosi_N_792 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i11_4_lut_LC_14_6_0.C_ON=1'b0;
    defparam i11_4_lut_LC_14_6_0.SEQ_MODE=4'b0000;
    defparam i11_4_lut_LC_14_6_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i11_4_lut_LC_14_6_0 (
            .in0(N__39722),
            .in1(N__39677),
            .in2(N__40113),
            .in3(N__40163),
            .lcout(n30_adj_1530),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i5_4_lut_LC_14_6_1.C_ON=1'b0;
    defparam i5_4_lut_LC_14_6_1.SEQ_MODE=4'b0000;
    defparam i5_4_lut_LC_14_6_1.LUT_INIT=16'b1000000000000000;
    LogicCell40 i5_4_lut_LC_14_6_1 (
            .in0(N__40358),
            .in1(N__40343),
            .in2(N__40131),
            .in3(N__40094),
            .lcout(),
            .ltout(n12_adj_1542_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6_4_lut_LC_14_6_2.C_ON=1'b0;
    defparam i6_4_lut_LC_14_6_2.SEQ_MODE=4'b0000;
    defparam i6_4_lut_LC_14_6_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 i6_4_lut_LC_14_6_2 (
            .in0(N__39980),
            .in1(N__40211),
            .in2(N__37149),
            .in3(N__40227),
            .lcout(),
            .ltout(n19986_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15_4_lut_LC_14_6_3.C_ON=1'b0;
    defparam i15_4_lut_LC_14_6_3.SEQ_MODE=4'b0000;
    defparam i15_4_lut_LC_14_6_3.LUT_INIT=16'b1111111111101111;
    LogicCell40 i15_4_lut_LC_14_6_3 (
            .in0(N__39944),
            .in1(N__40016),
            .in2(N__37146),
            .in3(N__37143),
            .lcout(),
            .ltout(n34_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18_4_lut_LC_14_6_4.C_ON=1'b0;
    defparam i18_4_lut_LC_14_6_4.SEQ_MODE=4'b0000;
    defparam i18_4_lut_LC_14_6_4.LUT_INIT=16'b1111111111111110;
    LogicCell40 i18_4_lut_LC_14_6_4 (
            .in0(N__37119),
            .in1(N__37137),
            .in2(N__37131),
            .in3(N__37128),
            .lcout(n49),
            .ltout(n49_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam wdtick_flag_289_LC_14_6_5.C_ON=1'b0;
    defparam wdtick_flag_289_LC_14_6_5.SEQ_MODE=4'b1010;
    defparam wdtick_flag_289_LC_14_6_5.LUT_INIT=16'b1111111100001111;
    LogicCell40 wdtick_flag_289_LC_14_6_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__37122),
            .in3(N__44815),
            .lcout(wdtick_flag),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50784),
            .ce(),
            .sr(N__42151));
    defparam i13_4_lut_LC_14_7_6.C_ON=1'b0;
    defparam i13_4_lut_LC_14_7_6.SEQ_MODE=4'b0000;
    defparam i13_4_lut_LC_14_7_6.LUT_INIT=16'b1111111111111110;
    LogicCell40 i13_4_lut_LC_14_7_6 (
            .in0(N__40178),
            .in1(N__40193),
            .in2(N__40149),
            .in3(N__40056),
            .lcout(n32),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.bit_cnt_3767__i3_LC_14_8_0 .C_ON=1'b0;
    defparam \comm_spi.bit_cnt_3767__i3_LC_14_8_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.bit_cnt_3767__i3_LC_14_8_0 .LUT_INIT=16'b0110110011001100;
    LogicCell40 \comm_spi.bit_cnt_3767__i3_LC_14_8_0  (
            .in0(N__37296),
            .in1(N__42791),
            .in2(N__37281),
            .in3(N__37314),
            .lcout(\comm_spi.bit_cnt_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.bit_cnt_3767__i3C_net ),
            .ce(),
            .sr(N__58165));
    defparam \comm_spi.bit_cnt_3767__i2_LC_14_8_1 .C_ON=1'b0;
    defparam \comm_spi.bit_cnt_3767__i2_LC_14_8_1 .SEQ_MODE=4'b1010;
    defparam \comm_spi.bit_cnt_3767__i2_LC_14_8_1 .LUT_INIT=16'b0111011110001000;
    LogicCell40 \comm_spi.bit_cnt_3767__i2_LC_14_8_1  (
            .in0(N__37313),
            .in1(N__37277),
            .in2(_gnd_net_),
            .in3(N__37295),
            .lcout(\comm_spi.bit_cnt_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.bit_cnt_3767__i3C_net ),
            .ce(),
            .sr(N__58165));
    defparam \comm_spi.bit_cnt_3767__i1_LC_14_8_2 .C_ON=1'b0;
    defparam \comm_spi.bit_cnt_3767__i1_LC_14_8_2 .SEQ_MODE=4'b1010;
    defparam \comm_spi.bit_cnt_3767__i1_LC_14_8_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \comm_spi.bit_cnt_3767__i1_LC_14_8_2  (
            .in0(N__37276),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37312),
            .lcout(\comm_spi.bit_cnt_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.bit_cnt_3767__i3C_net ),
            .ce(),
            .sr(N__58165));
    defparam \comm_spi.bit_cnt_3767__i0_LC_14_8_3 .C_ON=1'b0;
    defparam \comm_spi.bit_cnt_3767__i0_LC_14_8_3 .SEQ_MODE=4'b1010;
    defparam \comm_spi.bit_cnt_3767__i0_LC_14_8_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \comm_spi.bit_cnt_3767__i0_LC_14_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37275),
            .lcout(\comm_spi.bit_cnt_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.bit_cnt_3767__i3C_net ),
            .ce(),
            .sr(N__58165));
    defparam comm_cmd_1__bdd_4_lut_19721_LC_14_9_1.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19721_LC_14_9_1.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19721_LC_14_9_1.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_19721_LC_14_9_1 (
            .in0(N__37335),
            .in1(N__46462),
            .in2(N__37323),
            .in3(N__47697),
            .lcout(n22461),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i2_3_lut_LC_14_9_2 .C_ON=1'b0;
    defparam \comm_spi.i2_3_lut_LC_14_9_2 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i2_3_lut_LC_14_9_2 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \comm_spi.i2_3_lut_LC_14_9_2  (
            .in0(N__37311),
            .in1(N__37294),
            .in2(_gnd_net_),
            .in3(N__37274),
            .lcout(\comm_spi.n17254 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15452_2_lut_3_lut_LC_14_9_3.C_ON=1'b0;
    defparam i15452_2_lut_3_lut_LC_14_9_3.SEQ_MODE=4'b0000;
    defparam i15452_2_lut_3_lut_LC_14_9_3.LUT_INIT=16'b0000001000000010;
    LogicCell40 i15452_2_lut_3_lut_LC_14_9_3 (
            .in0(N__50414),
            .in1(N__54506),
            .in2(N__54853),
            .in3(_gnd_net_),
            .lcout(n14_adj_1579),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15462_2_lut_3_lut_LC_14_9_4.C_ON=1'b0;
    defparam i15462_2_lut_3_lut_LC_14_9_4.SEQ_MODE=4'b0000;
    defparam i15462_2_lut_3_lut_LC_14_9_4.LUT_INIT=16'b0001000100000000;
    LogicCell40 i15462_2_lut_3_lut_LC_14_9_4 (
            .in0(N__54504),
            .in1(N__54796),
            .in2(_gnd_net_),
            .in3(N__47786),
            .lcout(n14_adj_1572),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_4_lut_LC_14_9_5.C_ON=1'b0;
    defparam i1_2_lut_4_lut_LC_14_9_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_4_lut_LC_14_9_5.LUT_INIT=16'b1111111111111101;
    LogicCell40 i1_2_lut_4_lut_LC_14_9_5 (
            .in0(N__46461),
            .in1(N__47696),
            .in2(N__57262),
            .in3(N__53969),
            .lcout(n4_adj_1637),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15469_2_lut_3_lut_LC_14_9_6.C_ON=1'b0;
    defparam i15469_2_lut_3_lut_LC_14_9_6.SEQ_MODE=4'b0000;
    defparam i15469_2_lut_3_lut_LC_14_9_6.LUT_INIT=16'b0001000100000000;
    LogicCell40 i15469_2_lut_3_lut_LC_14_9_6 (
            .in0(N__54503),
            .in1(N__54795),
            .in2(_gnd_net_),
            .in3(N__42517),
            .lcout(n14_adj_1544),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15470_2_lut_3_lut_LC_14_9_7.C_ON=1'b0;
    defparam i15470_2_lut_3_lut_LC_14_9_7.SEQ_MODE=4'b0000;
    defparam i15470_2_lut_3_lut_LC_14_9_7.LUT_INIT=16'b0000001100000000;
    LogicCell40 i15470_2_lut_3_lut_LC_14_9_7 (
            .in0(_gnd_net_),
            .in1(N__54505),
            .in2(N__54852),
            .in3(N__53423),
            .lcout(n14_adj_1575),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19687_LC_14_10_0.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19687_LC_14_10_0.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19687_LC_14_10_0.LUT_INIT=16'b1111010110001000;
    LogicCell40 comm_cmd_1__bdd_4_lut_19687_LC_14_10_0 (
            .in0(N__47698),
            .in1(N__37431),
            .in2(N__37422),
            .in3(N__46463),
            .lcout(),
            .ltout(n22413_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22413_bdd_4_lut_LC_14_10_1.C_ON=1'b0;
    defparam n22413_bdd_4_lut_LC_14_10_1.SEQ_MODE=4'b0000;
    defparam n22413_bdd_4_lut_LC_14_10_1.LUT_INIT=16'b1111000011001010;
    LogicCell40 n22413_bdd_4_lut_LC_14_10_1 (
            .in0(N__37413),
            .in1(N__37407),
            .in2(N__37398),
            .in3(N__47699),
            .lcout(n22416),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19847_LC_14_10_3.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19847_LC_14_10_3.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19847_LC_14_10_3.LUT_INIT=16'b1101100010101010;
    LogicCell40 comm_cmd_1__bdd_4_lut_19847_LC_14_10_3 (
            .in0(N__46464),
            .in1(N__41754),
            .in2(N__37395),
            .in3(N__47700),
            .lcout(),
            .ltout(n22569_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22569_bdd_4_lut_LC_14_10_4.C_ON=1'b0;
    defparam n22569_bdd_4_lut_LC_14_10_4.SEQ_MODE=4'b0000;
    defparam n22569_bdd_4_lut_LC_14_10_4.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22569_bdd_4_lut_LC_14_10_4 (
            .in0(N__47701),
            .in1(N__37380),
            .in2(N__37365),
            .in3(N__37362),
            .lcout(),
            .ltout(n22572_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1565844_i1_3_lut_LC_14_10_5.C_ON=1'b0;
    defparam i1565844_i1_3_lut_LC_14_10_5.SEQ_MODE=4'b0000;
    defparam i1565844_i1_3_lut_LC_14_10_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 i1565844_i1_3_lut_LC_14_10_5 (
            .in0(_gnd_net_),
            .in1(N__37356),
            .in2(N__37350),
            .in3(N__47267),
            .lcout(),
            .ltout(n30_adj_1669_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_0__i5_LC_14_10_6.C_ON=1'b0;
    defparam comm_buf_0__i5_LC_14_10_6.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i5_LC_14_10_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 comm_buf_0__i5_LC_14_10_6 (
            .in0(_gnd_net_),
            .in1(N__53292),
            .in2(N__37347),
            .in3(N__54510),
            .lcout(comm_buf_0_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55959),
            .ce(N__43325),
            .sr(N__43249));
    defparam comm_buf_0__i7_LC_14_11_0.C_ON=1'b0;
    defparam comm_buf_0__i7_LC_14_11_0.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i7_LC_14_11_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 comm_buf_0__i7_LC_14_11_0 (
            .in0(N__48572),
            .in1(N__54509),
            .in2(_gnd_net_),
            .in3(N__37344),
            .lcout(comm_buf_0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55968),
            .ce(N__43338),
            .sr(N__43275));
    defparam comm_buf_0__i6_LC_14_11_1.C_ON=1'b0;
    defparam comm_buf_0__i6_LC_14_11_1.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i6_LC_14_11_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_0__i6_LC_14_11_1 (
            .in0(N__54507),
            .in1(N__53195),
            .in2(_gnd_net_),
            .in3(N__37629),
            .lcout(comm_buf_0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55968),
            .ce(N__43338),
            .sr(N__43275));
    defparam comm_buf_0__i3_LC_14_11_2.C_ON=1'b0;
    defparam comm_buf_0__i3_LC_14_11_2.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i3_LC_14_11_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 comm_buf_0__i3_LC_14_11_2 (
            .in0(N__49856),
            .in1(N__54508),
            .in2(_gnd_net_),
            .in3(N__37614),
            .lcout(comm_buf_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55968),
            .ce(N__43338),
            .sr(N__43275));
    defparam i22_4_lut_LC_14_12_0.C_ON=1'b0;
    defparam i22_4_lut_LC_14_12_0.SEQ_MODE=4'b0000;
    defparam i22_4_lut_LC_14_12_0.LUT_INIT=16'b1100111100001010;
    LogicCell40 i22_4_lut_LC_14_12_0 (
            .in0(N__52884),
            .in1(N__46038),
            .in2(N__54005),
            .in3(N__54737),
            .lcout(),
            .ltout(n8_adj_1689_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_i2_LC_14_12_1.C_ON=1'b0;
    defparam comm_state_i2_LC_14_12_1.SEQ_MODE=4'b1000;
    defparam comm_state_i2_LC_14_12_1.LUT_INIT=16'b0101000011001100;
    LogicCell40 comm_state_i2_LC_14_12_1 (
            .in0(N__52797),
            .in1(N__37545),
            .in2(N__37602),
            .in3(N__54494),
            .lcout(comm_state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55979),
            .ce(N__37596),
            .sr(N__55478));
    defparam i1_4_lut_adj_285_LC_14_12_2.C_ON=1'b0;
    defparam i1_4_lut_adj_285_LC_14_12_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_285_LC_14_12_2.LUT_INIT=16'b0010001100111000;
    LogicCell40 i1_4_lut_adj_285_LC_14_12_2 (
            .in0(N__52883),
            .in1(N__54685),
            .in2(N__54552),
            .in3(N__52799),
            .lcout(),
            .ltout(n26_adj_1595_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19442_2_lut_3_lut_LC_14_12_3.C_ON=1'b0;
    defparam i19442_2_lut_3_lut_LC_14_12_3.SEQ_MODE=4'b0000;
    defparam i19442_2_lut_3_lut_LC_14_12_3.LUT_INIT=16'b1100111111111111;
    LogicCell40 i19442_2_lut_3_lut_LC_14_12_3 (
            .in0(_gnd_net_),
            .in1(N__55183),
            .in2(N__37599),
            .in3(N__53982),
            .lcout(n18_adj_1615),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19360_4_lut_LC_14_12_4.C_ON=1'b0;
    defparam i19360_4_lut_LC_14_12_4.SEQ_MODE=4'b0000;
    defparam i19360_4_lut_LC_14_12_4.LUT_INIT=16'b0010000001110000;
    LogicCell40 i19360_4_lut_LC_14_12_4 (
            .in0(N__53981),
            .in1(N__52798),
            .in2(N__54810),
            .in3(N__37590),
            .lcout(n21714),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i22_4_lut_4_lut_LC_14_12_5.C_ON=1'b0;
    defparam i22_4_lut_4_lut_LC_14_12_5.SEQ_MODE=4'b0000;
    defparam i22_4_lut_4_lut_LC_14_12_5.LUT_INIT=16'b0100011001000100;
    LogicCell40 i22_4_lut_4_lut_LC_14_12_5 (
            .in0(N__54498),
            .in1(N__53980),
            .in2(N__52803),
            .in3(N__52882),
            .lcout(),
            .ltout(n7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_241_LC_14_12_6.C_ON=1'b0;
    defparam i1_4_lut_adj_241_LC_14_12_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_241_LC_14_12_6.LUT_INIT=16'b1011101000000000;
    LogicCell40 i1_4_lut_adj_241_LC_14_12_6 (
            .in0(N__55182),
            .in1(N__54684),
            .in2(N__37539),
            .in3(N__55553),
            .lcout(n12107),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_44_LC_14_12_7.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_44_LC_14_12_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_44_LC_14_12_7.LUT_INIT=16'b1111111111011101;
    LogicCell40 i1_2_lut_3_lut_adj_44_LC_14_12_7 (
            .in0(N__54683),
            .in1(N__55181),
            .in2(_gnd_net_),
            .in3(N__54490),
            .lcout(n21147),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_cntvec_i0_i0_LC_14_13_0.C_ON=1'b1;
    defparam data_cntvec_i0_i0_LC_14_13_0.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i0_LC_14_13_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i0_LC_14_13_0 (
            .in0(_gnd_net_),
            .in1(N__43840),
            .in2(N__37784),
            .in3(_gnd_net_),
            .lcout(data_cntvec_0),
            .ltout(),
            .carryin(bfn_14_13_0_),
            .carryout(n19774),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__37842),
            .sr(N__38151));
    defparam data_cntvec_i0_i1_LC_14_13_1.C_ON=1'b1;
    defparam data_cntvec_i0_i1_LC_14_13_1.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i1_LC_14_13_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i1_LC_14_13_1 (
            .in0(_gnd_net_),
            .in1(N__44195),
            .in2(_gnd_net_),
            .in3(N__37728),
            .lcout(data_cntvec_1),
            .ltout(),
            .carryin(n19774),
            .carryout(n19775),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__37842),
            .sr(N__38151));
    defparam data_cntvec_i0_i2_LC_14_13_2.C_ON=1'b1;
    defparam data_cntvec_i0_i2_LC_14_13_2.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i2_LC_14_13_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i2_LC_14_13_2 (
            .in0(_gnd_net_),
            .in1(N__37721),
            .in2(_gnd_net_),
            .in3(N__37701),
            .lcout(data_cntvec_2),
            .ltout(),
            .carryin(n19775),
            .carryout(n19776),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__37842),
            .sr(N__38151));
    defparam data_cntvec_i0_i3_LC_14_13_3.C_ON=1'b1;
    defparam data_cntvec_i0_i3_LC_14_13_3.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i3_LC_14_13_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i3_LC_14_13_3 (
            .in0(_gnd_net_),
            .in1(N__41219),
            .in2(_gnd_net_),
            .in3(N__37698),
            .lcout(data_cntvec_3),
            .ltout(),
            .carryin(n19776),
            .carryout(n19777),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__37842),
            .sr(N__38151));
    defparam data_cntvec_i0_i4_LC_14_13_4.C_ON=1'b1;
    defparam data_cntvec_i0_i4_LC_14_13_4.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i4_LC_14_13_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i4_LC_14_13_4 (
            .in0(_gnd_net_),
            .in1(N__37691),
            .in2(_gnd_net_),
            .in3(N__37671),
            .lcout(data_cntvec_4),
            .ltout(),
            .carryin(n19777),
            .carryout(n19778),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__37842),
            .sr(N__38151));
    defparam data_cntvec_i0_i5_LC_14_13_5.C_ON=1'b1;
    defparam data_cntvec_i0_i5_LC_14_13_5.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i5_LC_14_13_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i5_LC_14_13_5 (
            .in0(_gnd_net_),
            .in1(N__37660),
            .in2(_gnd_net_),
            .in3(N__37638),
            .lcout(data_cntvec_5),
            .ltout(),
            .carryin(n19778),
            .carryout(n19779),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__37842),
            .sr(N__38151));
    defparam data_cntvec_i0_i6_LC_14_13_6.C_ON=1'b1;
    defparam data_cntvec_i0_i6_LC_14_13_6.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i6_LC_14_13_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i6_LC_14_13_6 (
            .in0(_gnd_net_),
            .in1(N__43436),
            .in2(_gnd_net_),
            .in3(N__37635),
            .lcout(data_cntvec_6),
            .ltout(),
            .carryin(n19779),
            .carryout(n19780),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__37842),
            .sr(N__38151));
    defparam data_cntvec_i0_i7_LC_14_13_7.C_ON=1'b1;
    defparam data_cntvec_i0_i7_LC_14_13_7.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i7_LC_14_13_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i7_LC_14_13_7 (
            .in0(_gnd_net_),
            .in1(N__46519),
            .in2(_gnd_net_),
            .in3(N__37632),
            .lcout(data_cntvec_7),
            .ltout(),
            .carryin(n19780),
            .carryout(n19781),
            .clk(INVdata_cntvec_i0_i0C_net),
            .ce(N__37842),
            .sr(N__38151));
    defparam data_cntvec_i0_i8_LC_14_14_0.C_ON=1'b1;
    defparam data_cntvec_i0_i8_LC_14_14_0.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i8_LC_14_14_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i8_LC_14_14_0 (
            .in0(_gnd_net_),
            .in1(N__40901),
            .in2(_gnd_net_),
            .in3(N__37971),
            .lcout(data_cntvec_8),
            .ltout(),
            .carryin(bfn_14_14_0_),
            .carryout(n19782),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__37844),
            .sr(N__38150));
    defparam data_cntvec_i0_i9_LC_14_14_1.C_ON=1'b1;
    defparam data_cntvec_i0_i9_LC_14_14_1.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i9_LC_14_14_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i9_LC_14_14_1 (
            .in0(_gnd_net_),
            .in1(N__43078),
            .in2(_gnd_net_),
            .in3(N__37968),
            .lcout(data_cntvec_9),
            .ltout(),
            .carryin(n19782),
            .carryout(n19783),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__37844),
            .sr(N__38150));
    defparam data_cntvec_i0_i10_LC_14_14_2.C_ON=1'b1;
    defparam data_cntvec_i0_i10_LC_14_14_2.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i10_LC_14_14_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i10_LC_14_14_2 (
            .in0(_gnd_net_),
            .in1(N__40678),
            .in2(_gnd_net_),
            .in3(N__37965),
            .lcout(data_cntvec_10),
            .ltout(),
            .carryin(n19783),
            .carryout(n19784),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__37844),
            .sr(N__38150));
    defparam data_cntvec_i0_i11_LC_14_14_3.C_ON=1'b1;
    defparam data_cntvec_i0_i11_LC_14_14_3.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i11_LC_14_14_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i11_LC_14_14_3 (
            .in0(_gnd_net_),
            .in1(N__37954),
            .in2(_gnd_net_),
            .in3(N__37932),
            .lcout(data_cntvec_11),
            .ltout(),
            .carryin(n19784),
            .carryout(n19785),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__37844),
            .sr(N__38150));
    defparam data_cntvec_i0_i12_LC_14_14_4.C_ON=1'b1;
    defparam data_cntvec_i0_i12_LC_14_14_4.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i12_LC_14_14_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i12_LC_14_14_4 (
            .in0(_gnd_net_),
            .in1(N__37925),
            .in2(_gnd_net_),
            .in3(N__37911),
            .lcout(data_cntvec_12),
            .ltout(),
            .carryin(n19785),
            .carryout(n19786),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__37844),
            .sr(N__38150));
    defparam data_cntvec_i0_i13_LC_14_14_5.C_ON=1'b1;
    defparam data_cntvec_i0_i13_LC_14_14_5.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i13_LC_14_14_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i13_LC_14_14_5 (
            .in0(_gnd_net_),
            .in1(N__37904),
            .in2(_gnd_net_),
            .in3(N__37890),
            .lcout(data_cntvec_13),
            .ltout(),
            .carryin(n19786),
            .carryout(n19787),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__37844),
            .sr(N__38150));
    defparam data_cntvec_i0_i14_LC_14_14_6.C_ON=1'b1;
    defparam data_cntvec_i0_i14_LC_14_14_6.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i14_LC_14_14_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i14_LC_14_14_6 (
            .in0(_gnd_net_),
            .in1(N__37883),
            .in2(_gnd_net_),
            .in3(N__37869),
            .lcout(data_cntvec_14),
            .ltout(),
            .carryin(n19787),
            .carryout(n19788),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__37844),
            .sr(N__38150));
    defparam data_cntvec_i0_i15_LC_14_14_7.C_ON=1'b0;
    defparam data_cntvec_i0_i15_LC_14_14_7.SEQ_MODE=4'b1000;
    defparam data_cntvec_i0_i15_LC_14_14_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 data_cntvec_i0_i15_LC_14_14_7 (
            .in0(_gnd_net_),
            .in1(N__37859),
            .in2(_gnd_net_),
            .in3(N__37866),
            .lcout(data_cntvec_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVdata_cntvec_i0_i8C_net),
            .ce(N__37844),
            .sr(N__38150));
    defparam add_125_2_lut_LC_14_15_0.C_ON=1'b1;
    defparam add_125_2_lut_LC_14_15_0.SEQ_MODE=4'b0000;
    defparam add_125_2_lut_LC_14_15_0.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_125_2_lut_LC_14_15_0 (
            .in0(N__41141),
            .in1(N__41140),
            .in2(N__38927),
            .in3(N__38106),
            .lcout(n7_adj_1539),
            .ltout(),
            .carryin(bfn_14_15_0_),
            .carryout(n19804),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_125_3_lut_LC_14_15_1.C_ON=1'b1;
    defparam add_125_3_lut_LC_14_15_1.SEQ_MODE=4'b0000;
    defparam add_125_3_lut_LC_14_15_1.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_125_3_lut_LC_14_15_1 (
            .in0(N__39357),
            .in1(N__39356),
            .in2(N__38931),
            .in3(N__38103),
            .lcout(n7_adj_1569),
            .ltout(),
            .carryin(n19804),
            .carryout(n19805),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_125_4_lut_LC_14_15_2.C_ON=1'b1;
    defparam add_125_4_lut_LC_14_15_2.SEQ_MODE=4'b0000;
    defparam add_125_4_lut_LC_14_15_2.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_125_4_lut_LC_14_15_2 (
            .in0(N__39222),
            .in1(N__39221),
            .in2(N__38928),
            .in3(N__38100),
            .lcout(n7_adj_1567),
            .ltout(),
            .carryin(n19805),
            .carryout(n19806),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_125_5_lut_LC_14_15_3.C_ON=1'b1;
    defparam add_125_5_lut_LC_14_15_3.SEQ_MODE=4'b0000;
    defparam add_125_5_lut_LC_14_15_3.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_125_5_lut_LC_14_15_3 (
            .in0(N__38097),
            .in1(N__38095),
            .in2(N__38932),
            .in3(N__38067),
            .lcout(n7_adj_1565),
            .ltout(),
            .carryin(n19806),
            .carryout(n19807),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_125_6_lut_LC_14_15_4.C_ON=1'b1;
    defparam add_125_6_lut_LC_14_15_4.SEQ_MODE=4'b0000;
    defparam add_125_6_lut_LC_14_15_4.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_125_6_lut_LC_14_15_4 (
            .in0(N__38184),
            .in1(N__38183),
            .in2(N__38929),
            .in3(N__38064),
            .lcout(n7_adj_1563),
            .ltout(),
            .carryin(n19807),
            .carryout(n19808),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_125_7_lut_LC_14_15_5.C_ON=1'b1;
    defparam add_125_7_lut_LC_14_15_5.SEQ_MODE=4'b0000;
    defparam add_125_7_lut_LC_14_15_5.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_125_7_lut_LC_14_15_5 (
            .in0(N__39057),
            .in1(N__39056),
            .in2(N__38933),
            .in3(N__38061),
            .lcout(n17703),
            .ltout(),
            .carryin(n19808),
            .carryout(n19809),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_125_8_lut_LC_14_15_6.C_ON=1'b1;
    defparam add_125_8_lut_LC_14_15_6.SEQ_MODE=4'b0000;
    defparam add_125_8_lut_LC_14_15_6.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_125_8_lut_LC_14_15_6 (
            .in0(N__38058),
            .in1(N__38057),
            .in2(N__38930),
            .in3(N__38013),
            .lcout(n7_adj_1561),
            .ltout(),
            .carryin(n19809),
            .carryout(n19810),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_125_9_lut_LC_14_15_7.C_ON=1'b1;
    defparam add_125_9_lut_LC_14_15_7.SEQ_MODE=4'b0000;
    defparam add_125_9_lut_LC_14_15_7.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_125_9_lut_LC_14_15_7 (
            .in0(N__38010),
            .in1(N__38009),
            .in2(N__38934),
            .in3(N__37977),
            .lcout(n7_adj_1559),
            .ltout(),
            .carryin(n19810),
            .carryout(n19811),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_125_10_lut_LC_14_16_0.C_ON=1'b1;
    defparam add_125_10_lut_LC_14_16_0.SEQ_MODE=4'b0000;
    defparam add_125_10_lut_LC_14_16_0.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_125_10_lut_LC_14_16_0 (
            .in0(N__39177),
            .in1(N__39176),
            .in2(N__38944),
            .in3(N__37974),
            .lcout(n7_adj_1557),
            .ltout(),
            .carryin(bfn_14_16_0_),
            .carryout(n19812),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam add_125_11_lut_LC_14_16_1.C_ON=1'b0;
    defparam add_125_11_lut_LC_14_16_1.SEQ_MODE=4'b0000;
    defparam add_125_11_lut_LC_14_16_1.LUT_INIT=16'b1010001110101100;
    LogicCell40 add_125_11_lut_LC_14_16_1 (
            .in0(N__38962),
            .in1(N__38963),
            .in2(N__38945),
            .in3(N__38859),
            .lcout(n7_adj_1555),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_1_i30_3_lut_LC_14_16_2.C_ON=1'b0;
    defparam mux_130_Mux_1_i30_3_lut_LC_14_16_2.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_1_i30_3_lut_LC_14_16_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_130_Mux_1_i30_3_lut_LC_14_16_2 (
            .in0(N__38856),
            .in1(N__38835),
            .in2(_gnd_net_),
            .in3(N__47271),
            .lcout(n30_adj_1618),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam trig_dds1_305_LC_14_16_3.C_ON=1'b0;
    defparam trig_dds1_305_LC_14_16_3.SEQ_MODE=4'b1000;
    defparam trig_dds1_305_LC_14_16_3.LUT_INIT=16'b0110000001100100;
    LogicCell40 trig_dds1_305_LC_14_16_3 (
            .in0(N__49061),
            .in1(N__55459),
            .in2(N__38810),
            .in3(N__46938),
            .lcout(trig_dds1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56037),
            .ce(),
            .sr(_gnd_net_));
    defparam i15204_3_lut_LC_14_16_4.C_ON=1'b0;
    defparam i15204_3_lut_LC_14_16_4.SEQ_MODE=4'b0000;
    defparam i15204_3_lut_LC_14_16_4.LUT_INIT=16'b1100110010101010;
    LogicCell40 i15204_3_lut_LC_14_16_4 (
            .in0(N__50422),
            .in1(N__39055),
            .in2(_gnd_net_),
            .in3(N__41102),
            .lcout(n17705),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i6_LC_14_16_5.C_ON=1'b0;
    defparam buf_dds0_i6_LC_14_16_5.SEQ_MODE=4'b1000;
    defparam buf_dds0_i6_LC_14_16_5.LUT_INIT=16'b0101000011001100;
    LogicCell40 buf_dds0_i6_LC_14_16_5 (
            .in0(N__49059),
            .in1(N__41456),
            .in2(N__49495),
            .in3(N__41614),
            .lcout(buf_dds0_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56037),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i7_LC_14_16_7.C_ON=1'b0;
    defparam buf_dds0_i7_LC_14_16_7.SEQ_MODE=4'b1000;
    defparam buf_dds0_i7_LC_14_16_7.LUT_INIT=16'b0101000011001100;
    LogicCell40 buf_dds0_i7_LC_14_16_7 (
            .in0(N__49060),
            .in1(N__38790),
            .in2(N__44082),
            .in3(N__41615),
            .lcout(buf_dds0_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56037),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_IAC.ADC_DATA_i10_LC_14_17_1 .C_ON=1'b0;
    defparam \ADC_IAC.ADC_DATA_i10_LC_14_17_1 .SEQ_MODE=4'b1000;
    defparam \ADC_IAC.ADC_DATA_i10_LC_14_17_1 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \ADC_IAC.ADC_DATA_i10_LC_14_17_1  (
            .in0(N__38773),
            .in1(N__38570),
            .in2(N__38236),
            .in3(N__38263),
            .lcout(buf_adcdata_iac_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56053),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i4_LC_14_17_2.C_ON=1'b0;
    defparam data_index_i4_LC_14_17_2.SEQ_MODE=4'b1000;
    defparam data_index_i4_LC_14_17_2.LUT_INIT=16'b0011101100001000;
    LogicCell40 data_index_i4_LC_14_17_2 (
            .in0(N__38205),
            .in1(N__55294),
            .in2(N__49258),
            .in3(N__38199),
            .lcout(data_index_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56053),
            .ce(),
            .sr(_gnd_net_));
    defparam trig_dds0_304_LC_14_17_3.C_ON=1'b0;
    defparam trig_dds0_304_LC_14_17_3.SEQ_MODE=4'b1000;
    defparam trig_dds0_304_LC_14_17_3.LUT_INIT=16'b0010001011110000;
    LogicCell40 trig_dds0_304_LC_14_17_3 (
            .in0(N__55292),
            .in1(N__49127),
            .in2(N__43944),
            .in3(N__38163),
            .lcout(trig_dds0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56053),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19663_LC_14_17_4.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19663_LC_14_17_4.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19663_LC_14_17_4.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_cmd_0__bdd_4_lut_19663_LC_14_17_4 (
            .in0(N__39460),
            .in1(N__57212),
            .in2(N__39150),
            .in3(N__46467),
            .lcout(),
            .ltout(n22389_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22389_bdd_4_lut_LC_14_17_5.C_ON=1'b0;
    defparam n22389_bdd_4_lut_LC_14_17_5.SEQ_MODE=4'b0000;
    defparam n22389_bdd_4_lut_LC_14_17_5.LUT_INIT=16'b1110010111100000;
    LogicCell40 n22389_bdd_4_lut_LC_14_17_5 (
            .in0(N__46468),
            .in1(N__39111),
            .in2(N__39084),
            .in3(N__39077),
            .lcout(n22392),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i9_LC_14_17_6.C_ON=1'b0;
    defparam data_index_i9_LC_14_17_6.SEQ_MODE=4'b1000;
    defparam data_index_i9_LC_14_17_6.LUT_INIT=16'b0101000011001100;
    LogicCell40 data_index_i9_LC_14_17_6 (
            .in0(N__49126),
            .in1(N__41900),
            .in2(N__41922),
            .in3(N__55295),
            .lcout(data_index_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56053),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i5_LC_14_17_7.C_ON=1'b0;
    defparam data_index_i5_LC_14_17_7.SEQ_MODE=4'b1000;
    defparam data_index_i5_LC_14_17_7.LUT_INIT=16'b0101000011011000;
    LogicCell40 data_index_i5_LC_14_17_7 (
            .in0(N__55293),
            .in1(N__41439),
            .in2(N__41424),
            .in3(N__49131),
            .lcout(data_index_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56053),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.SCLK_27_LC_14_18_0 .C_ON=1'b0;
    defparam \SIG_DDS.SCLK_27_LC_14_18_0 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.SCLK_27_LC_14_18_0 .LUT_INIT=16'b0111001000110001;
    LogicCell40 \SIG_DDS.SCLK_27_LC_14_18_0  (
            .in0(N__44409),
            .in1(N__44670),
            .in2(N__39026),
            .in3(N__44752),
            .lcout(DDS_SCK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56066),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.MOSI_31_LC_14_18_1 .C_ON=1'b0;
    defparam \SIG_DDS.MOSI_31_LC_14_18_1 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.MOSI_31_LC_14_18_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \SIG_DDS.MOSI_31_LC_14_18_1  (
            .in0(N__39009),
            .in1(N__44408),
            .in2(_gnd_net_),
            .in3(N__38975),
            .lcout(DDS_MOSI),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56066),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i1_LC_14_18_3.C_ON=1'b0;
    defparam data_index_i1_LC_14_18_3.SEQ_MODE=4'b1000;
    defparam data_index_i1_LC_14_18_3.LUT_INIT=16'b0100111101000000;
    LogicCell40 data_index_i1_LC_14_18_3 (
            .in0(N__49124),
            .in1(N__39336),
            .in2(N__55479),
            .in3(N__39327),
            .lcout(data_index_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56066),
            .ce(),
            .sr(_gnd_net_));
    defparam i6294_3_lut_LC_14_18_4.C_ON=1'b0;
    defparam i6294_3_lut_LC_14_18_4.SEQ_MODE=4'b0000;
    defparam i6294_3_lut_LC_14_18_4.LUT_INIT=16'b1100110010101010;
    LogicCell40 i6294_3_lut_LC_14_18_4 (
            .in0(N__53437),
            .in1(N__38964),
            .in2(_gnd_net_),
            .in3(N__41119),
            .lcout(n8_adj_1556),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6364_3_lut_LC_14_18_5.C_ON=1'b0;
    defparam i6364_3_lut_LC_14_18_5.SEQ_MODE=4'b0000;
    defparam i6364_3_lut_LC_14_18_5.LUT_INIT=16'b1110111001000100;
    LogicCell40 i6364_3_lut_LC_14_18_5 (
            .in0(N__41120),
            .in1(N__45465),
            .in2(_gnd_net_),
            .in3(N__39214),
            .lcout(n8_adj_1568),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_cfgRTD_i1_LC_14_18_6.C_ON=1'b0;
    defparam buf_cfgRTD_i1_LC_14_18_6.SEQ_MODE=4'b1000;
    defparam buf_cfgRTD_i1_LC_14_18_6.LUT_INIT=16'b0011000010111000;
    LogicCell40 buf_cfgRTD_i1_LC_14_18_6 (
            .in0(N__53438),
            .in1(N__39662),
            .in2(N__39563),
            .in3(N__49125),
            .lcout(buf_cfgRTD_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56066),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_device_acadc_i1_LC_14_18_7.C_ON=1'b0;
    defparam buf_device_acadc_i1_LC_14_18_7.SEQ_MODE=4'b1000;
    defparam buf_device_acadc_i1_LC_14_18_7.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_device_acadc_i1_LC_14_18_7 (
            .in0(N__49123),
            .in1(N__39543),
            .in2(N__45635),
            .in3(N__39461),
            .lcout(IAC_OSR0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56066),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_354_Mux_8_i15_4_lut_LC_14_19_0.C_ON=1'b0;
    defparam comm_state_3__I_0_354_Mux_8_i15_4_lut_LC_14_19_0.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_354_Mux_8_i15_4_lut_LC_14_19_0.LUT_INIT=16'b0011101100001000;
    LogicCell40 comm_state_3__I_0_354_Mux_8_i15_4_lut_LC_14_19_0 (
            .in0(N__39197),
            .in1(N__55472),
            .in2(N__49242),
            .in3(N__39188),
            .lcout(data_index_9_N_212_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6304_3_lut_LC_14_19_2.C_ON=1'b0;
    defparam i6304_3_lut_LC_14_19_2.SEQ_MODE=4'b0000;
    defparam i6304_3_lut_LC_14_19_2.LUT_INIT=16'b1110111001000100;
    LogicCell40 i6304_3_lut_LC_14_19_2 (
            .in0(N__41121),
            .in1(N__45616),
            .in2(_gnd_net_),
            .in3(N__39169),
            .lcout(n8_adj_1558),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i6374_3_lut_LC_14_19_3.C_ON=1'b0;
    defparam i6374_3_lut_LC_14_19_3.SEQ_MODE=4'b0000;
    defparam i6374_3_lut_LC_14_19_3.LUT_INIT=16'b1100110010101010;
    LogicCell40 i6374_3_lut_LC_14_19_3 (
            .in0(N__53499),
            .in1(N__39355),
            .in2(_gnd_net_),
            .in3(N__41122),
            .lcout(n8_adj_1570),
            .ltout(n8_adj_1570_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_354_Mux_1_i15_4_lut_LC_14_19_4.C_ON=1'b0;
    defparam comm_state_3__I_0_354_Mux_1_i15_4_lut_LC_14_19_4.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_354_Mux_1_i15_4_lut_LC_14_19_4.LUT_INIT=16'b0111001101000000;
    LogicCell40 comm_state_3__I_0_354_Mux_1_i15_4_lut_LC_14_19_4 (
            .in0(N__49103),
            .in1(N__55471),
            .in2(N__39330),
            .in3(N__39326),
            .lcout(data_index_9_N_212_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i2_LC_14_19_5.C_ON=1'b0;
    defparam data_index_i2_LC_14_19_5.SEQ_MODE=4'b1000;
    defparam data_index_i2_LC_14_19_5.LUT_INIT=16'b0111010100100000;
    LogicCell40 data_index_i2_LC_14_19_5 (
            .in0(N__55473),
            .in1(N__49108),
            .in2(N__39930),
            .in3(N__39915),
            .lcout(data_index_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56079),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i8_LC_14_19_6.C_ON=1'b0;
    defparam data_index_i8_LC_14_19_6.SEQ_MODE=4'b1000;
    defparam data_index_i8_LC_14_19_6.LUT_INIT=16'b0011101100001000;
    LogicCell40 data_index_i8_LC_14_19_6 (
            .in0(N__39198),
            .in1(N__55474),
            .in2(N__49243),
            .in3(N__39189),
            .lcout(data_index_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56079),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_354_Mux_2_i15_4_lut_LC_14_19_7.C_ON=1'b0;
    defparam comm_state_3__I_0_354_Mux_2_i15_4_lut_LC_14_19_7.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_354_Mux_2_i15_4_lut_LC_14_19_7.LUT_INIT=16'b0111010100100000;
    LogicCell40 comm_state_3__I_0_354_Mux_2_i15_4_lut_LC_14_19_7 (
            .in0(N__55470),
            .in1(N__49104),
            .in2(N__39929),
            .in3(N__39914),
            .lcout(data_index_9_N_212_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.imiso_83_12297_12298_set_LC_15_3_6 .C_ON=1'b0;
    defparam \comm_spi.imiso_83_12297_12298_set_LC_15_3_6 .SEQ_MODE=4'b1011;
    defparam \comm_spi.imiso_83_12297_12298_set_LC_15_3_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.imiso_83_12297_12298_set_LC_15_3_6  (
            .in0(N__39812),
            .in1(N__39798),
            .in2(_gnd_net_),
            .in3(N__44323),
            .lcout(\comm_spi.n14818 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.imiso_83_12297_12298_setC_net ),
            .ce(),
            .sr(N__42837));
    defparam \comm_spi.RESET_I_0_87_2_lut_LC_15_4_5 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_87_2_lut_LC_15_4_5 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_87_2_lut_LC_15_4_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \comm_spi.RESET_I_0_87_2_lut_LC_15_4_5  (
            .in0(N__39786),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58158),
            .lcout(\comm_spi.DOUT_7__N_787 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam wdtick_cnt_3763_3764__i1_LC_15_5_0.C_ON=1'b1;
    defparam wdtick_cnt_3763_3764__i1_LC_15_5_0.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3763_3764__i1_LC_15_5_0.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3763_3764__i1_LC_15_5_0 (
            .in0(N__40321),
            .in1(N__39759),
            .in2(_gnd_net_),
            .in3(N__39747),
            .lcout(wdtick_cnt_0),
            .ltout(),
            .carryin(bfn_15_5_0_),
            .carryout(n19932),
            .clk(N__50785),
            .ce(N__42635),
            .sr(N__42153));
    defparam wdtick_cnt_3763_3764__i2_LC_15_5_1.C_ON=1'b1;
    defparam wdtick_cnt_3763_3764__i2_LC_15_5_1.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3763_3764__i2_LC_15_5_1.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3763_3764__i2_LC_15_5_1 (
            .in0(N__40313),
            .in1(N__39740),
            .in2(_gnd_net_),
            .in3(N__39726),
            .lcout(wdtick_cnt_1),
            .ltout(),
            .carryin(n19932),
            .carryout(n19933),
            .clk(N__50785),
            .ce(N__42635),
            .sr(N__42153));
    defparam wdtick_cnt_3763_3764__i3_LC_15_5_2.C_ON=1'b1;
    defparam wdtick_cnt_3763_3764__i3_LC_15_5_2.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3763_3764__i3_LC_15_5_2.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3763_3764__i3_LC_15_5_2 (
            .in0(N__40322),
            .in1(N__39723),
            .in2(_gnd_net_),
            .in3(N__39711),
            .lcout(wdtick_cnt_2),
            .ltout(),
            .carryin(n19933),
            .carryout(n19934),
            .clk(N__50785),
            .ce(N__42635),
            .sr(N__42153));
    defparam wdtick_cnt_3763_3764__i4_LC_15_5_3.C_ON=1'b1;
    defparam wdtick_cnt_3763_3764__i4_LC_15_5_3.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3763_3764__i4_LC_15_5_3.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3763_3764__i4_LC_15_5_3 (
            .in0(N__40314),
            .in1(N__39708),
            .in2(_gnd_net_),
            .in3(N__39696),
            .lcout(wdtick_cnt_3),
            .ltout(),
            .carryin(n19934),
            .carryout(n19935),
            .clk(N__50785),
            .ce(N__42635),
            .sr(N__42153));
    defparam wdtick_cnt_3763_3764__i5_LC_15_5_4.C_ON=1'b1;
    defparam wdtick_cnt_3763_3764__i5_LC_15_5_4.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3763_3764__i5_LC_15_5_4.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3763_3764__i5_LC_15_5_4 (
            .in0(N__40323),
            .in1(N__39693),
            .in2(_gnd_net_),
            .in3(N__39681),
            .lcout(wdtick_cnt_4),
            .ltout(),
            .carryin(n19935),
            .carryout(n19936),
            .clk(N__50785),
            .ce(N__42635),
            .sr(N__42153));
    defparam wdtick_cnt_3763_3764__i6_LC_15_5_5.C_ON=1'b1;
    defparam wdtick_cnt_3763_3764__i6_LC_15_5_5.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3763_3764__i6_LC_15_5_5.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3763_3764__i6_LC_15_5_5 (
            .in0(N__40315),
            .in1(N__39678),
            .in2(_gnd_net_),
            .in3(N__39666),
            .lcout(wdtick_cnt_5),
            .ltout(),
            .carryin(n19936),
            .carryout(n19937),
            .clk(N__50785),
            .ce(N__42635),
            .sr(N__42153));
    defparam wdtick_cnt_3763_3764__i7_LC_15_5_6.C_ON=1'b1;
    defparam wdtick_cnt_3763_3764__i7_LC_15_5_6.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3763_3764__i7_LC_15_5_6.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3763_3764__i7_LC_15_5_6 (
            .in0(N__40324),
            .in1(N__40073),
            .in2(_gnd_net_),
            .in3(N__40059),
            .lcout(wdtick_cnt_6),
            .ltout(),
            .carryin(n19937),
            .carryout(n19938),
            .clk(N__50785),
            .ce(N__42635),
            .sr(N__42153));
    defparam wdtick_cnt_3763_3764__i8_LC_15_5_7.C_ON=1'b1;
    defparam wdtick_cnt_3763_3764__i8_LC_15_5_7.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3763_3764__i8_LC_15_5_7.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3763_3764__i8_LC_15_5_7 (
            .in0(N__40316),
            .in1(N__40055),
            .in2(_gnd_net_),
            .in3(N__40041),
            .lcout(wdtick_cnt_7),
            .ltout(),
            .carryin(n19938),
            .carryout(n19939),
            .clk(N__50785),
            .ce(N__42635),
            .sr(N__42153));
    defparam wdtick_cnt_3763_3764__i9_LC_15_6_0.C_ON=1'b1;
    defparam wdtick_cnt_3763_3764__i9_LC_15_6_0.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3763_3764__i9_LC_15_6_0.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3763_3764__i9_LC_15_6_0 (
            .in0(N__40308),
            .in1(N__40034),
            .in2(_gnd_net_),
            .in3(N__40020),
            .lcout(wdtick_cnt_8),
            .ltout(),
            .carryin(bfn_15_6_0_),
            .carryout(n19940),
            .clk(N__50787),
            .ce(N__42631),
            .sr(N__42147));
    defparam wdtick_cnt_3763_3764__i10_LC_15_6_1.C_ON=1'b1;
    defparam wdtick_cnt_3763_3764__i10_LC_15_6_1.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3763_3764__i10_LC_15_6_1.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3763_3764__i10_LC_15_6_1 (
            .in0(N__40326),
            .in1(N__40017),
            .in2(_gnd_net_),
            .in3(N__40005),
            .lcout(wdtick_cnt_9),
            .ltout(),
            .carryin(n19940),
            .carryout(n19941),
            .clk(N__50787),
            .ce(N__42631),
            .sr(N__42147));
    defparam wdtick_cnt_3763_3764__i11_LC_15_6_2.C_ON=1'b1;
    defparam wdtick_cnt_3763_3764__i11_LC_15_6_2.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3763_3764__i11_LC_15_6_2.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3763_3764__i11_LC_15_6_2 (
            .in0(N__40305),
            .in1(N__39998),
            .in2(_gnd_net_),
            .in3(N__39984),
            .lcout(wdtick_cnt_10),
            .ltout(),
            .carryin(n19941),
            .carryout(n19942),
            .clk(N__50787),
            .ce(N__42631),
            .sr(N__42147));
    defparam wdtick_cnt_3763_3764__i12_LC_15_6_3.C_ON=1'b1;
    defparam wdtick_cnt_3763_3764__i12_LC_15_6_3.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3763_3764__i12_LC_15_6_3.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3763_3764__i12_LC_15_6_3 (
            .in0(N__40327),
            .in1(N__39981),
            .in2(_gnd_net_),
            .in3(N__39969),
            .lcout(wdtick_cnt_11),
            .ltout(),
            .carryin(n19942),
            .carryout(n19943),
            .clk(N__50787),
            .ce(N__42631),
            .sr(N__42147));
    defparam wdtick_cnt_3763_3764__i13_LC_15_6_4.C_ON=1'b1;
    defparam wdtick_cnt_3763_3764__i13_LC_15_6_4.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3763_3764__i13_LC_15_6_4.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3763_3764__i13_LC_15_6_4 (
            .in0(N__40306),
            .in1(N__39962),
            .in2(_gnd_net_),
            .in3(N__39948),
            .lcout(wdtick_cnt_12),
            .ltout(),
            .carryin(n19943),
            .carryout(n19944),
            .clk(N__50787),
            .ce(N__42631),
            .sr(N__42147));
    defparam wdtick_cnt_3763_3764__i14_LC_15_6_5.C_ON=1'b1;
    defparam wdtick_cnt_3763_3764__i14_LC_15_6_5.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3763_3764__i14_LC_15_6_5.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3763_3764__i14_LC_15_6_5 (
            .in0(N__40328),
            .in1(N__39945),
            .in2(_gnd_net_),
            .in3(N__39933),
            .lcout(wdtick_cnt_13),
            .ltout(),
            .carryin(n19944),
            .carryout(n19945),
            .clk(N__50787),
            .ce(N__42631),
            .sr(N__42147));
    defparam wdtick_cnt_3763_3764__i15_LC_15_6_6.C_ON=1'b1;
    defparam wdtick_cnt_3763_3764__i15_LC_15_6_6.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3763_3764__i15_LC_15_6_6.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3763_3764__i15_LC_15_6_6 (
            .in0(N__40307),
            .in1(N__40212),
            .in2(_gnd_net_),
            .in3(N__40197),
            .lcout(wdtick_cnt_14),
            .ltout(),
            .carryin(n19945),
            .carryout(n19946),
            .clk(N__50787),
            .ce(N__42631),
            .sr(N__42147));
    defparam wdtick_cnt_3763_3764__i16_LC_15_6_7.C_ON=1'b1;
    defparam wdtick_cnt_3763_3764__i16_LC_15_6_7.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3763_3764__i16_LC_15_6_7.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3763_3764__i16_LC_15_6_7 (
            .in0(N__40329),
            .in1(N__40194),
            .in2(_gnd_net_),
            .in3(N__40182),
            .lcout(wdtick_cnt_15),
            .ltout(),
            .carryin(n19946),
            .carryout(n19947),
            .clk(N__50787),
            .ce(N__42631),
            .sr(N__42147));
    defparam wdtick_cnt_3763_3764__i17_LC_15_7_0.C_ON=1'b1;
    defparam wdtick_cnt_3763_3764__i17_LC_15_7_0.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3763_3764__i17_LC_15_7_0.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3763_3764__i17_LC_15_7_0 (
            .in0(N__40317),
            .in1(N__40179),
            .in2(_gnd_net_),
            .in3(N__40167),
            .lcout(wdtick_cnt_16),
            .ltout(),
            .carryin(bfn_15_7_0_),
            .carryout(n19948),
            .clk(N__50789),
            .ce(N__42630),
            .sr(N__42143));
    defparam wdtick_cnt_3763_3764__i18_LC_15_7_1.C_ON=1'b1;
    defparam wdtick_cnt_3763_3764__i18_LC_15_7_1.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3763_3764__i18_LC_15_7_1.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3763_3764__i18_LC_15_7_1 (
            .in0(N__40309),
            .in1(N__40164),
            .in2(_gnd_net_),
            .in3(N__40152),
            .lcout(wdtick_cnt_17),
            .ltout(),
            .carryin(n19948),
            .carryout(n19949),
            .clk(N__50789),
            .ce(N__42630),
            .sr(N__42143));
    defparam wdtick_cnt_3763_3764__i19_LC_15_7_2.C_ON=1'b1;
    defparam wdtick_cnt_3763_3764__i19_LC_15_7_2.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3763_3764__i19_LC_15_7_2.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3763_3764__i19_LC_15_7_2 (
            .in0(N__40318),
            .in1(N__40148),
            .in2(_gnd_net_),
            .in3(N__40134),
            .lcout(wdtick_cnt_18),
            .ltout(),
            .carryin(n19949),
            .carryout(n19950),
            .clk(N__50789),
            .ce(N__42630),
            .sr(N__42143));
    defparam wdtick_cnt_3763_3764__i20_LC_15_7_3.C_ON=1'b1;
    defparam wdtick_cnt_3763_3764__i20_LC_15_7_3.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3763_3764__i20_LC_15_7_3.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3763_3764__i20_LC_15_7_3 (
            .in0(N__40310),
            .in1(N__40130),
            .in2(_gnd_net_),
            .in3(N__40116),
            .lcout(wdtick_cnt_19),
            .ltout(),
            .carryin(n19950),
            .carryout(n19951),
            .clk(N__50789),
            .ce(N__42630),
            .sr(N__42143));
    defparam wdtick_cnt_3763_3764__i21_LC_15_7_4.C_ON=1'b1;
    defparam wdtick_cnt_3763_3764__i21_LC_15_7_4.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3763_3764__i21_LC_15_7_4.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3763_3764__i21_LC_15_7_4 (
            .in0(N__40319),
            .in1(N__40112),
            .in2(_gnd_net_),
            .in3(N__40098),
            .lcout(wdtick_cnt_20),
            .ltout(),
            .carryin(n19951),
            .carryout(n19952),
            .clk(N__50789),
            .ce(N__42630),
            .sr(N__42143));
    defparam wdtick_cnt_3763_3764__i22_LC_15_7_5.C_ON=1'b1;
    defparam wdtick_cnt_3763_3764__i22_LC_15_7_5.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3763_3764__i22_LC_15_7_5.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3763_3764__i22_LC_15_7_5 (
            .in0(N__40311),
            .in1(N__40095),
            .in2(_gnd_net_),
            .in3(N__40083),
            .lcout(wdtick_cnt_21),
            .ltout(),
            .carryin(n19952),
            .carryout(n19953),
            .clk(N__50789),
            .ce(N__42630),
            .sr(N__42143));
    defparam wdtick_cnt_3763_3764__i23_LC_15_7_6.C_ON=1'b1;
    defparam wdtick_cnt_3763_3764__i23_LC_15_7_6.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3763_3764__i23_LC_15_7_6.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3763_3764__i23_LC_15_7_6 (
            .in0(N__40320),
            .in1(N__40359),
            .in2(_gnd_net_),
            .in3(N__40347),
            .lcout(wdtick_cnt_22),
            .ltout(),
            .carryin(n19953),
            .carryout(n19954),
            .clk(N__50789),
            .ce(N__42630),
            .sr(N__42143));
    defparam wdtick_cnt_3763_3764__i24_LC_15_7_7.C_ON=1'b1;
    defparam wdtick_cnt_3763_3764__i24_LC_15_7_7.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3763_3764__i24_LC_15_7_7.LUT_INIT=16'b1000001000101000;
    LogicCell40 wdtick_cnt_3763_3764__i24_LC_15_7_7 (
            .in0(N__40312),
            .in1(N__40344),
            .in2(_gnd_net_),
            .in3(N__40332),
            .lcout(wdtick_cnt_23),
            .ltout(),
            .carryin(n19954),
            .carryout(n19955),
            .clk(N__50789),
            .ce(N__42630),
            .sr(N__42143));
    defparam wdtick_cnt_3763_3764__i25_LC_15_8_0.C_ON=1'b0;
    defparam wdtick_cnt_3763_3764__i25_LC_15_8_0.SEQ_MODE=4'b1010;
    defparam wdtick_cnt_3763_3764__i25_LC_15_8_0.LUT_INIT=16'b1000010001001000;
    LogicCell40 wdtick_cnt_3763_3764__i25_LC_15_8_0 (
            .in0(N__40226),
            .in1(N__40325),
            .in2(_gnd_net_),
            .in3(N__40230),
            .lcout(wdtick_cnt_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50790),
            .ce(N__42636),
            .sr(N__42152));
    defparam \comm_spi.data_rx_i7_LC_15_9_0 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i7_LC_15_9_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i7_LC_15_9_0 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \comm_spi.data_rx_i7_LC_15_9_0  (
            .in0(N__53160),
            .in1(N__42781),
            .in2(_gnd_net_),
            .in3(N__42746),
            .lcout(comm_rx_buf_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__58402),
            .ce(),
            .sr(N__58145));
    defparam \comm_spi.data_rx_i6_LC_15_9_1 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i6_LC_15_9_1 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i6_LC_15_9_1 .LUT_INIT=16'b1100100011001000;
    LogicCell40 \comm_spi.data_rx_i6_LC_15_9_1  (
            .in0(N__42745),
            .in1(N__53291),
            .in2(N__42797),
            .in3(_gnd_net_),
            .lcout(comm_rx_buf_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__58402),
            .ce(),
            .sr(N__58145));
    defparam \comm_spi.data_rx_i5_LC_15_9_2 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i5_LC_15_9_2 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i5_LC_15_9_2 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \comm_spi.data_rx_i5_LC_15_9_2  (
            .in0(N__53584),
            .in1(N__42780),
            .in2(_gnd_net_),
            .in3(N__42744),
            .lcout(comm_rx_buf_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__58402),
            .ce(),
            .sr(N__58145));
    defparam \comm_spi.data_rx_i4_LC_15_9_3 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i4_LC_15_9_3 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i4_LC_15_9_3 .LUT_INIT=16'b1100100011001000;
    LogicCell40 \comm_spi.data_rx_i4_LC_15_9_3  (
            .in0(N__42743),
            .in1(N__49810),
            .in2(N__42796),
            .in3(_gnd_net_),
            .lcout(comm_rx_buf_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__58402),
            .ce(),
            .sr(N__58145));
    defparam \comm_spi.data_rx_i3_LC_15_9_4 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i3_LC_15_9_4 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i3_LC_15_9_4 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \comm_spi.data_rx_i3_LC_15_9_4  (
            .in0(N__50094),
            .in1(N__42779),
            .in2(_gnd_net_),
            .in3(N__42742),
            .lcout(comm_rx_buf_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__58402),
            .ce(),
            .sr(N__58145));
    defparam \comm_spi.data_rx_i2_LC_15_9_5 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i2_LC_15_9_5 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i2_LC_15_9_5 .LUT_INIT=16'b1111101000000000;
    LogicCell40 \comm_spi.data_rx_i2_LC_15_9_5  (
            .in0(N__42741),
            .in1(_gnd_net_),
            .in2(N__42795),
            .in3(N__49659),
            .lcout(comm_rx_buf_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__58402),
            .ce(),
            .sr(N__58145));
    defparam \comm_spi.data_rx_i1_LC_15_9_6 .C_ON=1'b0;
    defparam \comm_spi.data_rx_i1_LC_15_9_6 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_rx_i1_LC_15_9_6 .LUT_INIT=16'b1010101010001000;
    LogicCell40 \comm_spi.data_rx_i1_LC_15_9_6  (
            .in0(N__48677),
            .in1(N__42778),
            .in2(_gnd_net_),
            .in3(N__42740),
            .lcout(comm_rx_buf_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__58402),
            .ce(),
            .sr(N__58145));
    defparam clk_RTD_287_LC_15_10_0.C_ON=1'b0;
    defparam clk_RTD_287_LC_15_10_0.SEQ_MODE=4'b1000;
    defparam clk_RTD_287_LC_15_10_0.LUT_INIT=16'b0110011010101010;
    LogicCell40 clk_RTD_287_LC_15_10_0 (
            .in0(N__40473),
            .in1(N__45000),
            .in2(_gnd_net_),
            .in3(N__44976),
            .lcout(clk_RTD),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50792),
            .ce(),
            .sr(_gnd_net_));
    defparam i19121_2_lut_LC_15_10_1.C_ON=1'b0;
    defparam i19121_2_lut_LC_15_10_1.SEQ_MODE=4'b0000;
    defparam i19121_2_lut_LC_15_10_1.LUT_INIT=16'b0101010100000000;
    LogicCell40 i19121_2_lut_LC_15_10_1 (
            .in0(N__53965),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48188),
            .lcout(n21588),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19054_2_lut_3_lut_LC_15_10_2.C_ON=1'b0;
    defparam i19054_2_lut_3_lut_LC_15_10_2.SEQ_MODE=4'b0000;
    defparam i19054_2_lut_3_lut_LC_15_10_2.LUT_INIT=16'b1110111011111111;
    LogicCell40 i19054_2_lut_3_lut_LC_15_10_2 (
            .in0(N__46036),
            .in1(N__52762),
            .in2(_gnd_net_),
            .in3(N__53964),
            .lcout(n21586),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12442_2_lut_LC_15_10_3.C_ON=1'b0;
    defparam i12442_2_lut_LC_15_10_3.SEQ_MODE=4'b0000;
    defparam i12442_2_lut_LC_15_10_3.LUT_INIT=16'b1010101000000000;
    LogicCell40 i12442_2_lut_LC_15_10_3 (
            .in0(N__55068),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43305),
            .lcout(n14958),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15473_2_lut_3_lut_LC_15_10_4.C_ON=1'b0;
    defparam i15473_2_lut_3_lut_LC_15_10_4.SEQ_MODE=4'b0000;
    defparam i15473_2_lut_3_lut_LC_15_10_4.LUT_INIT=16'b0000000001000100;
    LogicCell40 i15473_2_lut_3_lut_LC_15_10_4 (
            .in0(N__54754),
            .in1(N__45620),
            .in2(_gnd_net_),
            .in3(N__54367),
            .lcout(n14_adj_1550),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18549_4_lut_LC_15_10_5.C_ON=1'b0;
    defparam i18549_4_lut_LC_15_10_5.SEQ_MODE=4'b0000;
    defparam i18549_4_lut_LC_15_10_5.LUT_INIT=16'b0010111000100010;
    LogicCell40 i18549_4_lut_LC_15_10_5 (
            .in0(N__42471),
            .in1(N__52382),
            .in2(N__53070),
            .in3(N__43559),
            .lcout(n21276),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_250_LC_15_10_6.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_250_LC_15_10_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_250_LC_15_10_6.LUT_INIT=16'b1110111011111111;
    LogicCell40 i1_2_lut_3_lut_adj_250_LC_15_10_6 (
            .in0(N__54753),
            .in1(N__54366),
            .in2(_gnd_net_),
            .in3(N__55067),
            .lcout(n12433),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22461_bdd_4_lut_LC_15_11_0.C_ON=1'b0;
    defparam n22461_bdd_4_lut_LC_15_11_0.SEQ_MODE=4'b0000;
    defparam n22461_bdd_4_lut_LC_15_11_0.LUT_INIT=16'b1100110010111000;
    LogicCell40 n22461_bdd_4_lut_LC_15_11_0 (
            .in0(N__40422),
            .in1(N__40413),
            .in2(N__40401),
            .in3(N__47530),
            .lcout(n22464),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19172_2_lut_LC_15_11_1.C_ON=1'b0;
    defparam i19172_2_lut_LC_15_11_1.SEQ_MODE=4'b0000;
    defparam i19172_2_lut_LC_15_11_1.LUT_INIT=16'b1100110000000000;
    LogicCell40 i19172_2_lut_LC_15_11_1 (
            .in0(_gnd_net_),
            .in1(N__40383),
            .in2(_gnd_net_),
            .in3(N__57179),
            .lcout(),
            .ltout(n21556_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19770_LC_15_11_2.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19770_LC_15_11_2.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19770_LC_15_11_2.LUT_INIT=16'b1011100011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_19770_LC_15_11_2 (
            .in0(N__42168),
            .in1(N__46471),
            .in2(N__40779),
            .in3(N__47529),
            .lcout(n22521),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22521_bdd_4_lut_LC_15_11_4.C_ON=1'b0;
    defparam n22521_bdd_4_lut_LC_15_11_4.SEQ_MODE=4'b0000;
    defparam n22521_bdd_4_lut_LC_15_11_4.LUT_INIT=16'b1100110010111000;
    LogicCell40 n22521_bdd_4_lut_LC_15_11_4 (
            .in0(N__40776),
            .in1(N__40764),
            .in2(N__41478),
            .in3(N__47531),
            .lcout(),
            .ltout(n22524_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1565241_i1_3_lut_LC_15_11_5.C_ON=1'b0;
    defparam i1565241_i1_3_lut_LC_15_11_5.SEQ_MODE=4'b0000;
    defparam i1565241_i1_3_lut_LC_15_11_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 i1565241_i1_3_lut_LC_15_11_5 (
            .in0(_gnd_net_),
            .in1(N__40758),
            .in2(N__40752),
            .in3(N__47163),
            .lcout(),
            .ltout(n30_adj_1676_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_0__i4_LC_15_11_6.C_ON=1'b0;
    defparam comm_buf_0__i4_LC_15_11_6.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i4_LC_15_11_6.LUT_INIT=16'b1010101011110000;
    LogicCell40 comm_buf_0__i4_LC_15_11_6 (
            .in0(N__53600),
            .in1(_gnd_net_),
            .in2(N__40749),
            .in3(N__54401),
            .lcout(comm_buf_0_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55980),
            .ce(N__43326),
            .sr(N__43250));
    defparam n22485_bdd_4_lut_LC_15_12_1.C_ON=1'b0;
    defparam n22485_bdd_4_lut_LC_15_12_1.SEQ_MODE=4'b0000;
    defparam n22485_bdd_4_lut_LC_15_12_1.LUT_INIT=16'b1110111000110000;
    LogicCell40 n22485_bdd_4_lut_LC_15_12_1 (
            .in0(N__40746),
            .in1(N__47691),
            .in2(N__40731),
            .in3(N__40716),
            .lcout(n22488),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_2_i26_3_lut_LC_15_12_2.C_ON=1'b0;
    defparam mux_128_Mux_2_i26_3_lut_LC_15_12_2.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_2_i26_3_lut_LC_15_12_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_128_Mux_2_i26_3_lut_LC_15_12_2 (
            .in0(N__40704),
            .in1(N__57114),
            .in2(_gnd_net_),
            .in3(N__40682),
            .lcout(),
            .ltout(n26_adj_1687_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19716_LC_15_12_3.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19716_LC_15_12_3.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19716_LC_15_12_3.LUT_INIT=16'b1011101111000000;
    LogicCell40 comm_cmd_1__bdd_4_lut_19716_LC_15_12_3 (
            .in0(N__52590),
            .in1(N__47692),
            .in2(N__40656),
            .in3(N__46485),
            .lcout(),
            .ltout(n22455_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22455_bdd_4_lut_LC_15_12_4.C_ON=1'b0;
    defparam n22455_bdd_4_lut_LC_15_12_4.SEQ_MODE=4'b0000;
    defparam n22455_bdd_4_lut_LC_15_12_4.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22455_bdd_4_lut_LC_15_12_4 (
            .in0(N__47693),
            .in1(N__45699),
            .in2(N__40653),
            .in3(N__40650),
            .lcout(),
            .ltout(n22458_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1564035_i1_3_lut_LC_15_12_5.C_ON=1'b0;
    defparam i1564035_i1_3_lut_LC_15_12_5.SEQ_MODE=4'b0000;
    defparam i1564035_i1_3_lut_LC_15_12_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 i1564035_i1_3_lut_LC_15_12_5 (
            .in0(_gnd_net_),
            .in1(N__40632),
            .in2(N__40626),
            .in3(N__47268),
            .lcout(),
            .ltout(n30_adj_1688_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_0__i2_LC_15_12_6.C_ON=1'b0;
    defparam comm_buf_0__i2_LC_15_12_6.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i2_LC_15_12_6.LUT_INIT=16'b1010101011110000;
    LogicCell40 comm_buf_0__i2_LC_15_12_6 (
            .in0(N__50108),
            .in1(_gnd_net_),
            .in2(N__40932),
            .in3(N__54402),
            .lcout(comm_buf_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55993),
            .ce(N__43336),
            .sr(N__43264));
    defparam mux_128_Mux_0_i26_3_lut_LC_15_13_2.C_ON=1'b0;
    defparam mux_128_Mux_0_i26_3_lut_LC_15_13_2.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_0_i26_3_lut_LC_15_13_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_128_Mux_0_i26_3_lut_LC_15_13_2 (
            .in0(N__40929),
            .in1(N__57109),
            .in2(_gnd_net_),
            .in3(N__40897),
            .lcout(),
            .ltout(n26_adj_1533_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18519_4_lut_LC_15_13_3.C_ON=1'b0;
    defparam i18519_4_lut_LC_15_13_3.SEQ_MODE=4'b0000;
    defparam i18519_4_lut_LC_15_13_3.LUT_INIT=16'b0100010011110000;
    LogicCell40 i18519_4_lut_LC_15_13_3 (
            .in0(N__57110),
            .in1(N__40881),
            .in2(N__40866),
            .in3(N__46409),
            .lcout(),
            .ltout(n21246_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_2__bdd_4_lut_19828_LC_15_13_4.C_ON=1'b0;
    defparam comm_cmd_2__bdd_4_lut_19828_LC_15_13_4.SEQ_MODE=4'b0000;
    defparam comm_cmd_2__bdd_4_lut_19828_LC_15_13_4.LUT_INIT=16'b1111010110001000;
    LogicCell40 comm_cmd_2__bdd_4_lut_19828_LC_15_13_4 (
            .in0(N__47250),
            .in1(N__40863),
            .in2(N__40854),
            .in3(N__47710),
            .lcout(),
            .ltout(n22581_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22581_bdd_4_lut_LC_15_13_5.C_ON=1'b0;
    defparam n22581_bdd_4_lut_LC_15_13_5.SEQ_MODE=4'b0000;
    defparam n22581_bdd_4_lut_LC_15_13_5.LUT_INIT=16'b1111000011001010;
    LogicCell40 n22581_bdd_4_lut_LC_15_13_5 (
            .in0(N__40851),
            .in1(N__40839),
            .in2(N__40824),
            .in3(N__47251),
            .lcout(),
            .ltout(n22584_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_0__i0_LC_15_13_6.C_ON=1'b0;
    defparam comm_buf_0__i0_LC_15_13_6.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i0_LC_15_13_6.LUT_INIT=16'b1111101001010000;
    LogicCell40 comm_buf_0__i0_LC_15_13_6 (
            .in0(N__54400),
            .in1(_gnd_net_),
            .in2(N__40821),
            .in3(N__48676),
            .lcout(comm_buf_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56007),
            .ce(N__43337),
            .sr(N__43263));
    defparam i19282_4_lut_4_lut_LC_15_13_7.C_ON=1'b0;
    defparam i19282_4_lut_4_lut_LC_15_13_7.SEQ_MODE=4'b0000;
    defparam i19282_4_lut_4_lut_LC_15_13_7.LUT_INIT=16'b1011111011110011;
    LogicCell40 i19282_4_lut_4_lut_LC_15_13_7 (
            .in0(N__47709),
            .in1(N__46408),
            .in2(N__57217),
            .in3(N__47249),
            .lcout(n21479),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i3_LC_15_14_0.C_ON=1'b0;
    defparam comm_buf_1__i3_LC_15_14_0.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i3_LC_15_14_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_1__i3_LC_15_14_0 (
            .in0(N__54556),
            .in1(N__49860),
            .in2(_gnd_net_),
            .in3(N__41250),
            .lcout(comm_buf_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56023),
            .ce(N__45199),
            .sr(N__44009));
    defparam comm_cmd_1__bdd_4_lut_19862_LC_15_14_1.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19862_LC_15_14_1.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19862_LC_15_14_1.LUT_INIT=16'b1101110110100000;
    LogicCell40 comm_cmd_1__bdd_4_lut_19862_LC_15_14_1 (
            .in0(N__47663),
            .in1(N__40818),
            .in2(N__40794),
            .in3(N__46479),
            .lcout(),
            .ltout(n22623_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22623_bdd_4_lut_LC_15_14_2.C_ON=1'b0;
    defparam n22623_bdd_4_lut_LC_15_14_2.SEQ_MODE=4'b0000;
    defparam n22623_bdd_4_lut_LC_15_14_2.LUT_INIT=16'b1111000010101100;
    LogicCell40 n22623_bdd_4_lut_LC_15_14_2 (
            .in0(N__41304),
            .in1(N__41265),
            .in2(N__41256),
            .in3(N__47664),
            .lcout(),
            .ltout(n22626_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1568859_i1_3_lut_LC_15_14_3.C_ON=1'b0;
    defparam i1568859_i1_3_lut_LC_15_14_3.SEQ_MODE=4'b0000;
    defparam i1568859_i1_3_lut_LC_15_14_3.LUT_INIT=16'b1111110000110000;
    LogicCell40 i1568859_i1_3_lut_LC_15_14_3 (
            .in0(_gnd_net_),
            .in1(N__47255),
            .in2(N__41253),
            .in3(N__41148),
            .lcout(n30_adj_1643),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_3_i26_3_lut_LC_15_14_4.C_ON=1'b0;
    defparam mux_129_Mux_3_i26_3_lut_LC_15_14_4.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_3_i26_3_lut_LC_15_14_4.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_129_Mux_3_i26_3_lut_LC_15_14_4 (
            .in0(N__41244),
            .in1(N__57128),
            .in2(_gnd_net_),
            .in3(N__41215),
            .lcout(),
            .ltout(n26_adj_1642_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19692_LC_15_14_5.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19692_LC_15_14_5.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19692_LC_15_14_5.LUT_INIT=16'b1101110110100000;
    LogicCell40 comm_cmd_1__bdd_4_lut_19692_LC_15_14_5 (
            .in0(N__47661),
            .in1(N__56601),
            .in2(N__41199),
            .in3(N__46478),
            .lcout(),
            .ltout(n22425_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22425_bdd_4_lut_LC_15_14_6.C_ON=1'b0;
    defparam n22425_bdd_4_lut_LC_15_14_6.SEQ_MODE=4'b0000;
    defparam n22425_bdd_4_lut_LC_15_14_6.LUT_INIT=16'b1110001111100000;
    LogicCell40 n22425_bdd_4_lut_LC_15_14_6 (
            .in0(N__41196),
            .in1(N__47662),
            .in2(N__41172),
            .in3(N__41169),
            .lcout(n22428),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam data_index_i0_LC_15_15_0.C_ON=1'b0;
    defparam data_index_i0_LC_15_15_0.SEQ_MODE=4'b1000;
    defparam data_index_i0_LC_15_15_0.LUT_INIT=16'b0000101011001100;
    LogicCell40 data_index_i0_LC_15_15_0 (
            .in0(N__41052),
            .in1(N__41046),
            .in2(N__49331),
            .in3(N__55288),
            .lcout(data_index_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56038),
            .ce(),
            .sr(_gnd_net_));
    defparam i4379_3_lut_LC_15_15_1.C_ON=1'b0;
    defparam i4379_3_lut_LC_15_15_1.SEQ_MODE=4'b0000;
    defparam i4379_3_lut_LC_15_15_1.LUT_INIT=16'b1100110010101010;
    LogicCell40 i4379_3_lut_LC_15_15_1 (
            .in0(N__45669),
            .in1(N__41142),
            .in2(_gnd_net_),
            .in3(N__41123),
            .lcout(n8_adj_1540),
            .ltout(n8_adj_1540_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_354_Mux_0_i15_4_lut_LC_15_15_2.C_ON=1'b0;
    defparam comm_state_3__I_0_354_Mux_0_i15_4_lut_LC_15_15_2.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_354_Mux_0_i15_4_lut_LC_15_15_2.LUT_INIT=16'b0101000011001100;
    LogicCell40 comm_state_3__I_0_354_Mux_0_i15_4_lut_LC_15_15_2 (
            .in0(N__49234),
            .in1(N__41045),
            .in2(N__41037),
            .in3(N__55287),
            .lcout(data_index_9_N_212_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i4_LC_15_15_3.C_ON=1'b0;
    defparam buf_control_i4_LC_15_15_3.SEQ_MODE=4'b1000;
    defparam buf_control_i4_LC_15_15_3.LUT_INIT=16'b0010111100100000;
    LogicCell40 buf_control_i4_LC_15_15_3 (
            .in0(N__47774),
            .in1(N__49235),
            .in2(N__42009),
            .in3(N__41497),
            .lcout(VDC_RNG0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56038),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i0_LC_15_15_4.C_ON=1'b0;
    defparam buf_dds1_i0_LC_15_15_4.SEQ_MODE=4'b1000;
    defparam buf_dds1_i0_LC_15_15_4.LUT_INIT=16'b1100101000000000;
    LogicCell40 buf_dds1_i0_LC_15_15_4 (
            .in0(N__41723),
            .in1(N__45670),
            .in2(N__46917),
            .in3(N__46745),
            .lcout(buf_dds1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56038),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_0_i16_3_lut_LC_15_15_5.C_ON=1'b0;
    defparam mux_129_Mux_0_i16_3_lut_LC_15_15_5.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_0_i16_3_lut_LC_15_15_5.LUT_INIT=16'b1110111001000100;
    LogicCell40 mux_129_Mux_0_i16_3_lut_LC_15_15_5 (
            .in0(N__57113),
            .in1(N__41530),
            .in2(_gnd_net_),
            .in3(N__41722),
            .lcout(),
            .ltout(n16_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18530_3_lut_LC_15_15_6.C_ON=1'b0;
    defparam i18530_3_lut_LC_15_15_6.SEQ_MODE=4'b0000;
    defparam i18530_3_lut_LC_15_15_6.LUT_INIT=16'b1111110000110000;
    LogicCell40 i18530_3_lut_LC_15_15_6 (
            .in0(_gnd_net_),
            .in1(N__46376),
            .in2(N__41709),
            .in3(N__41705),
            .lcout(n21257),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds0_i0_LC_15_15_7.C_ON=1'b0;
    defparam buf_dds0_i0_LC_15_15_7.SEQ_MODE=4'b1000;
    defparam buf_dds0_i0_LC_15_15_7.LUT_INIT=16'b1010101011001100;
    LogicCell40 buf_dds0_i0_LC_15_15_7 (
            .in0(N__43194),
            .in1(N__41531),
            .in2(_gnd_net_),
            .in3(N__41637),
            .lcout(buf_dds0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56038),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_4_i23_3_lut_LC_15_16_0.C_ON=1'b0;
    defparam mux_128_Mux_4_i23_3_lut_LC_15_16_0.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_4_i23_3_lut_LC_15_16_0.LUT_INIT=16'b1111110000110000;
    LogicCell40 mux_128_Mux_4_i23_3_lut_LC_15_16_0 (
            .in0(_gnd_net_),
            .in1(N__57111),
            .in2(N__41501),
            .in3(N__50649),
            .lcout(n23_adj_1675),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_6_i16_3_lut_LC_15_16_1.C_ON=1'b0;
    defparam mux_129_Mux_6_i16_3_lut_LC_15_16_1.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_6_i16_3_lut_LC_15_16_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_129_Mux_6_i16_3_lut_LC_15_16_1 (
            .in0(N__46958),
            .in1(N__41455),
            .in2(_gnd_net_),
            .in3(N__57112),
            .lcout(n16_adj_1624),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4272_2_lut_LC_15_16_4.C_ON=1'b0;
    defparam i4272_2_lut_LC_15_16_4.SEQ_MODE=4'b0000;
    defparam i4272_2_lut_LC_15_16_4.LUT_INIT=16'b1111111111001100;
    LogicCell40 i4272_2_lut_LC_15_16_4 (
            .in0(_gnd_net_),
            .in1(N__54827),
            .in2(_gnd_net_),
            .in3(N__54380),
            .lcout(n9342),
            .ltout(n9342_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15206_4_lut_LC_15_16_5.C_ON=1'b0;
    defparam i15206_4_lut_LC_15_16_5.SEQ_MODE=4'b0000;
    defparam i15206_4_lut_LC_15_16_5.LUT_INIT=16'b0101110100001000;
    LogicCell40 i15206_4_lut_LC_15_16_5 (
            .in0(N__55286),
            .in1(N__41438),
            .in2(N__41427),
            .in3(N__41417),
            .lcout(data_index_9_N_212_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18635_3_lut_LC_15_16_6.C_ON=1'b0;
    defparam i18635_3_lut_LC_15_16_6.SEQ_MODE=4'b0000;
    defparam i18635_3_lut_LC_15_16_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 i18635_3_lut_LC_15_16_6 (
            .in0(N__46477),
            .in1(N__42050),
            .in2(_gnd_net_),
            .in3(N__42021),
            .lcout(n21362),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_control_i6_LC_15_16_7.C_ON=1'b0;
    defparam buf_control_i6_LC_15_16_7.SEQ_MODE=4'b1000;
    defparam buf_control_i6_LC_15_16_7.LUT_INIT=16'b0111001101000000;
    LogicCell40 buf_control_i6_LC_15_16_7 (
            .in0(N__49062),
            .in1(N__42008),
            .in2(N__49585),
            .in3(N__50710),
            .lcout(buf_control_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56054),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.CS_28_LC_15_18_0 .C_ON=1'b0;
    defparam \SIG_DDS.CS_28_LC_15_18_0 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.CS_28_LC_15_18_0 .LUT_INIT=16'b0001000110111011;
    LogicCell40 \SIG_DDS.CS_28_LC_15_18_0  (
            .in0(N__44669),
            .in1(N__44726),
            .in2(_gnd_net_),
            .in3(N__44388),
            .lcout(DDS_CS),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56080),
            .ce(N__41934),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_354_Mux_9_i15_4_lut_LC_15_19_0.C_ON=1'b0;
    defparam comm_state_3__I_0_354_Mux_9_i15_4_lut_LC_15_19_0.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_354_Mux_9_i15_4_lut_LC_15_19_0.LUT_INIT=16'b0010111100100000;
    LogicCell40 comm_state_3__I_0_354_Mux_9_i15_4_lut_LC_15_19_0 (
            .in0(N__41915),
            .in1(N__49112),
            .in2(N__55463),
            .in3(N__41904),
            .lcout(data_index_9_N_212_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.MISO_48_12291_12292_reset_LC_16_2_0 .C_ON=1'b0;
    defparam \comm_spi.MISO_48_12291_12292_reset_LC_16_2_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.MISO_48_12291_12292_reset_LC_16_2_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.MISO_48_12291_12292_reset_LC_16_2_0  (
            .in0(N__41799),
            .in1(N__41783),
            .in2(_gnd_net_),
            .in3(N__44313),
            .lcout(\comm_spi.n14813 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.MISO_48_12291_12292_resetC_net ),
            .ce(),
            .sr(N__42880));
    defparam \comm_spi.MISO_48_12291_12292_set_LC_16_3_0 .C_ON=1'b0;
    defparam \comm_spi.MISO_48_12291_12292_set_LC_16_3_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.MISO_48_12291_12292_set_LC_16_3_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.MISO_48_12291_12292_set_LC_16_3_0  (
            .in0(N__41798),
            .in1(N__41787),
            .in2(_gnd_net_),
            .in3(N__44312),
            .lcout(\comm_spi.n14812 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.MISO_48_12291_12292_setC_net ),
            .ce(),
            .sr(N__42829));
    defparam i19344_2_lut_LC_16_4_1.C_ON=1'b0;
    defparam i19344_2_lut_LC_16_4_1.SEQ_MODE=4'b0000;
    defparam i19344_2_lut_LC_16_4_1.LUT_INIT=16'b0000000011001100;
    LogicCell40 i19344_2_lut_LC_16_4_1 (
            .in0(_gnd_net_),
            .in1(N__41769),
            .in2(_gnd_net_),
            .in3(N__57272),
            .lcout(n21672),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i19397_2_lut_LC_16_4_2 .C_ON=1'b0;
    defparam \ADC_VDC.i19397_2_lut_LC_16_4_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i19397_2_lut_LC_16_4_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \ADC_VDC.i19397_2_lut_LC_16_4_2  (
            .in0(N__51753),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51493),
            .lcout(),
            .ltout(\ADC_VDC.n22124_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.SCLK_46_LC_16_4_3 .C_ON=1'b0;
    defparam \ADC_VDC.SCLK_46_LC_16_4_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.SCLK_46_LC_16_4_3 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \ADC_VDC.SCLK_46_LC_16_4_3  (
            .in0(N__42446),
            .in1(N__44262),
            .in2(N__41739),
            .in3(N__51208),
            .lcout(VDC_SCLK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__42363),
            .ce(),
            .sr(_gnd_net_));
    defparam i19347_2_lut_LC_16_5_7.C_ON=1'b0;
    defparam i19347_2_lut_LC_16_5_7.SEQ_MODE=4'b0000;
    defparam i19347_2_lut_LC_16_5_7.LUT_INIT=16'b1111111111001100;
    LogicCell40 i19347_2_lut_LC_16_5_7 (
            .in0(_gnd_net_),
            .in1(N__42183),
            .in2(_gnd_net_),
            .in3(N__57270),
            .lcout(n21557),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam flagcntwd_303_LC_16_6_0.C_ON=1'b0;
    defparam flagcntwd_303_LC_16_6_0.SEQ_MODE=4'b1000;
    defparam flagcntwd_303_LC_16_6_0.LUT_INIT=16'b1111111101010101;
    LogicCell40 flagcntwd_303_LC_16_6_0 (
            .in0(N__53979),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__54486),
            .lcout(flagcntwd),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55945),
            .ce(N__42099),
            .sr(N__42083));
    defparam i18460_2_lut_LC_16_6_1.C_ON=1'b0;
    defparam i18460_2_lut_LC_16_6_1.SEQ_MODE=4'b0000;
    defparam i18460_2_lut_LC_16_6_1.LUT_INIT=16'b1100110000000000;
    LogicCell40 i18460_2_lut_LC_16_6_1 (
            .in0(_gnd_net_),
            .in1(N__54379),
            .in2(_gnd_net_),
            .in3(N__53978),
            .lcout(),
            .ltout(n21187_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_277_LC_16_6_2.C_ON=1'b0;
    defparam i1_4_lut_adj_277_LC_16_6_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_277_LC_16_6_2.LUT_INIT=16'b1010101100000000;
    LogicCell40 i1_4_lut_adj_277_LC_16_6_2 (
            .in0(N__55238),
            .in1(N__54862),
            .in2(N__42102),
            .in3(N__55572),
            .lcout(n11605),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_186_LC_16_6_3.C_ON=1'b0;
    defparam i1_2_lut_adj_186_LC_16_6_3.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_186_LC_16_6_3.LUT_INIT=16'b0000000010101010;
    LogicCell40 i1_2_lut_adj_186_LC_16_6_3 (
            .in0(N__54859),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55235),
            .lcout(n80),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_56_LC_16_6_4.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_56_LC_16_6_4.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_56_LC_16_6_4.LUT_INIT=16'b1010101010100000;
    LogicCell40 i1_2_lut_3_lut_adj_56_LC_16_6_4 (
            .in0(N__55236),
            .in1(_gnd_net_),
            .in2(N__54502),
            .in3(N__54861),
            .lcout(n20578),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_243_LC_16_6_5.C_ON=1'b0;
    defparam i1_2_lut_adj_243_LC_16_6_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_243_LC_16_6_5.LUT_INIT=16'b1111111110101010;
    LogicCell40 i1_2_lut_adj_243_LC_16_6_5 (
            .in0(N__54860),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53977),
            .lcout(),
            .ltout(n11576_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_289_LC_16_6_6.C_ON=1'b0;
    defparam i1_4_lut_adj_289_LC_16_6_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_289_LC_16_6_6.LUT_INIT=16'b1010111000000000;
    LogicCell40 i1_4_lut_adj_289_LC_16_6_6 (
            .in0(N__55237),
            .in1(N__54485),
            .in2(N__42072),
            .in3(N__55571),
            .lcout(n12148),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_45_LC_16_6_7.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_45_LC_16_6_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_45_LC_16_6_7.LUT_INIT=16'b1111111101110111;
    LogicCell40 i1_2_lut_3_lut_adj_45_LC_16_6_7 (
            .in0(N__54858),
            .in1(N__54375),
            .in2(_gnd_net_),
            .in3(N__55234),
            .lcout(n21143),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i4_12317_12318_set_LC_16_7_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i4_12317_12318_set_LC_16_7_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i4_12317_12318_set_LC_16_7_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i4_12317_12318_set_LC_16_7_0  (
            .in0(N__56504),
            .in1(N__56487),
            .in2(_gnd_net_),
            .in3(N__57378),
            .lcout(\comm_spi.n14838 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__58337),
            .ce(),
            .sr(N__56421));
    defparam i12470_2_lut_LC_16_7_1.C_ON=1'b0;
    defparam i12470_2_lut_LC_16_7_1.SEQ_MODE=4'b0000;
    defparam i12470_2_lut_LC_16_7_1.LUT_INIT=16'b1100110000000000;
    LogicCell40 i12470_2_lut_LC_16_7_1 (
            .in0(_gnd_net_),
            .in1(N__55251),
            .in2(_gnd_net_),
            .in3(N__45059),
            .lcout(n14986),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12477_2_lut_LC_16_7_2.C_ON=1'b0;
    defparam i12477_2_lut_LC_16_7_2.SEQ_MODE=4'b0000;
    defparam i12477_2_lut_LC_16_7_2.LUT_INIT=16'b1010000010100000;
    LogicCell40 i12477_2_lut_LC_16_7_2 (
            .in0(N__48293),
            .in1(_gnd_net_),
            .in2(N__55358),
            .in3(_gnd_net_),
            .lcout(n14993),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i9391_1_lut_LC_16_7_4.C_ON=1'b0;
    defparam i9391_1_lut_LC_16_7_4.SEQ_MODE=4'b0000;
    defparam i9391_1_lut_LC_16_7_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 i9391_1_lut_LC_16_7_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44822),
            .lcout(n11910),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15273_2_lut_LC_16_7_6.C_ON=1'b0;
    defparam i15273_2_lut_LC_16_7_6.SEQ_MODE=4'b0000;
    defparam i15273_2_lut_LC_16_7_6.LUT_INIT=16'b1100110000000000;
    LogicCell40 i15273_2_lut_LC_16_7_6 (
            .in0(_gnd_net_),
            .in1(N__44992),
            .in2(_gnd_net_),
            .in3(N__44967),
            .lcout(n17773),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19029_2_lut_LC_16_7_7.C_ON=1'b0;
    defparam i19029_2_lut_LC_16_7_7.SEQ_MODE=4'b0000;
    defparam i19029_2_lut_LC_16_7_7.LUT_INIT=16'b1111111110101010;
    LogicCell40 i19029_2_lut_LC_16_7_7 (
            .in0(N__57271),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42588),
            .lcout(n21385),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22539_bdd_4_lut_LC_16_8_1.C_ON=1'b0;
    defparam n22539_bdd_4_lut_LC_16_8_1.SEQ_MODE=4'b0000;
    defparam n22539_bdd_4_lut_LC_16_8_1.LUT_INIT=16'b1010101011011000;
    LogicCell40 n22539_bdd_4_lut_LC_16_8_1 (
            .in0(N__43215),
            .in1(N__44071),
            .in2(N__42550),
            .in3(N__52447),
            .lcout(),
            .ltout(n22542_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i7_LC_16_8_2.C_ON=1'b0;
    defparam comm_tx_buf_i7_LC_16_8_2.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i7_LC_16_8_2.LUT_INIT=16'b1101100011011000;
    LogicCell40 comm_tx_buf_i7_LC_16_8_2 (
            .in0(N__52555),
            .in1(N__42483),
            .in2(N__42474),
            .in3(_gnd_net_),
            .lcout(comm_tx_buf_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55960),
            .ce(N__50341),
            .sr(N__50261));
    defparam mux_137_Mux_7_i4_3_lut_LC_16_8_4.C_ON=1'b0;
    defparam mux_137_Mux_7_i4_3_lut_LC_16_8_4.SEQ_MODE=4'b0000;
    defparam mux_137_Mux_7_i4_3_lut_LC_16_8_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_137_Mux_7_i4_3_lut_LC_16_8_4 (
            .in0(N__48048),
            .in1(N__44907),
            .in2(_gnd_net_),
            .in3(N__53073),
            .lcout(n4_adj_1580),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i19490_4_lut_3_lut_LC_16_8_5 .C_ON=1'b0;
    defparam \comm_spi.i19490_4_lut_3_lut_LC_16_8_5 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19490_4_lut_3_lut_LC_16_8_5 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \comm_spi.i19490_4_lut_3_lut_LC_16_8_5  (
            .in0(N__44311),
            .in1(N__42847),
            .in2(N__58156),
            .in3(_gnd_net_),
            .lcout(\comm_spi.n14811 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_100_2_lut_LC_16_8_6 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_100_2_lut_LC_16_8_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_100_2_lut_LC_16_8_6 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \comm_spi.RESET_I_0_100_2_lut_LC_16_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__42852),
            .in3(N__58108),
            .lcout(\comm_spi.data_tx_7__N_814 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_92_2_lut_LC_16_8_7 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_92_2_lut_LC_16_8_7 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_92_2_lut_LC_16_8_7 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \comm_spi.RESET_I_0_92_2_lut_LC_16_8_7  (
            .in0(N__58109),
            .in1(N__42851),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\comm_spi.data_tx_7__N_806 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_valid_85_LC_16_9_0 .C_ON=1'b0;
    defparam \comm_spi.data_valid_85_LC_16_9_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_valid_85_LC_16_9_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \comm_spi.data_valid_85_LC_16_9_0  (
            .in0(N__42801),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__42750),
            .lcout(comm_data_vld),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcomm_spi.data_valid_85C_net ),
            .ce(),
            .sr(N__58122));
    defparam comm_index_0__bdd_4_lut_19794_LC_16_10_0.C_ON=1'b0;
    defparam comm_index_0__bdd_4_lut_19794_LC_16_10_0.SEQ_MODE=4'b0000;
    defparam comm_index_0__bdd_4_lut_19794_LC_16_10_0.LUT_INIT=16'b1101100010101010;
    LogicCell40 comm_index_0__bdd_4_lut_19794_LC_16_10_0 (
            .in0(N__53047),
            .in1(N__49890),
            .in2(N__45975),
            .in3(N__52379),
            .lcout(),
            .ltout(n22551_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22551_bdd_4_lut_LC_16_10_1.C_ON=1'b0;
    defparam n22551_bdd_4_lut_LC_16_10_1.SEQ_MODE=4'b0000;
    defparam n22551_bdd_4_lut_LC_16_10_1.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22551_bdd_4_lut_LC_16_10_1 (
            .in0(N__52380),
            .in1(N__47759),
            .in2(N__42717),
            .in3(N__42709),
            .lcout(n22554),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_137_Mux_4_i4_3_lut_LC_16_10_2.C_ON=1'b0;
    defparam mux_137_Mux_4_i4_3_lut_LC_16_10_2.SEQ_MODE=4'b0000;
    defparam mux_137_Mux_4_i4_3_lut_LC_16_10_2.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_137_Mux_4_i4_3_lut_LC_16_10_2 (
            .in0(N__53048),
            .in1(N__47985),
            .in2(_gnd_net_),
            .in3(N__44856),
            .lcout(),
            .ltout(n4_adj_1582_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18558_4_lut_LC_16_10_3.C_ON=1'b0;
    defparam i18558_4_lut_LC_16_10_3.SEQ_MODE=4'b0000;
    defparam i18558_4_lut_LC_16_10_3.LUT_INIT=16'b0101000011011000;
    LogicCell40 i18558_4_lut_LC_16_10_3 (
            .in0(N__52381),
            .in1(N__53556),
            .in2(N__42648),
            .in3(N__53049),
            .lcout(),
            .ltout(n21285_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i4_LC_16_10_4.C_ON=1'b0;
    defparam comm_tx_buf_i4_LC_16_10_4.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i4_LC_16_10_4.LUT_INIT=16'b1111010110100000;
    LogicCell40 comm_tx_buf_i4_LC_16_10_4 (
            .in0(N__52523),
            .in1(_gnd_net_),
            .in2(N__42645),
            .in3(N__42642),
            .lcout(comm_tx_buf_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55981),
            .ce(N__50334),
            .sr(N__50243));
    defparam i19295_2_lut_3_lut_LC_16_10_5.C_ON=1'b0;
    defparam i19295_2_lut_3_lut_LC_16_10_5.SEQ_MODE=4'b0000;
    defparam i19295_2_lut_3_lut_LC_16_10_5.LUT_INIT=16'b0001000100000000;
    LogicCell40 i19295_2_lut_3_lut_LC_16_10_5 (
            .in0(N__52378),
            .in1(N__52522),
            .in2(_gnd_net_),
            .in3(N__49932),
            .lcout(),
            .ltout(n21474_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19_4_lut_adj_290_LC_16_10_6.C_ON=1'b0;
    defparam i19_4_lut_adj_290_LC_16_10_6.SEQ_MODE=4'b0000;
    defparam i19_4_lut_adj_290_LC_16_10_6.LUT_INIT=16'b0100000001110011;
    LogicCell40 i19_4_lut_adj_290_LC_16_10_6 (
            .in0(N__53046),
            .in1(N__54374),
            .in2(N__43113),
            .in3(N__48241),
            .lcout(),
            .ltout(n12_adj_1596_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_291_LC_16_10_7.C_ON=1'b0;
    defparam i1_3_lut_adj_291_LC_16_10_7.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_291_LC_16_10_7.LUT_INIT=16'b1111110000000000;
    LogicCell40 i1_3_lut_adj_291_LC_16_10_7 (
            .in0(_gnd_net_),
            .in1(N__48411),
            .in2(N__43110),
            .in3(N__48749),
            .lcout(n12184),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_1_i26_3_lut_LC_16_11_0.C_ON=1'b0;
    defparam mux_128_Mux_1_i26_3_lut_LC_16_11_0.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_1_i26_3_lut_LC_16_11_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_128_Mux_1_i26_3_lut_LC_16_11_0 (
            .in0(N__43107),
            .in1(N__57162),
            .in2(_gnd_net_),
            .in3(N__43085),
            .lcout(),
            .ltout(n26_adj_1694_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18633_4_lut_LC_16_11_1.C_ON=1'b0;
    defparam i18633_4_lut_LC_16_11_1.SEQ_MODE=4'b0000;
    defparam i18633_4_lut_LC_16_11_1.LUT_INIT=16'b0010001011110000;
    LogicCell40 i18633_4_lut_LC_16_11_1 (
            .in0(N__43059),
            .in1(N__57180),
            .in2(N__43050),
            .in3(N__46472),
            .lcout(n21360),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_0__bdd_4_lut_19852_LC_16_11_2.C_ON=1'b0;
    defparam comm_cmd_0__bdd_4_lut_19852_LC_16_11_2.SEQ_MODE=4'b0000;
    defparam comm_cmd_0__bdd_4_lut_19852_LC_16_11_2.LUT_INIT=16'b1101101011010000;
    LogicCell40 comm_cmd_0__bdd_4_lut_19852_LC_16_11_2 (
            .in0(N__46473),
            .in1(N__43047),
            .in2(N__57258),
            .in3(N__43002),
            .lcout(),
            .ltout(n22617_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22617_bdd_4_lut_LC_16_11_3.C_ON=1'b0;
    defparam n22617_bdd_4_lut_LC_16_11_3.SEQ_MODE=4'b0000;
    defparam n22617_bdd_4_lut_LC_16_11_3.LUT_INIT=16'b1111000010101100;
    LogicCell40 n22617_bdd_4_lut_LC_16_11_3 (
            .in0(N__42981),
            .in1(N__42953),
            .in2(N__42918),
            .in3(N__46474),
            .lcout(),
            .ltout(n22620_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18634_3_lut_LC_16_11_4.C_ON=1'b0;
    defparam i18634_3_lut_LC_16_11_4.SEQ_MODE=4'b0000;
    defparam i18634_3_lut_LC_16_11_4.LUT_INIT=16'b1111101001010000;
    LogicCell40 i18634_3_lut_LC_16_11_4 (
            .in0(N__47517),
            .in1(_gnd_net_),
            .in2(N__42915),
            .in3(N__42912),
            .lcout(),
            .ltout(n21361_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1563432_i1_3_lut_LC_16_11_5.C_ON=1'b0;
    defparam i1563432_i1_3_lut_LC_16_11_5.SEQ_MODE=4'b0000;
    defparam i1563432_i1_3_lut_LC_16_11_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 i1563432_i1_3_lut_LC_16_11_5 (
            .in0(_gnd_net_),
            .in1(N__42906),
            .in2(N__42891),
            .in3(N__47154),
            .lcout(),
            .ltout(n30_adj_1695_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_0__i1_LC_16_11_6.C_ON=1'b0;
    defparam comm_buf_0__i1_LC_16_11_6.SEQ_MODE=4'b1000;
    defparam comm_buf_0__i1_LC_16_11_6.LUT_INIT=16'b1111101001010000;
    LogicCell40 comm_buf_0__i1_LC_16_11_6 (
            .in0(N__54484),
            .in1(_gnd_net_),
            .in2(N__43341),
            .in3(N__49678),
            .lcout(comm_buf_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55994),
            .ce(N__43324),
            .sr(N__43274));
    defparam i41_4_lut_LC_16_11_7.C_ON=1'b0;
    defparam i41_4_lut_LC_16_11_7.SEQ_MODE=4'b0000;
    defparam i41_4_lut_LC_16_11_7.LUT_INIT=16'b0001100100100000;
    LogicCell40 i41_4_lut_LC_16_11_7 (
            .in0(N__46470),
            .in1(N__47153),
            .in2(N__57249),
            .in3(N__47516),
            .lcout(n24_adj_1639),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_0__bdd_4_lut_19784_LC_16_12_0.C_ON=1'b0;
    defparam comm_index_0__bdd_4_lut_19784_LC_16_12_0.SEQ_MODE=4'b0000;
    defparam comm_index_0__bdd_4_lut_19784_LC_16_12_0.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_index_0__bdd_4_lut_19784_LC_16_12_0 (
            .in0(N__45507),
            .in1(N__52445),
            .in2(N__48510),
            .in3(N__53066),
            .lcout(n22539),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15538_2_lut_3_lut_LC_16_12_1.C_ON=1'b0;
    defparam i15538_2_lut_3_lut_LC_16_12_1.SEQ_MODE=4'b0000;
    defparam i15538_2_lut_3_lut_LC_16_12_1.LUT_INIT=16'b0000000000100010;
    LogicCell40 i15538_2_lut_3_lut_LC_16_12_1 (
            .in0(N__45677),
            .in1(N__54777),
            .in2(_gnd_net_),
            .in3(N__54438),
            .lcout(n14_adj_1541),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_4_lut_4_lut_LC_16_12_2.C_ON=1'b0;
    defparam i1_4_lut_4_lut_4_lut_LC_16_12_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_4_lut_4_lut_LC_16_12_2.LUT_INIT=16'b1101100011001000;
    LogicCell40 i1_4_lut_4_lut_4_lut_LC_16_12_2 (
            .in0(N__54437),
            .in1(N__55247),
            .in2(N__54842),
            .in3(N__53962),
            .lcout(n12541),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_130_Mux_0_i30_3_lut_LC_16_12_3.C_ON=1'b0;
    defparam mux_130_Mux_0_i30_3_lut_LC_16_12_3.SEQ_MODE=4'b0000;
    defparam mux_130_Mux_0_i30_3_lut_LC_16_12_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_130_Mux_0_i30_3_lut_LC_16_12_3 (
            .in0(N__47254),
            .in1(N__43152),
            .in2(_gnd_net_),
            .in3(N__43137),
            .lcout(n30_adj_1531),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_342_Mux_3_i7_4_lut_4_lut_LC_16_12_4.C_ON=1'b0;
    defparam comm_state_3__I_0_342_Mux_3_i7_4_lut_4_lut_LC_16_12_4.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_342_Mux_3_i7_4_lut_4_lut_LC_16_12_4.LUT_INIT=16'b1111011111100110;
    LogicCell40 comm_state_3__I_0_342_Mux_3_i7_4_lut_4_lut_LC_16_12_4 (
            .in0(N__54439),
            .in1(N__54787),
            .in2(N__43125),
            .in3(N__53963),
            .lcout(n18070),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12449_2_lut_LC_16_12_5.C_ON=1'b0;
    defparam i12449_2_lut_LC_16_12_5.SEQ_MODE=4'b0000;
    defparam i12449_2_lut_LC_16_12_5.LUT_INIT=16'b1010101000000000;
    LogicCell40 i12449_2_lut_LC_16_12_5 (
            .in0(N__45170),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__55249),
            .lcout(n14965),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12456_2_lut_LC_16_12_6.C_ON=1'b0;
    defparam i12456_2_lut_LC_16_12_6.SEQ_MODE=4'b0000;
    defparam i12456_2_lut_LC_16_12_6.LUT_INIT=16'b1010101000000000;
    LogicCell40 i12456_2_lut_LC_16_12_6 (
            .in0(N__55250),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45902),
            .lcout(n14972),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i7_LC_16_12_7.C_ON=1'b0;
    defparam comm_buf_6__i7_LC_16_12_7.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i7_LC_16_12_7.LUT_INIT=16'b0100010011110000;
    LogicCell40 comm_buf_6__i7_LC_16_12_7 (
            .in0(N__55248),
            .in1(N__48588),
            .in2(N__43560),
            .in3(N__53142),
            .lcout(comm_buf_6_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56008),
            .ce(),
            .sr(_gnd_net_));
    defparam n22515_bdd_4_lut_LC_16_13_0.C_ON=1'b0;
    defparam n22515_bdd_4_lut_LC_16_13_0.SEQ_MODE=4'b0000;
    defparam n22515_bdd_4_lut_LC_16_13_0.LUT_INIT=16'b1100111011000010;
    LogicCell40 n22515_bdd_4_lut_LC_16_13_0 (
            .in0(N__43542),
            .in1(N__43410),
            .in2(N__47728),
            .in3(N__43518),
            .lcout(n22518),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19804_LC_16_13_1.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19804_LC_16_13_1.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19804_LC_16_13_1.LUT_INIT=16'b1110001011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_19804_LC_16_13_1 (
            .in0(N__43497),
            .in1(N__46484),
            .in2(N__43488),
            .in3(N__47712),
            .lcout(n22527),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_6_i26_3_lut_LC_16_13_2.C_ON=1'b0;
    defparam mux_129_Mux_6_i26_3_lut_LC_16_13_2.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_6_i26_3_lut_LC_16_13_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_129_Mux_6_i26_3_lut_LC_16_13_2 (
            .in0(N__43461),
            .in1(N__57250),
            .in2(_gnd_net_),
            .in3(N__43432),
            .lcout(),
            .ltout(n26_adj_1626_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19765_LC_16_13_3.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19765_LC_16_13_3.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19765_LC_16_13_3.LUT_INIT=16'b1011100011001100;
    LogicCell40 comm_cmd_1__bdd_4_lut_19765_LC_16_13_3 (
            .in0(N__53244),
            .in1(N__46483),
            .in2(N__43413),
            .in3(N__47711),
            .lcout(n22515),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22527_bdd_4_lut_LC_16_13_4.C_ON=1'b0;
    defparam n22527_bdd_4_lut_LC_16_13_4.SEQ_MODE=4'b0000;
    defparam n22527_bdd_4_lut_LC_16_13_4.LUT_INIT=16'b1111101001000100;
    LogicCell40 n22527_bdd_4_lut_LC_16_13_4 (
            .in0(N__47716),
            .in1(N__43404),
            .in2(N__43388),
            .in3(N__43359),
            .lcout(),
            .ltout(n22530_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1570668_i1_3_lut_LC_16_13_5.C_ON=1'b0;
    defparam i1570668_i1_3_lut_LC_16_13_5.SEQ_MODE=4'b0000;
    defparam i1570668_i1_3_lut_LC_16_13_5.LUT_INIT=16'b1111110000110000;
    LogicCell40 i1570668_i1_3_lut_LC_16_13_5 (
            .in0(_gnd_net_),
            .in1(N__47256),
            .in2(N__43353),
            .in3(N__43350),
            .lcout(),
            .ltout(n30_adj_1627_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i6_LC_16_13_6.C_ON=1'b0;
    defparam comm_buf_1__i6_LC_16_13_6.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i6_LC_16_13_6.LUT_INIT=16'b1100110011110000;
    LogicCell40 comm_buf_1__i6_LC_16_13_6 (
            .in0(_gnd_net_),
            .in1(N__53217),
            .in2(N__43344),
            .in3(N__54542),
            .lcout(comm_buf_1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56024),
            .ce(N__45209),
            .sr(N__43962));
    defparam mux_129_Mux_0_i26_3_lut_LC_16_14_0.C_ON=1'b0;
    defparam mux_129_Mux_0_i26_3_lut_LC_16_14_0.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_0_i26_3_lut_LC_16_14_0.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_129_Mux_0_i26_3_lut_LC_16_14_0 (
            .in0(N__43869),
            .in1(N__57130),
            .in2(_gnd_net_),
            .in3(N__43845),
            .lcout(),
            .ltout(n26_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18534_4_lut_LC_16_14_1.C_ON=1'b0;
    defparam i18534_4_lut_LC_16_14_1.SEQ_MODE=4'b0000;
    defparam i18534_4_lut_LC_16_14_1.LUT_INIT=16'b0101000011011000;
    LogicCell40 i18534_4_lut_LC_16_14_1 (
            .in0(N__46482),
            .in1(N__43818),
            .in2(N__43803),
            .in3(N__57131),
            .lcout(),
            .ltout(n21261_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_2__bdd_4_lut_19814_LC_16_14_2.C_ON=1'b0;
    defparam comm_cmd_2__bdd_4_lut_19814_LC_16_14_2.SEQ_MODE=4'b0000;
    defparam comm_cmd_2__bdd_4_lut_19814_LC_16_14_2.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_cmd_2__bdd_4_lut_19814_LC_16_14_2 (
            .in0(N__43626),
            .in1(N__47196),
            .in2(N__43800),
            .in3(N__47717),
            .lcout(),
            .ltout(n22563_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22563_bdd_4_lut_LC_16_14_3.C_ON=1'b0;
    defparam n22563_bdd_4_lut_LC_16_14_3.SEQ_MODE=4'b0000;
    defparam n22563_bdd_4_lut_LC_16_14_3.LUT_INIT=16'b1110001111100000;
    LogicCell40 n22563_bdd_4_lut_LC_16_14_3 (
            .in0(N__43683),
            .in1(N__47257),
            .in2(N__43797),
            .in3(N__43794),
            .lcout(),
            .ltout(n22566_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i0_LC_16_14_4.C_ON=1'b0;
    defparam comm_buf_1__i0_LC_16_14_4.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i0_LC_16_14_4.LUT_INIT=16'b1100110011110000;
    LogicCell40 comm_buf_1__i0_LC_16_14_4 (
            .in0(_gnd_net_),
            .in1(N__48697),
            .in2(N__43785),
            .in3(N__54543),
            .lcout(comm_buf_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56039),
            .ce(N__45194),
            .sr(N__44001));
    defparam mux_129_Mux_0_i19_3_lut_LC_16_14_5.C_ON=1'b0;
    defparam mux_129_Mux_0_i19_3_lut_LC_16_14_5.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_0_i19_3_lut_LC_16_14_5.LUT_INIT=16'b1101100011011000;
    LogicCell40 mux_129_Mux_0_i19_3_lut_LC_16_14_5 (
            .in0(N__57129),
            .in1(N__43782),
            .in2(N__43757),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(n19_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18531_3_lut_LC_16_14_6.C_ON=1'b0;
    defparam i18531_3_lut_LC_16_14_6.SEQ_MODE=4'b0000;
    defparam i18531_3_lut_LC_16_14_6.LUT_INIT=16'b1010101011110000;
    LogicCell40 i18531_3_lut_LC_16_14_6 (
            .in0(N__43710),
            .in1(_gnd_net_),
            .in2(N__43686),
            .in3(N__46481),
            .lcout(n21258),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18533_3_lut_LC_16_14_7.C_ON=1'b0;
    defparam i18533_3_lut_LC_16_14_7.SEQ_MODE=4'b0000;
    defparam i18533_3_lut_LC_16_14_7.LUT_INIT=16'b1110111001000100;
    LogicCell40 i18533_3_lut_LC_16_14_7 (
            .in0(N__46480),
            .in1(N__43677),
            .in2(_gnd_net_),
            .in3(N__43656),
            .lcout(n21260),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22431_bdd_4_lut_LC_16_15_0.C_ON=1'b0;
    defparam n22431_bdd_4_lut_LC_16_15_0.SEQ_MODE=4'b0000;
    defparam n22431_bdd_4_lut_LC_16_15_0.LUT_INIT=16'b1110111001010000;
    LogicCell40 n22431_bdd_4_lut_LC_16_15_0 (
            .in0(N__47722),
            .in1(N__43613),
            .in2(N__43587),
            .in3(N__43575),
            .lcout(n22434),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_1_i26_3_lut_LC_16_15_2.C_ON=1'b0;
    defparam mux_129_Mux_1_i26_3_lut_LC_16_15_2.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_1_i26_3_lut_LC_16_15_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_129_Mux_1_i26_3_lut_LC_16_15_2 (
            .in0(N__44217),
            .in1(N__57251),
            .in2(_gnd_net_),
            .in3(N__44199),
            .lcout(),
            .ltout(n26_adj_1653_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_1__bdd_4_lut_19755_LC_16_15_3.C_ON=1'b0;
    defparam comm_cmd_1__bdd_4_lut_19755_LC_16_15_3.SEQ_MODE=4'b0000;
    defparam comm_cmd_1__bdd_4_lut_19755_LC_16_15_3.LUT_INIT=16'b1101100010101010;
    LogicCell40 comm_cmd_1__bdd_4_lut_19755_LC_16_15_3 (
            .in0(N__46476),
            .in1(N__57291),
            .in2(N__44175),
            .in3(N__47723),
            .lcout(),
            .ltout(n22497_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22497_bdd_4_lut_LC_16_15_4.C_ON=1'b0;
    defparam n22497_bdd_4_lut_LC_16_15_4.SEQ_MODE=4'b0000;
    defparam n22497_bdd_4_lut_LC_16_15_4.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22497_bdd_4_lut_LC_16_15_4 (
            .in0(N__47724),
            .in1(N__44172),
            .in2(N__44151),
            .in3(N__44148),
            .lcout(),
            .ltout(n22500_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1567653_i1_3_lut_LC_16_15_5.C_ON=1'b0;
    defparam i1567653_i1_3_lut_LC_16_15_5.SEQ_MODE=4'b0000;
    defparam i1567653_i1_3_lut_LC_16_15_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 i1567653_i1_3_lut_LC_16_15_5 (
            .in0(_gnd_net_),
            .in1(N__44127),
            .in2(N__44121),
            .in3(N__47253),
            .lcout(),
            .ltout(n30_adj_1654_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i1_LC_16_15_6.C_ON=1'b0;
    defparam comm_buf_1__i1_LC_16_15_6.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i1_LC_16_15_6.LUT_INIT=16'b1111110000110000;
    LogicCell40 comm_buf_1__i1_LC_16_15_6 (
            .in0(_gnd_net_),
            .in1(N__54541),
            .in2(N__44118),
            .in3(N__49722),
            .lcout(comm_buf_1_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56055),
            .ce(N__45211),
            .sr(N__44014));
    defparam i1_2_lut_4_lut_adj_230_LC_16_15_7.C_ON=1'b0;
    defparam i1_2_lut_4_lut_adj_230_LC_16_15_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_4_lut_adj_230_LC_16_15_7.LUT_INIT=16'b1111111111111110;
    LogicCell40 i1_2_lut_4_lut_adj_230_LC_16_15_7 (
            .in0(N__46475),
            .in1(N__47252),
            .in2(N__44115),
            .in3(N__47721),
            .lcout(n68),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_1__i7_LC_16_16_0.C_ON=1'b0;
    defparam comm_buf_1__i7_LC_16_16_0.SEQ_MODE=4'b1000;
    defparam comm_buf_1__i7_LC_16_16_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_1__i7_LC_16_16_0 (
            .in0(N__54567),
            .in1(N__48599),
            .in2(_gnd_net_),
            .in3(N__46971),
            .lcout(comm_buf_1_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56067),
            .ce(N__45210),
            .sr(N__44013));
    defparam \SIG_DDS.i19394_4_lut_LC_16_17_4 .C_ON=1'b0;
    defparam \SIG_DDS.i19394_4_lut_LC_16_17_4 .SEQ_MODE=4'b0000;
    defparam \SIG_DDS.i19394_4_lut_LC_16_17_4 .LUT_INIT=16'b1010101000100110;
    LogicCell40 \SIG_DDS.i19394_4_lut_LC_16_17_4  (
            .in0(N__44657),
            .in1(N__44748),
            .in2(N__43943),
            .in3(N__44376),
            .lcout(\SIG_DDS.n12895 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15221_2_lut_2_lut_LC_16_17_5.C_ON=1'b0;
    defparam i15221_2_lut_2_lut_LC_16_17_5.SEQ_MODE=4'b0000;
    defparam i15221_2_lut_2_lut_LC_16_17_5.LUT_INIT=16'b0101010100000000;
    LogicCell40 i15221_2_lut_2_lut_LC_16_17_5 (
            .in0(N__44829),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44799),
            .lcout(CONT_SD),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \SIG_DDS.dds_state_i1_LC_16_18_0 .C_ON=1'b0;
    defparam \SIG_DDS.dds_state_i1_LC_16_18_0 .SEQ_MODE=4'b1000;
    defparam \SIG_DDS.dds_state_i1_LC_16_18_0 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \SIG_DDS.dds_state_i1_LC_16_18_0  (
            .in0(N__44754),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44668),
            .lcout(dds_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56087),
            .ce(N__44543),
            .sr(N__44503));
    defparam \comm_spi.i12293_3_lut_LC_17_2_4 .C_ON=1'b0;
    defparam \comm_spi.i12293_3_lut_LC_17_2_4 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i12293_3_lut_LC_17_2_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \comm_spi.i12293_3_lut_LC_17_2_4  (
            .in0(N__44343),
            .in1(N__44337),
            .in2(_gnd_net_),
            .in3(N__44330),
            .lcout(ICE_SPI_MISO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i19395_4_lut_4_lut_LC_17_4_2 .C_ON=1'b0;
    defparam \ADC_VDC.i19395_4_lut_4_lut_LC_17_4_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i19395_4_lut_4_lut_LC_17_4_2 .LUT_INIT=16'b1111101011111001;
    LogicCell40 \ADC_VDC.i19395_4_lut_4_lut_LC_17_4_2  (
            .in0(N__51492),
            .in1(N__51895),
            .in2(N__51761),
            .in3(N__51213),
            .lcout(\ADC_VDC.n11895 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i19480_4_lut_3_lut_LC_17_4_6 .C_ON=1'b0;
    defparam \comm_spi.i19480_4_lut_3_lut_LC_17_4_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19480_4_lut_3_lut_LC_17_4_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \comm_spi.i19480_4_lut_3_lut_LC_17_4_6  (
            .in0(N__44256),
            .in1(N__48140),
            .in2(_gnd_net_),
            .in3(N__58159),
            .lcout(\comm_spi.n23086 ),
            .ltout(\comm_spi.n23086_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i12285_3_lut_LC_17_4_7 .C_ON=1'b0;
    defparam \comm_spi.i12285_3_lut_LC_17_4_7 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i12285_3_lut_LC_17_4_7 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \comm_spi.i12285_3_lut_LC_17_4_7  (
            .in0(N__46653),
            .in1(N__44247),
            .in2(N__44250),
            .in3(_gnd_net_),
            .lcout(\comm_spi.iclk ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.iclk_40_12283_12284_set_LC_17_5_0 .C_ON=1'b0;
    defparam \comm_spi.iclk_40_12283_12284_set_LC_17_5_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.iclk_40_12283_12284_set_LC_17_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \comm_spi.iclk_40_12283_12284_set_LC_17_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48141),
            .lcout(\comm_spi.n14804 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55946),
            .ce(),
            .sr(N__46647));
    defparam i19131_4_lut_LC_17_6_2.C_ON=1'b0;
    defparam i19131_4_lut_LC_17_6_2.SEQ_MODE=4'b0000;
    defparam i19131_4_lut_LC_17_6_2.LUT_INIT=16'b1000000000000000;
    LogicCell40 i19131_4_lut_LC_17_6_2 (
            .in0(N__44241),
            .in1(N__47270),
            .in2(N__44235),
            .in3(N__47642),
            .lcout(n21481),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i19510_4_lut_3_lut_LC_17_6_4 .C_ON=1'b0;
    defparam \comm_spi.i19510_4_lut_3_lut_LC_17_6_4 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19510_4_lut_3_lut_LC_17_6_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \comm_spi.i19510_4_lut_3_lut_LC_17_6_4  (
            .in0(N__56503),
            .in1(N__56140),
            .in2(_gnd_net_),
            .in3(N__57988),
            .lcout(\comm_spi.n23101 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i19485_4_lut_3_lut_LC_17_6_6 .C_ON=1'b0;
    defparam \comm_spi.i19485_4_lut_3_lut_LC_17_6_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19485_4_lut_3_lut_LC_17_6_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \comm_spi.i19485_4_lut_3_lut_LC_17_6_6  (
            .in0(N__45016),
            .in1(N__50869),
            .in2(_gnd_net_),
            .in3(N__57987),
            .lcout(\comm_spi.n23092 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_cnt_3761_3762__i2_LC_17_7_0.C_ON=1'b0;
    defparam clk_cnt_3761_3762__i2_LC_17_7_0.SEQ_MODE=4'b1000;
    defparam clk_cnt_3761_3762__i2_LC_17_7_0.LUT_INIT=16'b0101010110101010;
    LogicCell40 clk_cnt_3761_3762__i2_LC_17_7_0 (
            .in0(N__44969),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44993),
            .lcout(clk_cnt_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50791),
            .ce(),
            .sr(N__44949));
    defparam clk_cnt_3761_3762__i1_LC_17_7_1.C_ON=1'b0;
    defparam clk_cnt_3761_3762__i1_LC_17_7_1.SEQ_MODE=4'b1000;
    defparam clk_cnt_3761_3762__i1_LC_17_7_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 clk_cnt_3761_3762__i1_LC_17_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44968),
            .lcout(clk_cnt_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__50791),
            .ce(),
            .sr(N__44949));
    defparam comm_buf_4__i0_LC_17_8_0.C_ON=1'b0;
    defparam comm_buf_4__i0_LC_17_8_0.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i0_LC_17_8_0.LUT_INIT=16'b1110111000100010;
    LogicCell40 comm_buf_4__i0_LC_17_8_0 (
            .in0(N__44940),
            .in1(N__54335),
            .in2(_gnd_net_),
            .in3(N__48703),
            .lcout(comm_buf_4_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55970),
            .ce(N__45060),
            .sr(N__45090));
    defparam comm_buf_4__i7_LC_17_8_1.C_ON=1'b0;
    defparam comm_buf_4__i7_LC_17_8_1.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i7_LC_17_8_1.LUT_INIT=16'b1111010110100000;
    LogicCell40 comm_buf_4__i7_LC_17_8_1 (
            .in0(N__54334),
            .in1(_gnd_net_),
            .in2(N__48596),
            .in3(N__44922),
            .lcout(comm_buf_4_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55970),
            .ce(N__45060),
            .sr(N__45090));
    defparam comm_buf_4__i6_LC_17_8_2.C_ON=1'b0;
    defparam comm_buf_4__i6_LC_17_8_2.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i6_LC_17_8_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_4__i6_LC_17_8_2 (
            .in0(N__53227),
            .in1(N__44901),
            .in2(_gnd_net_),
            .in3(N__54338),
            .lcout(comm_buf_4_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55970),
            .ce(N__45060),
            .sr(N__45090));
    defparam comm_buf_4__i5_LC_17_8_3.C_ON=1'b0;
    defparam comm_buf_4__i5_LC_17_8_3.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i5_LC_17_8_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_4__i5_LC_17_8_3 (
            .in0(N__54333),
            .in1(N__53331),
            .in2(_gnd_net_),
            .in3(N__44889),
            .lcout(comm_buf_4_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55970),
            .ce(N__45060),
            .sr(N__45090));
    defparam comm_buf_4__i4_LC_17_8_4.C_ON=1'b0;
    defparam comm_buf_4__i4_LC_17_8_4.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i4_LC_17_8_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_4__i4_LC_17_8_4 (
            .in0(N__53619),
            .in1(N__44874),
            .in2(_gnd_net_),
            .in3(N__54337),
            .lcout(comm_buf_4_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55970),
            .ce(N__45060),
            .sr(N__45090));
    defparam comm_buf_4__i3_LC_17_8_5.C_ON=1'b0;
    defparam comm_buf_4__i3_LC_17_8_5.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i3_LC_17_8_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_4__i3_LC_17_8_5 (
            .in0(N__54332),
            .in1(N__49867),
            .in2(_gnd_net_),
            .in3(N__44847),
            .lcout(comm_buf_4_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55970),
            .ce(N__45060),
            .sr(N__45090));
    defparam comm_buf_4__i2_LC_17_8_6.C_ON=1'b0;
    defparam comm_buf_4__i2_LC_17_8_6.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i2_LC_17_8_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_4__i2_LC_17_8_6 (
            .in0(N__50145),
            .in1(N__45126),
            .in2(_gnd_net_),
            .in3(N__54336),
            .lcout(comm_buf_4_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55970),
            .ce(N__45060),
            .sr(N__45090));
    defparam comm_buf_4__i1_LC_17_8_7.C_ON=1'b0;
    defparam comm_buf_4__i1_LC_17_8_7.SEQ_MODE=4'b1000;
    defparam comm_buf_4__i1_LC_17_8_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_4__i1_LC_17_8_7 (
            .in0(N__54331),
            .in1(N__49717),
            .in2(_gnd_net_),
            .in3(N__45108),
            .lcout(comm_buf_4_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55970),
            .ce(N__45060),
            .sr(N__45090));
    defparam i18541_4_lut_LC_17_9_0.C_ON=1'b0;
    defparam i18541_4_lut_LC_17_9_0.SEQ_MODE=4'b0000;
    defparam i18541_4_lut_LC_17_9_0.LUT_INIT=16'b1110111011110000;
    LogicCell40 i18541_4_lut_LC_17_9_0 (
            .in0(N__52151),
            .in1(N__45075),
            .in2(N__45069),
            .in3(N__54841),
            .lcout(),
            .ltout(n21268_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_i0_LC_17_9_1.C_ON=1'b0;
    defparam comm_state_i0_LC_17_9_1.SEQ_MODE=4'b1000;
    defparam comm_state_i0_LC_17_9_1.LUT_INIT=16'b0011001111110000;
    LogicCell40 comm_state_i0_LC_17_9_1 (
            .in0(_gnd_net_),
            .in1(N__49374),
            .in2(N__45078),
            .in3(N__55066),
            .lcout(comm_state_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55982),
            .ce(N__48453),
            .sr(_gnd_net_));
    defparam i19367_3_lut_LC_17_9_2.C_ON=1'b0;
    defparam i19367_3_lut_LC_17_9_2.SEQ_MODE=4'b0000;
    defparam i19367_3_lut_LC_17_9_2.LUT_INIT=16'b1110111000000000;
    LogicCell40 i19367_3_lut_LC_17_9_2 (
            .in0(N__50003),
            .in1(N__46037),
            .in2(_gnd_net_),
            .in3(N__54191),
            .lcout(n22094),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18539_3_lut_LC_17_9_3.C_ON=1'b0;
    defparam i18539_3_lut_LC_17_9_3.SEQ_MODE=4'b0000;
    defparam i18539_3_lut_LC_17_9_3.LUT_INIT=16'b1010101011011101;
    LogicCell40 i18539_3_lut_LC_17_9_3 (
            .in0(N__54192),
            .in1(N__52782),
            .in2(_gnd_net_),
            .in3(N__53869),
            .lcout(n21266),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_301_LC_17_9_4.C_ON=1'b0;
    defparam i1_4_lut_adj_301_LC_17_9_4.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_301_LC_17_9_4.LUT_INIT=16'b1010001010100000;
    LogicCell40 i1_4_lut_adj_301_LC_17_9_4 (
            .in0(N__48764),
            .in1(N__53071),
            .in2(N__45390),
            .in3(N__45039),
            .lcout(n12407),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_4_lut_adj_304_LC_17_9_5.C_ON=1'b0;
    defparam i1_3_lut_4_lut_adj_304_LC_17_9_5.SEQ_MODE=4'b0000;
    defparam i1_3_lut_4_lut_adj_304_LC_17_9_5.LUT_INIT=16'b0000000000010000;
    LogicCell40 i1_3_lut_4_lut_adj_304_LC_17_9_5 (
            .in0(N__52783),
            .in1(N__50002),
            .in2(N__52855),
            .in3(N__53868),
            .lcout(n21085),
            .ltout(n21085_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_262_LC_17_9_6.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_262_LC_17_9_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_262_LC_17_9_6.LUT_INIT=16'b0101000000000000;
    LogicCell40 i1_2_lut_3_lut_adj_262_LC_17_9_6 (
            .in0(N__52446),
            .in1(_gnd_net_),
            .in2(N__45042),
            .in3(N__52553),
            .lcout(n19188),
            .ltout(n19188_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_309_LC_17_9_7.C_ON=1'b0;
    defparam i1_4_lut_adj_309_LC_17_9_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_309_LC_17_9_7.LUT_INIT=16'b1110110000000000;
    LogicCell40 i1_4_lut_adj_309_LC_17_9_7 (
            .in0(N__53072),
            .in1(N__45388),
            .in2(N__45360),
            .in3(N__48765),
            .lcout(n12431),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_0__bdd_4_lut_LC_17_10_0.C_ON=1'b0;
    defparam comm_index_0__bdd_4_lut_LC_17_10_0.SEQ_MODE=4'b0000;
    defparam comm_index_0__bdd_4_lut_LC_17_10_0.LUT_INIT=16'b1110010010101010;
    LogicCell40 comm_index_0__bdd_4_lut_LC_17_10_0 (
            .in0(N__52990),
            .in1(N__45948),
            .in2(N__49776),
            .in3(N__52409),
            .lcout(),
            .ltout(n22557_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22557_bdd_4_lut_LC_17_10_1.C_ON=1'b0;
    defparam n22557_bdd_4_lut_LC_17_10_1.SEQ_MODE=4'b0000;
    defparam n22557_bdd_4_lut_LC_17_10_1.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22557_bdd_4_lut_LC_17_10_1 (
            .in0(N__52410),
            .in1(N__45334),
            .in2(N__45285),
            .in3(N__45280),
            .lcout(n22560),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_137_Mux_3_i4_3_lut_LC_17_10_2.C_ON=1'b0;
    defparam mux_137_Mux_3_i4_3_lut_LC_17_10_2.SEQ_MODE=4'b0000;
    defparam mux_137_Mux_3_i4_3_lut_LC_17_10_2.LUT_INIT=16'b1111010110100000;
    LogicCell40 mux_137_Mux_3_i4_3_lut_LC_17_10_2 (
            .in0(N__52991),
            .in1(_gnd_net_),
            .in2(N__47961),
            .in3(N__45252),
            .lcout(),
            .ltout(n4_adj_1583_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18561_4_lut_LC_17_10_3.C_ON=1'b0;
    defparam i18561_4_lut_LC_17_10_3.SEQ_MODE=4'b0000;
    defparam i18561_4_lut_LC_17_10_3.LUT_INIT=16'b0101000011011000;
    LogicCell40 i18561_4_lut_LC_17_10_3 (
            .in0(N__52411),
            .in1(N__46620),
            .in2(N__45243),
            .in3(N__52992),
            .lcout(),
            .ltout(n21288_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i3_LC_17_10_4.C_ON=1'b0;
    defparam comm_tx_buf_i3_LC_17_10_4.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i3_LC_17_10_4.LUT_INIT=16'b1111000011001100;
    LogicCell40 comm_tx_buf_i3_LC_17_10_4 (
            .in0(_gnd_net_),
            .in1(N__45240),
            .in2(N__45234),
            .in3(N__52521),
            .lcout(comm_tx_buf_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55995),
            .ce(N__50333),
            .sr(N__50254));
    defparam i19129_3_lut_4_lut_LC_17_10_5.C_ON=1'b0;
    defparam i19129_3_lut_4_lut_LC_17_10_5.SEQ_MODE=4'b0000;
    defparam i19129_3_lut_4_lut_LC_17_10_5.LUT_INIT=16'b0000010000000000;
    LogicCell40 i19129_3_lut_4_lut_LC_17_10_5 (
            .in0(N__52520),
            .in1(N__52989),
            .in2(N__52439),
            .in3(N__49931),
            .lcout(),
            .ltout(n21477_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i48_4_lut_LC_17_10_6.C_ON=1'b0;
    defparam i48_4_lut_LC_17_10_6.SEQ_MODE=4'b0000;
    defparam i48_4_lut_LC_17_10_6.LUT_INIT=16'b1100000011100010;
    LogicCell40 i48_4_lut_LC_17_10_6 (
            .in0(N__45231),
            .in1(N__54440),
            .in2(N__45219),
            .in3(N__48257),
            .lcout(),
            .ltout(n44_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_294_LC_17_10_7.C_ON=1'b0;
    defparam i1_3_lut_adj_294_LC_17_10_7.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_294_LC_17_10_7.LUT_INIT=16'b1111110000000000;
    LogicCell40 i1_3_lut_adj_294_LC_17_10_7 (
            .in0(_gnd_net_),
            .in1(N__48409),
            .in2(N__45216),
            .in3(N__48742),
            .lcout(n12260),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_137_Mux_2_i1_3_lut_LC_17_11_0.C_ON=1'b0;
    defparam mux_137_Mux_2_i1_3_lut_LC_17_11_0.SEQ_MODE=4'b0000;
    defparam mux_137_Mux_2_i1_3_lut_LC_17_11_0.LUT_INIT=16'b1100110010101010;
    LogicCell40 mux_137_Mux_2_i1_3_lut_LC_17_11_0 (
            .in0(N__45829),
            .in1(N__45475),
            .in2(_gnd_net_),
            .in3(N__53065),
            .lcout(),
            .ltout(n1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i2_LC_17_11_1.C_ON=1'b0;
    defparam comm_tx_buf_i2_LC_17_11_1.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i2_LC_17_11_1.LUT_INIT=16'b1110111001010000;
    LogicCell40 comm_tx_buf_i2_LC_17_11_1 (
            .in0(N__52560),
            .in1(N__45420),
            .in2(N__45423),
            .in3(N__45396),
            .lcout(comm_tx_buf_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56009),
            .ce(N__50355),
            .sr(N__50265));
    defparam i19154_2_lut_LC_17_11_2.C_ON=1'b0;
    defparam i19154_2_lut_LC_17_11_2.SEQ_MODE=4'b0000;
    defparam i19154_2_lut_LC_17_11_2.LUT_INIT=16'b0000000010101010;
    LogicCell40 i19154_2_lut_LC_17_11_2 (
            .in0(N__50072),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__53062),
            .lcout(n21528),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_137_Mux_2_i2_3_lut_LC_17_11_3.C_ON=1'b0;
    defparam mux_137_Mux_2_i2_3_lut_LC_17_11_3.SEQ_MODE=4'b0000;
    defparam mux_137_Mux_2_i2_3_lut_LC_17_11_3.LUT_INIT=16'b1111010110100000;
    LogicCell40 mux_137_Mux_2_i2_3_lut_LC_17_11_3 (
            .in0(N__53064),
            .in1(_gnd_net_),
            .in2(N__49755),
            .in3(N__45927),
            .lcout(n2_adj_1584),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_137_Mux_2_i4_3_lut_LC_17_11_4.C_ON=1'b0;
    defparam mux_137_Mux_2_i4_3_lut_LC_17_11_4.SEQ_MODE=4'b0000;
    defparam mux_137_Mux_2_i4_3_lut_LC_17_11_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_137_Mux_2_i4_3_lut_LC_17_11_4 (
            .in0(N__47937),
            .in1(N__45414),
            .in2(_gnd_net_),
            .in3(N__53063),
            .lcout(),
            .ltout(n4_adj_1585_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_1__bdd_4_lut_LC_17_11_5.C_ON=1'b0;
    defparam comm_index_1__bdd_4_lut_LC_17_11_5.SEQ_MODE=4'b0000;
    defparam comm_index_1__bdd_4_lut_LC_17_11_5.LUT_INIT=16'b1101110110100000;
    LogicCell40 comm_index_1__bdd_4_lut_LC_17_11_5 (
            .in0(N__52559),
            .in1(N__45405),
            .in2(N__45399),
            .in3(N__52444),
            .lcout(n22491),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_281_LC_17_11_6.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_281_LC_17_11_6.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_281_LC_17_11_6.LUT_INIT=16'b0010001000000000;
    LogicCell40 i1_2_lut_3_lut_adj_281_LC_17_11_6 (
            .in0(N__52443),
            .in1(N__52558),
            .in2(_gnd_net_),
            .in3(N__49943),
            .lcout(),
            .ltout(n19193_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_299_LC_17_11_7.C_ON=1'b0;
    defparam i1_4_lut_adj_299_LC_17_11_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_299_LC_17_11_7.LUT_INIT=16'b1110110000000000;
    LogicCell40 i1_4_lut_adj_299_LC_17_11_7 (
            .in0(N__53061),
            .in1(N__45389),
            .in2(N__45363),
            .in3(N__48763),
            .lcout(n12353),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i0_LC_17_12_0.C_ON=1'b0;
    defparam comm_tx_buf_i0_LC_17_12_0.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i0_LC_17_12_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_tx_buf_i0_LC_17_12_0 (
            .in0(N__45687),
            .in1(N__45549),
            .in2(_gnd_net_),
            .in3(N__52557),
            .lcout(comm_tx_buf_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56025),
            .ce(N__50305),
            .sr(N__50231));
    defparam i18546_4_lut_LC_17_12_1.C_ON=1'b0;
    defparam i18546_4_lut_LC_17_12_1.SEQ_MODE=4'b0000;
    defparam i18546_4_lut_LC_17_12_1.LUT_INIT=16'b0100010011100100;
    LogicCell40 i18546_4_lut_LC_17_12_1 (
            .in0(N__52434),
            .in1(N__50037),
            .in2(N__46641),
            .in3(N__53052),
            .lcout(n21273),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_0__bdd_4_lut_19779_LC_17_12_2.C_ON=1'b0;
    defparam comm_index_0__bdd_4_lut_19779_LC_17_12_2.SEQ_MODE=4'b0000;
    defparam comm_index_0__bdd_4_lut_19779_LC_17_12_2.LUT_INIT=16'b1110010010101010;
    LogicCell40 comm_index_0__bdd_4_lut_19779_LC_17_12_2 (
            .in0(N__53051),
            .in1(N__45525),
            .in2(N__48624),
            .in3(N__52432),
            .lcout(),
            .ltout(n22533_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22533_bdd_4_lut_LC_17_12_3.C_ON=1'b0;
    defparam n22533_bdd_4_lut_LC_17_12_3.SEQ_MODE=4'b0000;
    defparam n22533_bdd_4_lut_LC_17_12_3.LUT_INIT=16'b1110010111100000;
    LogicCell40 n22533_bdd_4_lut_LC_17_12_3 (
            .in0(N__52433),
            .in1(N__45681),
            .in2(N__45651),
            .in3(N__45621),
            .lcout(n22536),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19137_3_lut_4_lut_LC_17_12_5.C_ON=1'b0;
    defparam i19137_3_lut_4_lut_LC_17_12_5.SEQ_MODE=4'b0000;
    defparam i19137_3_lut_4_lut_LC_17_12_5.LUT_INIT=16'b0001000000000000;
    LogicCell40 i19137_3_lut_4_lut_LC_17_12_5 (
            .in0(N__52556),
            .in1(N__53050),
            .in2(N__52448),
            .in3(N__49942),
            .lcout(),
            .ltout(n21497_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i39_4_lut_LC_17_12_6.C_ON=1'b0;
    defparam i39_4_lut_LC_17_12_6.SEQ_MODE=4'b0000;
    defparam i39_4_lut_LC_17_12_6.LUT_INIT=16'b1100000011100010;
    LogicCell40 i39_4_lut_LC_17_12_6 (
            .in0(N__45543),
            .in1(N__54525),
            .in2(N__45537),
            .in3(N__48258),
            .lcout(),
            .ltout(n34_adj_1649_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_296_LC_17_12_7.C_ON=1'b0;
    defparam i1_3_lut_adj_296_LC_17_12_7.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_296_LC_17_12_7.LUT_INIT=16'b1010101010100000;
    LogicCell40 i1_3_lut_adj_296_LC_17_12_7 (
            .in0(N__48750),
            .in1(_gnd_net_),
            .in2(N__45534),
            .in3(N__48410),
            .lcout(n12314),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_2__i0_LC_17_13_0.C_ON=1'b0;
    defparam comm_buf_2__i0_LC_17_13_0.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i0_LC_17_13_0.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_2__i0_LC_17_13_0 (
            .in0(N__48699),
            .in1(N__45531),
            .in2(_gnd_net_),
            .in3(N__54548),
            .lcout(comm_buf_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56040),
            .ce(N__45906),
            .sr(N__45891));
    defparam comm_buf_2__i7_LC_17_13_1.C_ON=1'b0;
    defparam comm_buf_2__i7_LC_17_13_1.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i7_LC_17_13_1.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_2__i7_LC_17_13_1 (
            .in0(N__54547),
            .in1(N__48595),
            .in2(_gnd_net_),
            .in3(N__45519),
            .lcout(comm_buf_2_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56040),
            .ce(N__45906),
            .sr(N__45891));
    defparam comm_buf_2__i6_LC_17_13_2.C_ON=1'b0;
    defparam comm_buf_2__i6_LC_17_13_2.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i6_LC_17_13_2.LUT_INIT=16'b1110111000100010;
    LogicCell40 comm_buf_2__i6_LC_17_13_2 (
            .in0(N__45501),
            .in1(N__54551),
            .in2(_gnd_net_),
            .in3(N__53218),
            .lcout(comm_buf_2_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56040),
            .ce(N__45906),
            .sr(N__45891));
    defparam comm_buf_2__i5_LC_17_13_3.C_ON=1'b0;
    defparam comm_buf_2__i5_LC_17_13_3.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i5_LC_17_13_3.LUT_INIT=16'b1111010110100000;
    LogicCell40 comm_buf_2__i5_LC_17_13_3 (
            .in0(N__54546),
            .in1(_gnd_net_),
            .in2(N__53345),
            .in3(N__46005),
            .lcout(comm_buf_2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56040),
            .ce(N__45906),
            .sr(N__45891));
    defparam comm_buf_2__i4_LC_17_13_4.C_ON=1'b0;
    defparam comm_buf_2__i4_LC_17_13_4.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i4_LC_17_13_4.LUT_INIT=16'b1100110010101010;
    LogicCell40 comm_buf_2__i4_LC_17_13_4 (
            .in0(N__45990),
            .in1(N__53649),
            .in2(_gnd_net_),
            .in3(N__54550),
            .lcout(comm_buf_2_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56040),
            .ce(N__45906),
            .sr(N__45891));
    defparam comm_buf_2__i3_LC_17_13_5.C_ON=1'b0;
    defparam comm_buf_2__i3_LC_17_13_5.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i3_LC_17_13_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_2__i3_LC_17_13_5 (
            .in0(N__54545),
            .in1(N__49868),
            .in2(_gnd_net_),
            .in3(N__45963),
            .lcout(comm_buf_2_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56040),
            .ce(N__45906),
            .sr(N__45891));
    defparam comm_buf_2__i2_LC_17_13_6.C_ON=1'b0;
    defparam comm_buf_2__i2_LC_17_13_6.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i2_LC_17_13_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_2__i2_LC_17_13_6 (
            .in0(N__50165),
            .in1(N__45939),
            .in2(_gnd_net_),
            .in3(N__54549),
            .lcout(comm_buf_2_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56040),
            .ce(N__45906),
            .sr(N__45891));
    defparam comm_buf_2__i1_LC_17_13_7.C_ON=1'b0;
    defparam comm_buf_2__i1_LC_17_13_7.SEQ_MODE=4'b1000;
    defparam comm_buf_2__i1_LC_17_13_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_2__i1_LC_17_13_7 (
            .in0(N__54544),
            .in1(N__49723),
            .in2(_gnd_net_),
            .in3(N__45918),
            .lcout(comm_buf_2_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56040),
            .ce(N__45906),
            .sr(N__45891));
    defparam i1_2_lut_3_lut_adj_57_LC_17_14_1.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_57_LC_17_14_1.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_57_LC_17_14_1.LUT_INIT=16'b1010101000100010;
    LogicCell40 i1_2_lut_3_lut_adj_57_LC_17_14_1 (
            .in0(N__52090),
            .in1(N__54847),
            .in2(_gnd_net_),
            .in3(N__55270),
            .lcout(n16824),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i10_LC_17_14_2.C_ON=1'b0;
    defparam acadc_skipCount_i10_LC_17_14_2.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i10_LC_17_14_2.LUT_INIT=16'b0111001101000000;
    LogicCell40 acadc_skipCount_i10_LC_17_14_2 (
            .in0(N__49310),
            .in1(N__47920),
            .in2(N__45864),
            .in3(N__50607),
            .lcout(acadc_skipCount_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56056),
            .ce(),
            .sr(_gnd_net_));
    defparam i19161_2_lut_LC_17_14_3.C_ON=1'b0;
    defparam i19161_2_lut_LC_17_14_3.SEQ_MODE=4'b0000;
    defparam i19161_2_lut_LC_17_14_3.LUT_INIT=16'b0000000011001100;
    LogicCell40 i19161_2_lut_LC_17_14_3 (
            .in0(_gnd_net_),
            .in1(N__45768),
            .in2(_gnd_net_),
            .in3(N__57210),
            .lcout(n21543),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_128_Mux_2_i23_3_lut_LC_17_14_4.C_ON=1'b0;
    defparam mux_128_Mux_2_i23_3_lut_LC_17_14_4.SEQ_MODE=4'b0000;
    defparam mux_128_Mux_2_i23_3_lut_LC_17_14_4.LUT_INIT=16'b1110111001000100;
    LogicCell40 mux_128_Mux_2_i23_3_lut_LC_17_14_4 (
            .in0(N__57211),
            .in1(N__45728),
            .in2(_gnd_net_),
            .in3(N__50606),
            .lcout(n23_adj_1685),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i0_LC_17_14_6.C_ON=1'b0;
    defparam comm_buf_6__i0_LC_17_14_6.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i0_LC_17_14_6.LUT_INIT=16'b0100010011110000;
    LogicCell40 comm_buf_6__i0_LC_17_14_6 (
            .in0(N__55271),
            .in1(N__48698),
            .in2(N__46640),
            .in3(N__53128),
            .lcout(comm_buf_6_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56056),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i3_LC_17_14_7.C_ON=1'b0;
    defparam comm_buf_6__i3_LC_17_14_7.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i3_LC_17_14_7.LUT_INIT=16'b0100111001000100;
    LogicCell40 comm_buf_6__i3_LC_17_14_7 (
            .in0(N__53129),
            .in1(N__46616),
            .in2(N__55388),
            .in3(N__49877),
            .lcout(comm_buf_6_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56056),
            .ce(),
            .sr(_gnd_net_));
    defparam i18641_3_lut_LC_17_15_1.C_ON=1'b0;
    defparam i18641_3_lut_LC_17_15_1.SEQ_MODE=4'b0000;
    defparam i18641_3_lut_LC_17_15_1.LUT_INIT=16'b1110111001000100;
    LogicCell40 i18641_3_lut_LC_17_15_1 (
            .in0(N__46372),
            .in1(N__46602),
            .in2(_gnd_net_),
            .in3(N__46578),
            .lcout(n21368),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_129_Mux_7_i26_3_lut_LC_17_15_2.C_ON=1'b0;
    defparam mux_129_Mux_7_i26_3_lut_LC_17_15_2.SEQ_MODE=4'b0000;
    defparam mux_129_Mux_7_i26_3_lut_LC_17_15_2.LUT_INIT=16'b1011101110001000;
    LogicCell40 mux_129_Mux_7_i26_3_lut_LC_17_15_2 (
            .in0(N__46551),
            .in1(N__57252),
            .in2(_gnd_net_),
            .in3(N__46526),
            .lcout(),
            .ltout(n26_adj_1622_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18642_4_lut_LC_17_15_3.C_ON=1'b0;
    defparam i18642_4_lut_LC_17_15_3.SEQ_MODE=4'b0000;
    defparam i18642_4_lut_LC_17_15_3.LUT_INIT=16'b0100010011110000;
    LogicCell40 i18642_4_lut_LC_17_15_3 (
            .in0(N__57253),
            .in1(N__46500),
            .in2(N__46488),
            .in3(N__46373),
            .lcout(n21369),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_length_i0_LC_17_15_4.C_ON=1'b0;
    defparam comm_length_i0_LC_17_15_4.SEQ_MODE=4'b1000;
    defparam comm_length_i0_LC_17_15_4.LUT_INIT=16'b0001101000110110;
    LogicCell40 comm_length_i0_LC_17_15_4 (
            .in0(N__46374),
            .in1(N__47195),
            .in2(N__47708),
            .in3(N__57257),
            .lcout(comm_length_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56068),
            .ce(N__52095),
            .sr(N__46059));
    defparam comm_length_i1_LC_17_15_5.C_ON=1'b0;
    defparam comm_length_i1_LC_17_15_5.SEQ_MODE=4'b1000;
    defparam comm_length_i1_LC_17_15_5.LUT_INIT=16'b1101101011111101;
    LogicCell40 comm_length_i1_LC_17_15_5 (
            .in0(N__47194),
            .in1(N__47638),
            .in2(N__57273),
            .in3(N__46375),
            .lcout(comm_length_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56068),
            .ce(N__52095),
            .sr(N__46059));
    defparam i2_3_lut_adj_298_LC_17_15_7.C_ON=1'b0;
    defparam i2_3_lut_adj_298_LC_17_15_7.SEQ_MODE=4'b0000;
    defparam i2_3_lut_adj_298_LC_17_15_7.LUT_INIT=16'b1111111101100110;
    LogicCell40 i2_3_lut_adj_298_LC_17_15_7 (
            .in0(N__46047),
            .in1(N__52449),
            .in2(_gnd_net_),
            .in3(N__48429),
            .lcout(n5_adj_1524),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam acadc_skipCount_i12_LC_17_16_0.C_ON=1'b0;
    defparam acadc_skipCount_i12_LC_17_16_0.SEQ_MODE=4'b1000;
    defparam acadc_skipCount_i12_LC_17_16_0.LUT_INIT=16'b0111001101000000;
    LogicCell40 acadc_skipCount_i12_LC_17_16_0 (
            .in0(N__49309),
            .in1(N__47925),
            .in2(N__47815),
            .in3(N__50648),
            .lcout(acadc_skipCount_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56081),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_cmd_2__bdd_4_lut_LC_17_16_2.C_ON=1'b0;
    defparam comm_cmd_2__bdd_4_lut_LC_17_16_2.SEQ_MODE=4'b0000;
    defparam comm_cmd_2__bdd_4_lut_LC_17_16_2.LUT_INIT=16'b1110110001100100;
    LogicCell40 comm_cmd_2__bdd_4_lut_LC_17_16_2 (
            .in0(N__47262),
            .in1(N__47637),
            .in2(N__47316),
            .in3(N__47307),
            .lcout(),
            .ltout(n22599_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22599_bdd_4_lut_LC_17_16_3.C_ON=1'b0;
    defparam n22599_bdd_4_lut_LC_17_16_3.SEQ_MODE=4'b0000;
    defparam n22599_bdd_4_lut_LC_17_16_3.LUT_INIT=16'b1111000011001010;
    LogicCell40 n22599_bdd_4_lut_LC_17_16_3 (
            .in0(N__47301),
            .in1(N__47292),
            .in2(N__47274),
            .in3(N__47263),
            .lcout(n22602),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam buf_dds1_i6_LC_17_16_4.C_ON=1'b0;
    defparam buf_dds1_i6_LC_17_16_4.SEQ_MODE=4'b1000;
    defparam buf_dds1_i6_LC_17_16_4.LUT_INIT=16'b1110001000000000;
    LogicCell40 buf_dds1_i6_LC_17_16_4 (
            .in0(N__46957),
            .in1(N__46810),
            .in2(N__49487),
            .in3(N__46696),
            .lcout(buf_dds1_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56081),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_245_LC_17_16_6.C_ON=1'b0;
    defparam i1_4_lut_adj_245_LC_17_16_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_245_LC_17_16_6.LUT_INIT=16'b1011101100001011;
    LogicCell40 i1_4_lut_adj_245_LC_17_16_6 (
            .in0(N__55268),
            .in1(N__53775),
            .in2(N__46934),
            .in3(N__55574),
            .lcout(n12048),
            .ltout(n12048_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_4_lut_LC_17_16_7.C_ON=1'b0;
    defparam i1_2_lut_3_lut_4_lut_LC_17_16_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_4_lut_LC_17_16_7.LUT_INIT=16'b0001111100001111;
    LogicCell40 i1_2_lut_3_lut_4_lut_LC_17_16_7 (
            .in0(N__54843),
            .in1(N__54534),
            .in2(N__46770),
            .in3(N__55269),
            .lcout(n16971),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_clear_301_LC_17_17_0.C_ON=1'b0;
    defparam comm_clear_301_LC_17_17_0.SEQ_MODE=4'b1000;
    defparam comm_clear_301_LC_17_17_0.LUT_INIT=16'b0111011101010101;
    LogicCell40 comm_clear_301_LC_17_17_0 (
            .in0(N__54566),
            .in1(N__55387),
            .in2(_gnd_net_),
            .in3(N__53947),
            .lcout(comm_clear),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56088),
            .ce(N__50580),
            .sr(_gnd_net_));
    defparam \comm_spi.iclk_40_12283_12284_reset_LC_18_4_6 .C_ON=1'b0;
    defparam \comm_spi.iclk_40_12283_12284_reset_LC_18_4_6 .SEQ_MODE=4'b1010;
    defparam \comm_spi.iclk_40_12283_12284_reset_LC_18_4_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \comm_spi.iclk_40_12283_12284_reset_LC_18_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48137),
            .lcout(\comm_spi.n14805 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55947),
            .ce(),
            .sr(N__48090));
    defparam \comm_spi.RESET_I_0_90_2_lut_LC_18_5_5 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_90_2_lut_LC_18_5_5 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_90_2_lut_LC_18_5_5 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \comm_spi.RESET_I_0_90_2_lut_LC_18_5_5  (
            .in0(N__58054),
            .in1(N__48138),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\comm_spi.iclk_N_802 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_91_2_lut_LC_18_5_6 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_91_2_lut_LC_18_5_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_91_2_lut_LC_18_5_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \comm_spi.RESET_I_0_91_2_lut_LC_18_5_6  (
            .in0(_gnd_net_),
            .in1(N__58053),
            .in2(_gnd_net_),
            .in3(N__48139),
            .lcout(\comm_spi.iclk_N_803 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_adj_213_LC_18_6_5.C_ON=1'b0;
    defparam i1_2_lut_adj_213_LC_18_6_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_adj_213_LC_18_6_5.LUT_INIT=16'b1111111100110011;
    LogicCell40 i1_2_lut_adj_213_LC_18_6_5 (
            .in0(_gnd_net_),
            .in1(N__54874),
            .in2(_gnd_net_),
            .in3(N__55104),
            .lcout(n21110),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_5__i0_LC_18_7_0.C_ON=1'b0;
    defparam comm_buf_5__i0_LC_18_7_0.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i0_LC_18_7_0.LUT_INIT=16'b1110111000100010;
    LogicCell40 comm_buf_5__i0_LC_18_7_0 (
            .in0(N__48078),
            .in1(N__54197),
            .in2(_gnd_net_),
            .in3(N__48708),
            .lcout(comm_buf_5_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55971),
            .ce(N__48297),
            .sr(N__48276));
    defparam comm_buf_5__i7_LC_18_7_1.C_ON=1'b0;
    defparam comm_buf_5__i7_LC_18_7_1.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i7_LC_18_7_1.LUT_INIT=16'b1111010110100000;
    LogicCell40 comm_buf_5__i7_LC_18_7_1 (
            .in0(N__54196),
            .in1(_gnd_net_),
            .in2(N__48597),
            .in3(N__48066),
            .lcout(comm_buf_5_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55971),
            .ce(N__48297),
            .sr(N__48276));
    defparam comm_buf_5__i6_LC_18_7_2.C_ON=1'b0;
    defparam comm_buf_5__i6_LC_18_7_2.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i6_LC_18_7_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_5__i6_LC_18_7_2 (
            .in0(N__53226),
            .in1(N__48036),
            .in2(_gnd_net_),
            .in3(N__54200),
            .lcout(comm_buf_5_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55971),
            .ce(N__48297),
            .sr(N__48276));
    defparam comm_buf_5__i5_LC_18_7_3.C_ON=1'b0;
    defparam comm_buf_5__i5_LC_18_7_3.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i5_LC_18_7_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_5__i5_LC_18_7_3 (
            .in0(N__54195),
            .in1(N__53332),
            .in2(_gnd_net_),
            .in3(N__48021),
            .lcout(comm_buf_5_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55971),
            .ce(N__48297),
            .sr(N__48276));
    defparam comm_buf_5__i4_LC_18_7_4.C_ON=1'b0;
    defparam comm_buf_5__i4_LC_18_7_4.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i4_LC_18_7_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_5__i4_LC_18_7_4 (
            .in0(N__53645),
            .in1(N__48003),
            .in2(_gnd_net_),
            .in3(N__54199),
            .lcout(comm_buf_5_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55971),
            .ce(N__48297),
            .sr(N__48276));
    defparam comm_buf_5__i3_LC_18_7_5.C_ON=1'b0;
    defparam comm_buf_5__i3_LC_18_7_5.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i3_LC_18_7_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_5__i3_LC_18_7_5 (
            .in0(N__54194),
            .in1(N__49876),
            .in2(_gnd_net_),
            .in3(N__47973),
            .lcout(comm_buf_5_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55971),
            .ce(N__48297),
            .sr(N__48276));
    defparam comm_buf_5__i2_LC_18_7_6.C_ON=1'b0;
    defparam comm_buf_5__i2_LC_18_7_6.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i2_LC_18_7_6.LUT_INIT=16'b1100110010101010;
    LogicCell40 comm_buf_5__i2_LC_18_7_6 (
            .in0(N__47949),
            .in1(N__50146),
            .in2(_gnd_net_),
            .in3(N__54198),
            .lcout(comm_buf_5_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55971),
            .ce(N__48297),
            .sr(N__48276));
    defparam comm_buf_5__i1_LC_18_7_7.C_ON=1'b0;
    defparam comm_buf_5__i1_LC_18_7_7.SEQ_MODE=4'b1000;
    defparam comm_buf_5__i1_LC_18_7_7.LUT_INIT=16'b1111101001010000;
    LogicCell40 comm_buf_5__i1_LC_18_7_7 (
            .in0(N__54193),
            .in1(_gnd_net_),
            .in2(N__48309),
            .in3(N__49721),
            .lcout(comm_buf_5_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55971),
            .ce(N__48297),
            .sr(N__48276));
    defparam comm_state_1__bdd_4_lut_LC_18_8_0.C_ON=1'b0;
    defparam comm_state_1__bdd_4_lut_LC_18_8_0.SEQ_MODE=4'b0000;
    defparam comm_state_1__bdd_4_lut_LC_18_8_0.LUT_INIT=16'b1110011011000100;
    LogicCell40 comm_state_1__bdd_4_lut_LC_18_8_0 (
            .in0(N__54891),
            .in1(N__54173),
            .in2(N__52152),
            .in3(N__48267),
            .lcout(n22611),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_342_Mux_1_i2_3_lut_4_lut_LC_18_8_1.C_ON=1'b0;
    defparam comm_state_3__I_0_342_Mux_1_i2_3_lut_4_lut_LC_18_8_1.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_342_Mux_1_i2_3_lut_4_lut_LC_18_8_1.LUT_INIT=16'b0101000011001100;
    LogicCell40 comm_state_3__I_0_342_Mux_1_i2_3_lut_4_lut_LC_18_8_1 (
            .in0(N__48162),
            .in1(N__52690),
            .in2(N__54339),
            .in3(N__53872),
            .lcout(),
            .ltout(n2_adj_1576_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22611_bdd_4_lut_LC_18_8_2.C_ON=1'b0;
    defparam n22611_bdd_4_lut_LC_18_8_2.SEQ_MODE=4'b0000;
    defparam n22611_bdd_4_lut_LC_18_8_2.LUT_INIT=16'b1111101001000100;
    LogicCell40 n22611_bdd_4_lut_LC_18_8_2 (
            .in0(N__54892),
            .in1(N__53946),
            .in2(N__48201),
            .in3(N__48198),
            .lcout(n22614),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i227_2_lut_LC_18_8_3.C_ON=1'b0;
    defparam i227_2_lut_LC_18_8_3.SEQ_MODE=4'b0000;
    defparam i227_2_lut_LC_18_8_3.LUT_INIT=16'b0000000011001100;
    LogicCell40 i227_2_lut_LC_18_8_3 (
            .in0(_gnd_net_),
            .in1(N__52691),
            .in2(_gnd_net_),
            .in3(N__52881),
            .lcout(n1348),
            .ltout(n1348_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_3__I_0_342_Mux_1_i8_3_lut_4_lut_LC_18_8_4.C_ON=1'b0;
    defparam comm_state_3__I_0_342_Mux_1_i8_3_lut_4_lut_LC_18_8_4.SEQ_MODE=4'b0000;
    defparam comm_state_3__I_0_342_Mux_1_i8_3_lut_4_lut_LC_18_8_4.LUT_INIT=16'b0001101100010001;
    LogicCell40 comm_state_3__I_0_342_Mux_1_i8_3_lut_4_lut_LC_18_8_4 (
            .in0(N__53873),
            .in1(N__48192),
            .in2(N__48168),
            .in3(N__54177),
            .lcout(n8_adj_1577),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_4_lut_LC_18_8_5.C_ON=1'b0;
    defparam i2_3_lut_4_lut_LC_18_8_5.SEQ_MODE=4'b0000;
    defparam i2_3_lut_4_lut_LC_18_8_5.LUT_INIT=16'b1111111111111101;
    LogicCell40 i2_3_lut_4_lut_LC_18_8_5 (
            .in0(N__54172),
            .in1(N__53870),
            .in2(N__48408),
            .in3(N__52044),
            .lcout(),
            .ltout(n21139_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_302_LC_18_8_6.C_ON=1'b0;
    defparam i1_4_lut_adj_302_LC_18_8_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_302_LC_18_8_6.LUT_INIT=16'b1111000011010000;
    LogicCell40 i1_4_lut_adj_302_LC_18_8_6 (
            .in0(N__53871),
            .in1(N__55564),
            .in2(N__48165),
            .in3(N__48161),
            .lcout(n4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_i1_LC_18_8_7.C_ON=1'b0;
    defparam comm_state_i1_LC_18_8_7.SEQ_MODE=4'b1000;
    defparam comm_state_i1_LC_18_8_7.LUT_INIT=16'b0101110100001000;
    LogicCell40 comm_state_i1_LC_18_8_7 (
            .in0(N__55120),
            .in1(N__48153),
            .in2(N__49375),
            .in3(N__48147),
            .lcout(comm_state_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__55983),
            .ce(N__52113),
            .sr(_gnd_net_));
    defparam i2_4_lut_adj_303_LC_18_9_0.C_ON=1'b0;
    defparam i2_4_lut_adj_303_LC_18_9_0.SEQ_MODE=4'b0000;
    defparam i2_4_lut_adj_303_LC_18_9_0.LUT_INIT=16'b1110111100000000;
    LogicCell40 i2_4_lut_adj_303_LC_18_9_0 (
            .in0(N__48417),
            .in1(N__48358),
            .in2(N__52796),
            .in3(N__48462),
            .lcout(n21013),
            .ltout(n21013_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_LC_18_9_1.C_ON=1'b0;
    defparam i1_4_lut_LC_18_9_1.SEQ_MODE=4'b0000;
    defparam i1_4_lut_LC_18_9_1.LUT_INIT=16'b1110000000000000;
    LogicCell40 i1_4_lut_LC_18_9_1 (
            .in0(N__48359),
            .in1(N__52038),
            .in2(N__48456),
            .in3(N__48315),
            .lcout(n21035),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_4_lut_adj_312_LC_18_9_2.C_ON=1'b0;
    defparam i1_4_lut_4_lut_adj_312_LC_18_9_2.SEQ_MODE=4'b0000;
    defparam i1_4_lut_4_lut_adj_312_LC_18_9_2.LUT_INIT=16'b0111001111111011;
    LogicCell40 i1_4_lut_4_lut_adj_312_LC_18_9_2 (
            .in0(N__52863),
            .in1(N__54179),
            .in2(N__52795),
            .in3(N__53923),
            .lcout(n4_adj_1589),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_297_LC_18_9_3.C_ON=1'b0;
    defparam i1_4_lut_adj_297_LC_18_9_3.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_297_LC_18_9_3.LUT_INIT=16'b0111110110111110;
    LogicCell40 i1_4_lut_adj_297_LC_18_9_3 (
            .in0(N__52513),
            .in1(N__52938),
            .in2(N__48444),
            .in3(N__52055),
            .lcout(n4_adj_1623),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15288_2_lut_LC_18_9_4.C_ON=1'b0;
    defparam i15288_2_lut_LC_18_9_4.SEQ_MODE=4'b0000;
    defparam i15288_2_lut_LC_18_9_4.LUT_INIT=16'b1100110011111111;
    LogicCell40 i15288_2_lut_LC_18_9_4 (
            .in0(_gnd_net_),
            .in1(N__54178),
            .in2(_gnd_net_),
            .in3(N__53922),
            .lcout(n3),
            .ltout(n3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_4_lut_adj_305_LC_18_9_5.C_ON=1'b0;
    defparam i2_3_lut_4_lut_adj_305_LC_18_9_5.SEQ_MODE=4'b0000;
    defparam i2_3_lut_4_lut_adj_305_LC_18_9_5.LUT_INIT=16'b1111111011111111;
    LogicCell40 i2_3_lut_4_lut_adj_305_LC_18_9_5 (
            .in0(N__52781),
            .in1(N__48407),
            .in2(N__48363),
            .in3(N__52862),
            .lcout(),
            .ltout(n20095_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_46_LC_18_9_6.C_ON=1'b0;
    defparam i1_4_lut_adj_46_LC_18_9_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_46_LC_18_9_6.LUT_INIT=16'b1110000000000000;
    LogicCell40 i1_4_lut_adj_46_LC_18_9_6 (
            .in0(N__48360),
            .in1(N__48330),
            .in2(N__48324),
            .in3(N__48321),
            .lcout(n21033),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_3_lut_adj_314_LC_18_9_7.C_ON=1'b0;
    defparam i2_3_lut_adj_314_LC_18_9_7.SEQ_MODE=4'b0000;
    defparam i2_3_lut_adj_314_LC_18_9_7.LUT_INIT=16'b1110111011111111;
    LogicCell40 i2_3_lut_adj_314_LC_18_9_7 (
            .in0(N__52150),
            .in1(N__48792),
            .in2(_gnd_net_),
            .in3(N__52861),
            .lcout(n11619),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_4_lut_LC_18_10_3.C_ON=1'b0;
    defparam i1_3_lut_4_lut_LC_18_10_3.SEQ_MODE=4'b0000;
    defparam i1_3_lut_4_lut_LC_18_10_3.LUT_INIT=16'b1100100011111010;
    LogicCell40 i1_3_lut_4_lut_LC_18_10_3 (
            .in0(N__55537),
            .in1(N__55028),
            .in2(N__53986),
            .in3(N__54840),
            .lcout(n11600),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_state_i3_LC_18_10_4.C_ON=1'b0;
    defparam comm_state_i3_LC_18_10_4.SEQ_MODE=4'b1000;
    defparam comm_state_i3_LC_18_10_4.LUT_INIT=16'b0000100001011101;
    LogicCell40 comm_state_i3_LC_18_10_4 (
            .in0(N__55029),
            .in1(N__49401),
            .in2(N__49386),
            .in3(N__48891),
            .lcout(comm_state_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56010),
            .ce(N__48879),
            .sr(_gnd_net_));
    defparam i18492_3_lut_LC_18_10_5.C_ON=1'b0;
    defparam i18492_3_lut_LC_18_10_5.SEQ_MODE=4'b0000;
    defparam i18492_3_lut_LC_18_10_5.LUT_INIT=16'b1111111111101110;
    LogicCell40 i18492_3_lut_LC_18_10_5 (
            .in0(N__48870),
            .in1(N__48858),
            .in2(_gnd_net_),
            .in3(N__48831),
            .lcout(),
            .ltout(n21219_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_308_LC_18_10_6.C_ON=1'b0;
    defparam i1_4_lut_adj_308_LC_18_10_6.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_308_LC_18_10_6.LUT_INIT=16'b1100111000000000;
    LogicCell40 i1_4_lut_adj_308_LC_18_10_6 (
            .in0(N__48807),
            .in1(N__48791),
            .in2(N__48768),
            .in3(N__48741),
            .lcout(n21089),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_49_LC_18_10_7.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_49_LC_18_10_7.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_49_LC_18_10_7.LUT_INIT=16'b1010101010001000;
    LogicCell40 i1_2_lut_3_lut_adj_49_LC_18_10_7 (
            .in0(N__55536),
            .in1(N__54839),
            .in2(_gnd_net_),
            .in3(N__55027),
            .lcout(n21043),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_3__i0_LC_18_11_0.C_ON=1'b0;
    defparam comm_buf_3__i0_LC_18_11_0.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i0_LC_18_11_0.LUT_INIT=16'b1110111000100010;
    LogicCell40 comm_buf_3__i0_LC_18_11_0 (
            .in0(N__48720),
            .in1(N__54433),
            .in2(_gnd_net_),
            .in3(N__48707),
            .lcout(comm_buf_3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56026),
            .ce(N__49428),
            .sr(N__49413));
    defparam comm_buf_3__i7_LC_18_11_1.C_ON=1'b0;
    defparam comm_buf_3__i7_LC_18_11_1.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i7_LC_18_11_1.LUT_INIT=16'b1110111001000100;
    LogicCell40 comm_buf_3__i7_LC_18_11_1 (
            .in0(N__54432),
            .in1(N__48615),
            .in2(_gnd_net_),
            .in3(N__48600),
            .lcout(comm_buf_3_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56026),
            .ce(N__49428),
            .sr(N__49413));
    defparam comm_buf_3__i6_LC_18_11_2.C_ON=1'b0;
    defparam comm_buf_3__i6_LC_18_11_2.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i6_LC_18_11_2.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_3__i6_LC_18_11_2 (
            .in0(N__53225),
            .in1(N__48492),
            .in2(_gnd_net_),
            .in3(N__54436),
            .lcout(comm_buf_3_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56026),
            .ce(N__49428),
            .sr(N__49413));
    defparam comm_buf_3__i5_LC_18_11_3.C_ON=1'b0;
    defparam comm_buf_3__i5_LC_18_11_3.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i5_LC_18_11_3.LUT_INIT=16'b1111010110100000;
    LogicCell40 comm_buf_3__i5_LC_18_11_3 (
            .in0(N__54431),
            .in1(_gnd_net_),
            .in2(N__53344),
            .in3(N__48477),
            .lcout(comm_buf_3_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56026),
            .ce(N__49428),
            .sr(N__49413));
    defparam comm_buf_3__i4_LC_18_11_4.C_ON=1'b0;
    defparam comm_buf_3__i4_LC_18_11_4.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i4_LC_18_11_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_3__i4_LC_18_11_4 (
            .in0(N__53636),
            .in1(N__49905),
            .in2(_gnd_net_),
            .in3(N__54435),
            .lcout(comm_buf_3_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56026),
            .ce(N__49428),
            .sr(N__49413));
    defparam comm_buf_3__i3_LC_18_11_5.C_ON=1'b0;
    defparam comm_buf_3__i3_LC_18_11_5.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i3_LC_18_11_5.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_3__i3_LC_18_11_5 (
            .in0(N__54430),
            .in1(N__49875),
            .in2(_gnd_net_),
            .in3(N__49788),
            .lcout(comm_buf_3_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56026),
            .ce(N__49428),
            .sr(N__49413));
    defparam comm_buf_3__i2_LC_18_11_6.C_ON=1'b0;
    defparam comm_buf_3__i2_LC_18_11_6.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i2_LC_18_11_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_buf_3__i2_LC_18_11_6 (
            .in0(N__50156),
            .in1(N__49767),
            .in2(_gnd_net_),
            .in3(N__54434),
            .lcout(comm_buf_3_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56026),
            .ce(N__49428),
            .sr(N__49413));
    defparam comm_buf_3__i1_LC_18_11_7.C_ON=1'b0;
    defparam comm_buf_3__i1_LC_18_11_7.SEQ_MODE=4'b1000;
    defparam comm_buf_3__i1_LC_18_11_7.LUT_INIT=16'b1101110110001000;
    LogicCell40 comm_buf_3__i1_LC_18_11_7 (
            .in0(N__54429),
            .in1(N__49704),
            .in2(_gnd_net_),
            .in3(N__49632),
            .lcout(comm_buf_3_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56026),
            .ce(N__49428),
            .sr(N__49413));
    defparam mux_137_Mux_6_i4_3_lut_LC_18_12_0.C_ON=1'b0;
    defparam mux_137_Mux_6_i4_3_lut_LC_18_12_0.SEQ_MODE=4'b0000;
    defparam mux_137_Mux_6_i4_3_lut_LC_18_12_0.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_137_Mux_6_i4_3_lut_LC_18_12_0 (
            .in0(N__53031),
            .in1(N__49623),
            .in2(_gnd_net_),
            .in3(N__49614),
            .lcout(n4_adj_1581),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_0__bdd_4_lut_19789_LC_18_12_1.C_ON=1'b0;
    defparam comm_index_0__bdd_4_lut_19789_LC_18_12_1.SEQ_MODE=4'b0000;
    defparam comm_index_0__bdd_4_lut_19789_LC_18_12_1.LUT_INIT=16'b1111001110001000;
    LogicCell40 comm_index_0__bdd_4_lut_19789_LC_18_12_1 (
            .in0(N__49602),
            .in1(N__52394),
            .in2(N__49596),
            .in3(N__53032),
            .lcout(),
            .ltout(n22545_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22545_bdd_4_lut_LC_18_12_2.C_ON=1'b0;
    defparam n22545_bdd_4_lut_LC_18_12_2.SEQ_MODE=4'b0000;
    defparam n22545_bdd_4_lut_LC_18_12_2.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22545_bdd_4_lut_LC_18_12_2 (
            .in0(N__52395),
            .in1(N__49557),
            .in2(N__49500),
            .in3(N__49486),
            .lcout(n22548),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12463_2_lut_LC_18_12_3.C_ON=1'b0;
    defparam i12463_2_lut_LC_18_12_3.SEQ_MODE=4'b0000;
    defparam i12463_2_lut_LC_18_12_3.LUT_INIT=16'b1100110000000000;
    LogicCell40 i12463_2_lut_LC_18_12_3 (
            .in0(_gnd_net_),
            .in1(N__55164),
            .in2(_gnd_net_),
            .in3(N__49424),
            .lcout(n14979),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i2_LC_18_12_4.C_ON=1'b0;
    defparam comm_buf_6__i2_LC_18_12_4.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i2_LC_18_12_4.LUT_INIT=16'b0101000011001100;
    LogicCell40 comm_buf_6__i2_LC_18_12_4 (
            .in0(N__55165),
            .in1(N__50073),
            .in2(N__50169),
            .in3(N__53126),
            .lcout(comm_buf_6_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56041),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_137_Mux_0_i4_3_lut_LC_18_12_5.C_ON=1'b0;
    defparam mux_137_Mux_0_i4_3_lut_LC_18_12_5.SEQ_MODE=4'b0000;
    defparam mux_137_Mux_0_i4_3_lut_LC_18_12_5.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_137_Mux_0_i4_3_lut_LC_18_12_5 (
            .in0(N__50061),
            .in1(N__50049),
            .in2(_gnd_net_),
            .in3(N__53030),
            .lcout(n4_adj_1457),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_137_Mux_1_i4_3_lut_LC_18_12_6.C_ON=1'b0;
    defparam mux_137_Mux_1_i4_3_lut_LC_18_12_6.SEQ_MODE=4'b0000;
    defparam mux_137_Mux_1_i4_3_lut_LC_18_12_6.LUT_INIT=16'b1101110110001000;
    LogicCell40 mux_137_Mux_1_i4_3_lut_LC_18_12_6 (
            .in0(N__53033),
            .in1(N__50031),
            .in2(_gnd_net_),
            .in3(N__50019),
            .lcout(n4_adj_1588),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i12491_3_lut_LC_18_12_7.C_ON=1'b0;
    defparam i12491_3_lut_LC_18_12_7.SEQ_MODE=4'b0000;
    defparam i12491_3_lut_LC_18_12_7.LUT_INIT=16'b1000100010101010;
    LogicCell40 i12491_3_lut_LC_18_12_7 (
            .in0(N__50321),
            .in1(N__55163),
            .in2(_gnd_net_),
            .in3(N__50007),
            .lcout(n15007),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19086_2_lut_LC_18_13_3.C_ON=1'b0;
    defparam i19086_2_lut_LC_18_13_3.SEQ_MODE=4'b0000;
    defparam i19086_2_lut_LC_18_13_3.LUT_INIT=16'b0000000011001100;
    LogicCell40 i19086_2_lut_LC_18_13_3 (
            .in0(_gnd_net_),
            .in1(N__49977),
            .in2(_gnd_net_),
            .in3(N__53067),
            .lcout(),
            .ltout(n21433_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_1__bdd_4_lut_19741_LC_18_13_4.C_ON=1'b0;
    defparam comm_index_1__bdd_4_lut_19741_LC_18_13_4.SEQ_MODE=4'b0000;
    defparam comm_index_1__bdd_4_lut_19741_LC_18_13_4.LUT_INIT=16'b1110010010101010;
    LogicCell40 comm_index_1__bdd_4_lut_19741_LC_18_13_4 (
            .in0(N__52436),
            .in1(N__49959),
            .in2(N__49953),
            .in3(N__52562),
            .lcout(),
            .ltout(n22419_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i1_LC_18_13_5.C_ON=1'b0;
    defparam comm_tx_buf_i1_LC_18_13_5.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i1_LC_18_13_5.LUT_INIT=16'b1111010010100100;
    LogicCell40 comm_tx_buf_i1_LC_18_13_5 (
            .in0(N__52563),
            .in1(N__53358),
            .in2(N__49950),
            .in3(N__53517),
            .lcout(comm_tx_buf_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56057),
            .ce(N__50354),
            .sr(N__50227));
    defparam i2_2_lut_3_lut_adj_284_LC_18_13_6.C_ON=1'b0;
    defparam i2_2_lut_3_lut_adj_284_LC_18_13_6.SEQ_MODE=4'b0000;
    defparam i2_2_lut_3_lut_adj_284_LC_18_13_6.LUT_INIT=16'b1000100000000000;
    LogicCell40 i2_2_lut_3_lut_adj_284_LC_18_13_6 (
            .in0(N__52435),
            .in1(N__52561),
            .in2(_gnd_net_),
            .in3(N__49947),
            .lcout(),
            .ltout(n7_adj_1458_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_4_lut_adj_232_LC_18_13_7.C_ON=1'b0;
    defparam i1_4_lut_adj_232_LC_18_13_7.SEQ_MODE=4'b0000;
    defparam i1_4_lut_adj_232_LC_18_13_7.LUT_INIT=16'b1100110010000000;
    LogicCell40 i1_4_lut_adj_232_LC_18_13_7 (
            .in0(N__52890),
            .in1(N__55573),
            .in2(N__49908),
            .in3(N__55108),
            .lcout(n12477),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18555_4_lut_LC_18_14_1.C_ON=1'b0;
    defparam i18555_4_lut_LC_18_14_1.SEQ_MODE=4'b0000;
    defparam i18555_4_lut_LC_18_14_1.LUT_INIT=16'b0100010011100100;
    LogicCell40 i18555_4_lut_LC_18_14_1 (
            .in0(N__52438),
            .in1(N__50487),
            .in2(N__53088),
            .in3(N__53068),
            .lcout(),
            .ltout(n21282_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i6_LC_18_14_2.C_ON=1'b0;
    defparam comm_tx_buf_i6_LC_18_14_2.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i6_LC_18_14_2.LUT_INIT=16'b1111001111000000;
    LogicCell40 comm_tx_buf_i6_LC_18_14_2 (
            .in0(_gnd_net_),
            .in1(N__52566),
            .in2(N__50478),
            .in3(N__50475),
            .lcout(comm_tx_buf_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56069),
            .ce(N__50342),
            .sr(N__50250));
    defparam i15197_3_lut_LC_18_14_3.C_ON=1'b0;
    defparam i15197_3_lut_LC_18_14_3.SEQ_MODE=4'b0000;
    defparam i15197_3_lut_LC_18_14_3.LUT_INIT=16'b1101110110001000;
    LogicCell40 i15197_3_lut_LC_18_14_3 (
            .in0(N__52564),
            .in1(N__50433),
            .in2(_gnd_net_),
            .in3(N__50423),
            .lcout(),
            .ltout(n17698_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i18543_4_lut_LC_18_14_4.C_ON=1'b0;
    defparam i18543_4_lut_LC_18_14_4.SEQ_MODE=4'b0000;
    defparam i18543_4_lut_LC_18_14_4.LUT_INIT=16'b0010001011110000;
    LogicCell40 i18543_4_lut_LC_18_14_4 (
            .in0(N__50370),
            .in1(N__52565),
            .in2(N__50361),
            .in3(N__52437),
            .lcout(),
            .ltout(n21270_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_tx_buf_i5_LC_18_14_5.C_ON=1'b0;
    defparam comm_tx_buf_i5_LC_18_14_5.SEQ_MODE=4'b1000;
    defparam comm_tx_buf_i5_LC_18_14_5.LUT_INIT=16'b1111000011001100;
    LogicCell40 comm_tx_buf_i5_LC_18_14_5 (
            .in0(_gnd_net_),
            .in1(N__52182),
            .in2(N__50358),
            .in3(N__53069),
            .lcout(comm_tx_buf_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56069),
            .ce(N__50342),
            .sr(N__50250));
    defparam i6_4_lut_adj_274_LC_18_15_0.C_ON=1'b0;
    defparam i6_4_lut_adj_274_LC_18_15_0.SEQ_MODE=4'b0000;
    defparam i6_4_lut_adj_274_LC_18_15_0.LUT_INIT=16'b1111111111111110;
    LogicCell40 i6_4_lut_adj_274_LC_18_15_0 (
            .in0(N__50567),
            .in1(N__51005),
            .in2(N__50535),
            .in3(N__50181),
            .lcout(n20996),
            .ltout(n20996_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i15361_2_lut_LC_18_15_1.C_ON=1'b0;
    defparam i15361_2_lut_LC_18_15_1.SEQ_MODE=4'b0000;
    defparam i15361_2_lut_LC_18_15_1.LUT_INIT=16'b1010000010100000;
    LogicCell40 i15361_2_lut_LC_18_15_1 (
            .in0(N__51020),
            .in1(_gnd_net_),
            .in2(N__50184),
            .in3(_gnd_net_),
            .lcout(n10_adj_1528),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i5_4_lut_adj_273_LC_18_15_2.C_ON=1'b0;
    defparam i5_4_lut_adj_273_LC_18_15_2.SEQ_MODE=4'b0000;
    defparam i5_4_lut_adj_273_LC_18_15_2.LUT_INIT=16'b1111111111111110;
    LogicCell40 i5_4_lut_adj_273_LC_18_15_2 (
            .in0(N__50501),
            .in1(N__50516),
            .in2(N__50553),
            .in3(N__51044),
            .lcout(n12_adj_1663),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclk_294_LC_18_15_3.C_ON=1'b0;
    defparam dds0_mclk_294_LC_18_15_3.SEQ_MODE=4'b1000;
    defparam dds0_mclk_294_LC_18_15_3.LUT_INIT=16'b1010101001011010;
    LogicCell40 dds0_mclk_294_LC_18_15_3 (
            .in0(N__50729),
            .in1(_gnd_net_),
            .in2(N__51024),
            .in3(N__50175),
            .lcout(dds0_mclk),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVdds0_mclk_294C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_16MHz_I_0_3_lut_LC_18_15_4.C_ON=1'b0;
    defparam clk_16MHz_I_0_3_lut_LC_18_15_4.SEQ_MODE=4'b0000;
    defparam clk_16MHz_I_0_3_lut_LC_18_15_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 clk_16MHz_I_0_3_lut_LC_18_15_4 (
            .in0(N__50811),
            .in1(N__50730),
            .in2(_gnd_net_),
            .in3(N__50721),
            .lcout(DDS_MCLK),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i5_4_lut_adj_65_LC_18_15_6.C_ON=1'b0;
    defparam i5_4_lut_adj_65_LC_18_15_6.SEQ_MODE=4'b0000;
    defparam i5_4_lut_adj_65_LC_18_15_6.LUT_INIT=16'b0111110110111110;
    LogicCell40 i5_4_lut_adj_65_LC_18_15_6 (
            .in0(N__50670),
            .in1(N__50644),
            .in2(N__50628),
            .in3(N__50605),
            .lcout(n21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_3_lut_adj_272_LC_18_15_7.C_ON=1'b0;
    defparam i2_2_lut_3_lut_adj_272_LC_18_15_7.SEQ_MODE=4'b0000;
    defparam i2_2_lut_3_lut_adj_272_LC_18_15_7.LUT_INIT=16'b1111111110111011;
    LogicCell40 i2_2_lut_3_lut_adj_272_LC_18_15_7 (
            .in0(N__54342),
            .in1(N__55272),
            .in2(_gnd_net_),
            .in3(N__53987),
            .lcout(n11590),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3772__i0_LC_18_16_0.C_ON=1'b1;
    defparam dds0_mclkcnt_i7_3772__i0_LC_18_16_0.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3772__i0_LC_18_16_0.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3772__i0_LC_18_16_0 (
            .in0(_gnd_net_),
            .in1(N__50568),
            .in2(_gnd_net_),
            .in3(N__50556),
            .lcout(dds0_mclkcnt_0),
            .ltout(),
            .carryin(bfn_18_16_0_),
            .carryout(n19925),
            .clk(INVdds0_mclkcnt_i7_3772__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3772__i1_LC_18_16_1.C_ON=1'b1;
    defparam dds0_mclkcnt_i7_3772__i1_LC_18_16_1.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3772__i1_LC_18_16_1.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3772__i1_LC_18_16_1 (
            .in0(_gnd_net_),
            .in1(N__50552),
            .in2(_gnd_net_),
            .in3(N__50538),
            .lcout(dds0_mclkcnt_1),
            .ltout(),
            .carryin(n19925),
            .carryout(n19926),
            .clk(INVdds0_mclkcnt_i7_3772__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3772__i2_LC_18_16_2.C_ON=1'b1;
    defparam dds0_mclkcnt_i7_3772__i2_LC_18_16_2.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3772__i2_LC_18_16_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3772__i2_LC_18_16_2 (
            .in0(_gnd_net_),
            .in1(N__50534),
            .in2(_gnd_net_),
            .in3(N__50520),
            .lcout(dds0_mclkcnt_2),
            .ltout(),
            .carryin(n19926),
            .carryout(n19927),
            .clk(INVdds0_mclkcnt_i7_3772__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3772__i3_LC_18_16_3.C_ON=1'b1;
    defparam dds0_mclkcnt_i7_3772__i3_LC_18_16_3.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3772__i3_LC_18_16_3.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3772__i3_LC_18_16_3 (
            .in0(_gnd_net_),
            .in1(N__50517),
            .in2(_gnd_net_),
            .in3(N__50505),
            .lcout(dds0_mclkcnt_3),
            .ltout(),
            .carryin(n19927),
            .carryout(n19928),
            .clk(INVdds0_mclkcnt_i7_3772__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3772__i4_LC_18_16_4.C_ON=1'b1;
    defparam dds0_mclkcnt_i7_3772__i4_LC_18_16_4.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3772__i4_LC_18_16_4.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3772__i4_LC_18_16_4 (
            .in0(_gnd_net_),
            .in1(N__50502),
            .in2(_gnd_net_),
            .in3(N__50490),
            .lcout(dds0_mclkcnt_4),
            .ltout(),
            .carryin(n19928),
            .carryout(n19929),
            .clk(INVdds0_mclkcnt_i7_3772__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3772__i5_LC_18_16_5.C_ON=1'b1;
    defparam dds0_mclkcnt_i7_3772__i5_LC_18_16_5.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3772__i5_LC_18_16_5.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3772__i5_LC_18_16_5 (
            .in0(_gnd_net_),
            .in1(N__51045),
            .in2(_gnd_net_),
            .in3(N__51033),
            .lcout(dds0_mclkcnt_5),
            .ltout(),
            .carryin(n19929),
            .carryout(n19930),
            .clk(INVdds0_mclkcnt_i7_3772__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3772__i6_LC_18_16_6.C_ON=1'b1;
    defparam dds0_mclkcnt_i7_3772__i6_LC_18_16_6.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3772__i6_LC_18_16_6.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3772__i6_LC_18_16_6 (
            .in0(_gnd_net_),
            .in1(N__51030),
            .in2(_gnd_net_),
            .in3(N__51012),
            .lcout(dds0_mclkcnt_6),
            .ltout(),
            .carryin(n19930),
            .carryout(n19931),
            .clk(INVdds0_mclkcnt_i7_3772__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam dds0_mclkcnt_i7_3772__i7_LC_18_16_7.C_ON=1'b0;
    defparam dds0_mclkcnt_i7_3772__i7_LC_18_16_7.SEQ_MODE=4'b1000;
    defparam dds0_mclkcnt_i7_3772__i7_LC_18_16_7.LUT_INIT=16'b1100001100111100;
    LogicCell40 dds0_mclkcnt_i7_3772__i7_LC_18_16_7 (
            .in0(_gnd_net_),
            .in1(N__51006),
            .in2(_gnd_net_),
            .in3(N__51009),
            .lcout(dds0_mclkcnt_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVdds0_mclkcnt_i7_3772__i0C_net),
            .ce(),
            .sr(_gnd_net_));
    defparam i12205_2_lut_LC_18_17_3.C_ON=1'b0;
    defparam i12205_2_lut_LC_18_17_3.SEQ_MODE=4'b0000;
    defparam i12205_2_lut_LC_18_17_3.LUT_INIT=16'b0000000011001100;
    LogicCell40 i12205_2_lut_LC_18_17_3 (
            .in0(_gnd_net_),
            .in1(N__54516),
            .in2(_gnd_net_),
            .in3(N__55233),
            .lcout(n14716),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i3_12313_12314_set_LC_19_5_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i3_12313_12314_set_LC_19_5_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i3_12313_12314_set_LC_19_5_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \comm_spi.data_tx_i3_12313_12314_set_LC_19_5_0  (
            .in0(N__57417),
            .in1(N__57441),
            .in2(_gnd_net_),
            .in3(N__57399),
            .lcout(\comm_spi.n14834 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__58328),
            .ce(),
            .sr(N__50820));
    defparam \comm_spi.RESET_I_0_89_2_lut_LC_19_5_1 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_89_2_lut_LC_19_5_1 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_89_2_lut_LC_19_5_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \comm_spi.RESET_I_0_89_2_lut_LC_19_5_1  (
            .in0(_gnd_net_),
            .in1(N__50875),
            .in2(_gnd_net_),
            .in3(N__58051),
            .lcout(\comm_spi.imosi_N_793 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_96_2_lut_LC_19_5_2 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_96_2_lut_LC_19_5_2 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_96_2_lut_LC_19_5_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \comm_spi.RESET_I_0_96_2_lut_LC_19_5_2  (
            .in0(N__58052),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56154),
            .lcout(\comm_spi.data_tx_7__N_810 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.div_state_i1_LC_19_6_1 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.div_state_i1_LC_19_6_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.div_state_i1_LC_19_6_1 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \ADC_VDC.genclk.div_state_i1_LC_19_6_1  (
            .in0(N__56230),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56574),
            .lcout(\ADC_VDC.genclk.div_state_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVADC_VDC.genclk.div_state_i1C_net ),
            .ce(N__53691),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i19403_2_lut_LC_19_6_3 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i19403_2_lut_LC_19_6_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i19403_2_lut_LC_19_6_3 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \ADC_VDC.genclk.i19403_2_lut_LC_19_6_3  (
            .in0(N__56229),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56573),
            .lcout(\ADC_VDC.genclk.n11900 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i1_2_lut_adj_26_LC_19_6_4 .C_ON=1'b0;
    defparam \ADC_VDC.i1_2_lut_adj_26_LC_19_6_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i1_2_lut_adj_26_LC_19_6_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \ADC_VDC.i1_2_lut_adj_26_LC_19_6_4  (
            .in0(N__52005),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51903),
            .lcout(),
            .ltout(\ADC_VDC.n52_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.i16282_4_lut_LC_19_6_5 .C_ON=1'b0;
    defparam \ADC_VDC.i16282_4_lut_LC_19_6_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.i16282_4_lut_LC_19_6_5 .LUT_INIT=16'b1001100011011100;
    LogicCell40 \ADC_VDC.i16282_4_lut_LC_19_6_5  (
            .in0(N__51760),
            .in1(N__51479),
            .in2(N__51216),
            .in3(N__51204),
            .lcout(\ADC_VDC.n11905 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.t0off_i0_LC_19_7_0 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i0_LC_19_7_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i0_LC_19_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i0_LC_19_7_0  (
            .in0(_gnd_net_),
            .in1(N__56340),
            .in2(_gnd_net_),
            .in3(N__51063),
            .lcout(\ADC_VDC.genclk.t0off_0 ),
            .ltout(),
            .carryin(bfn_19_7_0_),
            .carryout(\ADC_VDC.genclk.n19888 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__52169),
            .sr(N__58977));
    defparam \ADC_VDC.genclk.t0off_i1_LC_19_7_1 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i1_LC_19_7_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i1_LC_19_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i1_LC_19_7_1  (
            .in0(_gnd_net_),
            .in1(N__56370),
            .in2(N__58743),
            .in3(N__51060),
            .lcout(\ADC_VDC.genclk.t0off_1 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19888 ),
            .carryout(\ADC_VDC.genclk.n19889 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__52169),
            .sr(N__58977));
    defparam \ADC_VDC.genclk.t0off_i2_LC_19_7_2 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i2_LC_19_7_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i2_LC_19_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i2_LC_19_7_2  (
            .in0(_gnd_net_),
            .in1(N__58656),
            .in2(N__53742),
            .in3(N__51057),
            .lcout(\ADC_VDC.genclk.t0off_2 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19889 ),
            .carryout(\ADC_VDC.genclk.n19890 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__52169),
            .sr(N__58977));
    defparam \ADC_VDC.genclk.t0off_i3_LC_19_7_3 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i3_LC_19_7_3 .SEQ_MODE=4'b1001;
    defparam \ADC_VDC.genclk.t0off_i3_LC_19_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i3_LC_19_7_3  (
            .in0(_gnd_net_),
            .in1(N__56279),
            .in2(N__58744),
            .in3(N__51054),
            .lcout(\ADC_VDC.genclk.t0off_3 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19890 ),
            .carryout(\ADC_VDC.genclk.n19891 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__52169),
            .sr(N__58977));
    defparam \ADC_VDC.genclk.t0off_i4_LC_19_7_4 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i4_LC_19_7_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i4_LC_19_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i4_LC_19_7_4  (
            .in0(_gnd_net_),
            .in1(N__58660),
            .in2(N__56358),
            .in3(N__51051),
            .lcout(\ADC_VDC.genclk.t0off_4 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19891 ),
            .carryout(\ADC_VDC.genclk.n19892 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__52169),
            .sr(N__58977));
    defparam \ADC_VDC.genclk.t0off_i5_LC_19_7_5 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i5_LC_19_7_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i5_LC_19_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i5_LC_19_7_5  (
            .in0(_gnd_net_),
            .in1(N__56264),
            .in2(N__58745),
            .in3(N__51048),
            .lcout(\ADC_VDC.genclk.t0off_5 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19892 ),
            .carryout(\ADC_VDC.genclk.n19893 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__52169),
            .sr(N__58977));
    defparam \ADC_VDC.genclk.t0off_i6_LC_19_7_6 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i6_LC_19_7_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i6_LC_19_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i6_LC_19_7_6  (
            .in0(_gnd_net_),
            .in1(N__58664),
            .in2(N__56385),
            .in3(N__52032),
            .lcout(\ADC_VDC.genclk.t0off_6 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19893 ),
            .carryout(\ADC_VDC.genclk.n19894 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__52169),
            .sr(N__58977));
    defparam \ADC_VDC.genclk.t0off_i7_LC_19_7_7 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i7_LC_19_7_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i7_LC_19_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i7_LC_19_7_7  (
            .in0(_gnd_net_),
            .in1(N__53726),
            .in2(N__58746),
            .in3(N__52029),
            .lcout(\ADC_VDC.genclk.t0off_7 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19894 ),
            .carryout(\ADC_VDC.genclk.n19895 ),
            .clk(\INVADC_VDC.genclk.t0off_i0C_net ),
            .ce(N__52169),
            .sr(N__58977));
    defparam \ADC_VDC.genclk.t0off_i8_LC_19_8_0 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i8_LC_19_8_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i8_LC_19_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i8_LC_19_8_0  (
            .in0(_gnd_net_),
            .in1(N__56250),
            .in2(N__58718),
            .in3(N__52026),
            .lcout(\ADC_VDC.genclk.t0off_8 ),
            .ltout(),
            .carryin(bfn_19_8_0_),
            .carryout(\ADC_VDC.genclk.n19896 ),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__52170),
            .sr(N__58972));
    defparam \ADC_VDC.genclk.t0off_i9_LC_19_8_1 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i9_LC_19_8_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i9_LC_19_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i9_LC_19_8_1  (
            .in0(_gnd_net_),
            .in1(N__58626),
            .in2(N__56184),
            .in3(N__52023),
            .lcout(\ADC_VDC.genclk.t0off_9 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19896 ),
            .carryout(\ADC_VDC.genclk.n19897 ),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__52170),
            .sr(N__58972));
    defparam \ADC_VDC.genclk.t0off_i10_LC_19_8_2 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i10_LC_19_8_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i10_LC_19_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i10_LC_19_8_2  (
            .in0(_gnd_net_),
            .in1(N__53711),
            .in2(N__58715),
            .in3(N__52020),
            .lcout(\ADC_VDC.genclk.t0off_10 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19897 ),
            .carryout(\ADC_VDC.genclk.n19898 ),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__52170),
            .sr(N__58972));
    defparam \ADC_VDC.genclk.t0off_i11_LC_19_8_3 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i11_LC_19_8_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i11_LC_19_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i11_LC_19_8_3  (
            .in0(_gnd_net_),
            .in1(N__58614),
            .in2(N__56541),
            .in3(N__52017),
            .lcout(\ADC_VDC.genclk.t0off_11 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19898 ),
            .carryout(\ADC_VDC.genclk.n19899 ),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__52170),
            .sr(N__58972));
    defparam \ADC_VDC.genclk.t0off_i12_LC_19_8_4 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i12_LC_19_8_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i12_LC_19_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i12_LC_19_8_4  (
            .in0(_gnd_net_),
            .in1(N__53756),
            .in2(N__58716),
            .in3(N__52014),
            .lcout(\ADC_VDC.genclk.t0off_12 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19899 ),
            .carryout(\ADC_VDC.genclk.n19900 ),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__52170),
            .sr(N__58972));
    defparam \ADC_VDC.genclk.t0off_i13_LC_19_8_5 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i13_LC_19_8_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i13_LC_19_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i13_LC_19_8_5  (
            .in0(_gnd_net_),
            .in1(N__58618),
            .in2(N__56298),
            .in3(N__52011),
            .lcout(\ADC_VDC.genclk.t0off_13 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19900 ),
            .carryout(\ADC_VDC.genclk.n19901 ),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__52170),
            .sr(N__58972));
    defparam \ADC_VDC.genclk.t0off_i14_LC_19_8_6 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0off_i14_LC_19_8_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i14_LC_19_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0off_i14_LC_19_8_6  (
            .in0(_gnd_net_),
            .in1(N__56199),
            .in2(N__58717),
            .in3(N__52008),
            .lcout(\ADC_VDC.genclk.t0off_14 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19901 ),
            .carryout(\ADC_VDC.genclk.n19902 ),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__52170),
            .sr(N__58972));
    defparam \ADC_VDC.genclk.t0off_i15_LC_19_8_7 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.t0off_i15_LC_19_8_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0off_i15_LC_19_8_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ADC_VDC.genclk.t0off_i15_LC_19_8_7  (
            .in0(N__56168),
            .in1(N__58622),
            .in2(_gnd_net_),
            .in3(N__52173),
            .lcout(\ADC_VDC.genclk.t0off_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVADC_VDC.genclk.t0off_i8C_net ),
            .ce(N__52170),
            .sr(N__58972));
    defparam i19104_2_lut_3_lut_LC_19_9_0.C_ON=1'b0;
    defparam i19104_2_lut_3_lut_LC_19_9_0.SEQ_MODE=4'b0000;
    defparam i19104_2_lut_3_lut_LC_19_9_0.LUT_INIT=16'b0000000001000100;
    LogicCell40 i19104_2_lut_3_lut_LC_19_9_0 (
            .in0(N__52763),
            .in1(N__54183),
            .in2(_gnd_net_),
            .in3(N__52857),
            .lcout(n21453),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_2_lut_adj_306_LC_19_9_1.C_ON=1'b0;
    defparam i2_2_lut_adj_306_LC_19_9_1.SEQ_MODE=4'b0000;
    defparam i2_2_lut_adj_306_LC_19_9_1.LUT_INIT=16'b1100110011111111;
    LogicCell40 i2_2_lut_adj_306_LC_19_9_1 (
            .in0(_gnd_net_),
            .in1(N__52767),
            .in2(_gnd_net_),
            .in3(N__53919),
            .lcout(n14350),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19264_4_lut_4_lut_LC_19_9_2.C_ON=1'b0;
    defparam i19264_4_lut_4_lut_LC_19_9_2.SEQ_MODE=4'b0000;
    defparam i19264_4_lut_4_lut_LC_19_9_2.LUT_INIT=16'b0001001000010000;
    LogicCell40 i19264_4_lut_4_lut_LC_19_9_2 (
            .in0(N__54875),
            .in1(N__54184),
            .in2(N__52793),
            .in3(N__52858),
            .lcout(),
            .ltout(n21454_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19433_4_lut_LC_19_9_3.C_ON=1'b0;
    defparam i19433_4_lut_LC_19_9_3.SEQ_MODE=4'b0000;
    defparam i19433_4_lut_LC_19_9_3.LUT_INIT=16'b1100111111011101;
    LogicCell40 i19433_4_lut_LC_19_9_3 (
            .in0(N__52122),
            .in1(N__55065),
            .in2(N__52116),
            .in3(N__53921),
            .lcout(n14_adj_1638),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_length_i2_LC_19_9_4.C_ON=1'b0;
    defparam comm_length_i2_LC_19_9_4.SEQ_MODE=4'b1000;
    defparam comm_length_i2_LC_19_9_4.LUT_INIT=16'b1010101011001100;
    LogicCell40 comm_length_i2_LC_19_9_4 (
            .in0(N__52107),
            .in1(N__52056),
            .in2(_gnd_net_),
            .in3(N__52094),
            .lcout(comm_length_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56011),
            .ce(),
            .sr(_gnd_net_));
    defparam i3881_2_lut_3_lut_LC_19_9_5.C_ON=1'b0;
    defparam i3881_2_lut_3_lut_LC_19_9_5.SEQ_MODE=4'b0000;
    defparam i3881_2_lut_3_lut_LC_19_9_5.LUT_INIT=16'b0010001000000000;
    LogicCell40 i3881_2_lut_3_lut_LC_19_9_5 (
            .in0(N__52860),
            .in1(N__52769),
            .in2(_gnd_net_),
            .in3(N__52986),
            .lcout(n6401),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i4211_2_lut_LC_19_9_6.C_ON=1'b0;
    defparam i4211_2_lut_LC_19_9_6.SEQ_MODE=4'b0000;
    defparam i4211_2_lut_LC_19_9_6.LUT_INIT=16'b1111111110101010;
    LogicCell40 i4211_2_lut_LC_19_9_6 (
            .in0(N__52770),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__52856),
            .lcout(n6541),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i2_4_lut_4_lut_LC_19_9_7.C_ON=1'b0;
    defparam i2_4_lut_4_lut_LC_19_9_7.SEQ_MODE=4'b0000;
    defparam i2_4_lut_4_lut_LC_19_9_7.LUT_INIT=16'b0100111111101111;
    LogicCell40 i2_4_lut_4_lut_LC_19_9_7 (
            .in0(N__52859),
            .in1(N__52768),
            .in2(N__54340),
            .in3(N__53920),
            .lcout(n21154),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_i1_LC_19_10_0.C_ON=1'b0;
    defparam comm_index_i1_LC_19_10_0.SEQ_MODE=4'b1000;
    defparam comm_index_i1_LC_19_10_0.LUT_INIT=16'b1100011011001100;
    LogicCell40 comm_index_i1_LC_19_10_0 (
            .in0(N__52987),
            .in1(N__52376),
            .in2(N__52794),
            .in3(N__52880),
            .lcout(comm_index_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56027),
            .ce(N__54903),
            .sr(N__52647));
    defparam comm_index_i0_LC_19_10_1.C_ON=1'b0;
    defparam comm_index_i0_LC_19_10_1.SEQ_MODE=4'b1000;
    defparam comm_index_i0_LC_19_10_1.LUT_INIT=16'b1101110100100010;
    LogicCell40 comm_index_i0_LC_19_10_1 (
            .in0(N__52879),
            .in1(N__52771),
            .in2(_gnd_net_),
            .in3(N__52988),
            .lcout(comm_index_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56027),
            .ce(N__54903),
            .sr(N__52647));
    defparam comm_index_i2_LC_19_10_2.C_ON=1'b0;
    defparam comm_index_i2_LC_19_10_2.SEQ_MODE=4'b1000;
    defparam comm_index_i2_LC_19_10_2.LUT_INIT=16'b0111011110001000;
    LogicCell40 comm_index_i2_LC_19_10_2 (
            .in0(N__52653),
            .in1(N__52377),
            .in2(_gnd_net_),
            .in3(N__52512),
            .lcout(comm_index_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56027),
            .ce(N__54903),
            .sr(N__52647));
    defparam \comm_spi.data_tx_i5_12321_12322_set_LC_19_11_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i5_12321_12322_set_LC_19_11_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i5_12321_12322_set_LC_19_11_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \comm_spi.data_tx_i5_12321_12322_set_LC_19_11_0  (
            .in0(N__57492),
            .in1(N__57537),
            .in2(_gnd_net_),
            .in3(N__57515),
            .lcout(\comm_spi.n14842 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__58392),
            .ce(),
            .sr(N__53655));
    defparam i19106_2_lut_LC_19_11_2.C_ON=1'b0;
    defparam i19106_2_lut_LC_19_11_2.SEQ_MODE=4'b0000;
    defparam i19106_2_lut_LC_19_11_2.LUT_INIT=16'b0000000011001100;
    LogicCell40 i19106_2_lut_LC_19_11_2 (
            .in0(_gnd_net_),
            .in1(N__52602),
            .in2(_gnd_net_),
            .in3(N__57267),
            .lcout(n21460),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_102_2_lut_LC_19_12_0 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_102_2_lut_LC_19_12_0 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_102_2_lut_LC_19_12_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \comm_spi.RESET_I_0_102_2_lut_LC_19_12_0  (
            .in0(N__53674),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58126),
            .lcout(\comm_spi.data_tx_7__N_820 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i19515_4_lut_3_lut_LC_19_12_1 .C_ON=1'b0;
    defparam \comm_spi.i19515_4_lut_3_lut_LC_19_12_1 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19515_4_lut_3_lut_LC_19_12_1 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \comm_spi.i19515_4_lut_3_lut_LC_19_12_1  (
            .in0(N__56448),
            .in1(_gnd_net_),
            .in2(N__58160),
            .in3(N__57535),
            .lcout(\comm_spi.n23098 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_index_2__bdd_4_lut_LC_19_12_2.C_ON=1'b0;
    defparam comm_index_2__bdd_4_lut_LC_19_12_2.SEQ_MODE=4'b0000;
    defparam comm_index_2__bdd_4_lut_LC_19_12_2.LUT_INIT=16'b1111100000111000;
    LogicCell40 comm_index_2__bdd_4_lut_LC_19_12_2 (
            .in0(N__52578),
            .in1(N__52392),
            .in2(N__52554),
            .in3(N__53267),
            .lcout(),
            .ltout(n22503_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam n22503_bdd_4_lut_LC_19_12_3.C_ON=1'b0;
    defparam n22503_bdd_4_lut_LC_19_12_3.SEQ_MODE=4'b0000;
    defparam n22503_bdd_4_lut_LC_19_12_3.LUT_INIT=16'b1111010010100100;
    LogicCell40 n22503_bdd_4_lut_LC_19_12_3 (
            .in0(N__52393),
            .in1(N__52278),
            .in2(N__52200),
            .in3(N__52197),
            .lcout(n22506),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_94_2_lut_LC_19_12_4 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_94_2_lut_LC_19_12_4 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_94_2_lut_LC_19_12_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \comm_spi.RESET_I_0_94_2_lut_LC_19_12_4  (
            .in0(N__53675),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58127),
            .lcout(\comm_spi.data_tx_7__N_808 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i4_LC_19_12_5.C_ON=1'b0;
    defparam comm_buf_6__i4_LC_19_12_5.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i4_LC_19_12_5.LUT_INIT=16'b0000110010101010;
    LogicCell40 comm_buf_6__i4_LC_19_12_5 (
            .in0(N__53552),
            .in1(N__53620),
            .in2(N__55285),
            .in3(N__53130),
            .lcout(comm_buf_6_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56058),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_137_Mux_1_i2_3_lut_LC_19_12_6.C_ON=1'b0;
    defparam mux_137_Mux_1_i2_3_lut_LC_19_12_6.SEQ_MODE=4'b0000;
    defparam mux_137_Mux_1_i2_3_lut_LC_19_12_6.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_137_Mux_1_i2_3_lut_LC_19_12_6 (
            .in0(N__53538),
            .in1(N__53529),
            .in2(_gnd_net_),
            .in3(N__53042),
            .lcout(n2_adj_1587),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam mux_137_Mux_1_i1_3_lut_LC_19_13_1.C_ON=1'b0;
    defparam mux_137_Mux_1_i1_3_lut_LC_19_13_1.SEQ_MODE=4'b0000;
    defparam mux_137_Mux_1_i1_3_lut_LC_19_13_1.LUT_INIT=16'b1010101011001100;
    LogicCell40 mux_137_Mux_1_i1_3_lut_LC_19_13_1 (
            .in0(N__53503),
            .in1(N__53424),
            .in2(_gnd_net_),
            .in3(N__53029),
            .lcout(n1_adj_1586),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i5_LC_19_13_5.C_ON=1'b0;
    defparam comm_buf_6__i5_LC_19_13_5.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i5_LC_19_13_5.LUT_INIT=16'b0011000010101010;
    LogicCell40 comm_buf_6__i5_LC_19_13_5 (
            .in0(N__53268),
            .in1(N__55180),
            .in2(N__53349),
            .in3(N__53127),
            .lcout(comm_buf_6_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56070),
            .ce(),
            .sr(_gnd_net_));
    defparam i19164_2_lut_LC_19_13_6.C_ON=1'b0;
    defparam i19164_2_lut_LC_19_13_6.SEQ_MODE=4'b0000;
    defparam i19164_2_lut_LC_19_13_6.LUT_INIT=16'b0000000011001100;
    LogicCell40 i19164_2_lut_LC_19_13_6 (
            .in0(_gnd_net_),
            .in1(N__53256),
            .in2(_gnd_net_),
            .in3(N__57266),
            .lcout(n21547),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_buf_6__i6_LC_19_14_0.C_ON=1'b0;
    defparam comm_buf_6__i6_LC_19_14_0.SEQ_MODE=4'b1000;
    defparam comm_buf_6__i6_LC_19_14_0.LUT_INIT=16'b0011000010101010;
    LogicCell40 comm_buf_6__i6_LC_19_14_0 (
            .in0(N__53087),
            .in1(N__55281),
            .in2(N__53234),
            .in3(N__53131),
            .lcout(comm_buf_6_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56082),
            .ce(),
            .sr(_gnd_net_));
    defparam i3_3_lut_LC_19_14_4.C_ON=1'b0;
    defparam i3_3_lut_LC_19_14_4.SEQ_MODE=4'b0000;
    defparam i3_3_lut_LC_19_14_4.LUT_INIT=16'b0011000000000000;
    LogicCell40 i3_3_lut_LC_19_14_4 (
            .in0(_gnd_net_),
            .in1(N__53028),
            .in2(N__54894),
            .in3(N__54417),
            .lcout(n8_adj_1456),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_104_2_lut_LC_19_14_6 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_104_2_lut_LC_19_14_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_104_2_lut_LC_19_14_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \comm_spi.RESET_I_0_104_2_lut_LC_19_14_6  (
            .in0(N__56147),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58113),
            .lcout(\comm_spi.data_tx_7__N_826 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam comm_response_302_LC_19_15_0.C_ON=1'b0;
    defparam comm_response_302_LC_19_15_0.SEQ_MODE=4'b1000;
    defparam comm_response_302_LC_19_15_0.LUT_INIT=16'b0000001101010000;
    LogicCell40 comm_response_302_LC_19_15_0 (
            .in0(N__54004),
            .in1(N__54887),
            .in2(N__54515),
            .in3(N__55280),
            .lcout(ICE_GPMI_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__56089),
            .ce(N__55599),
            .sr(_gnd_net_));
    defparam i17_3_lut_3_lut_LC_19_15_3.C_ON=1'b0;
    defparam i17_3_lut_3_lut_LC_19_15_3.SEQ_MODE=4'b0000;
    defparam i17_3_lut_3_lut_LC_19_15_3.LUT_INIT=16'b0001000110001000;
    LogicCell40 i17_3_lut_3_lut_LC_19_15_3 (
            .in0(N__54886),
            .in1(N__54410),
            .in2(_gnd_net_),
            .in3(N__54003),
            .lcout(),
            .ltout(n10_adj_1619_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_3_lut_adj_288_LC_19_15_4.C_ON=1'b0;
    defparam i1_3_lut_adj_288_LC_19_15_4.SEQ_MODE=4'b0000;
    defparam i1_3_lut_adj_288_LC_19_15_4.LUT_INIT=16'b1100110011000000;
    LogicCell40 i1_3_lut_adj_288_LC_19_15_4 (
            .in0(_gnd_net_),
            .in1(N__55578),
            .in2(N__55482),
            .in3(N__55279),
            .lcout(n12079),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i1_2_lut_3_lut_adj_227_LC_19_15_5.C_ON=1'b0;
    defparam i1_2_lut_3_lut_adj_227_LC_19_15_5.SEQ_MODE=4'b0000;
    defparam i1_2_lut_3_lut_adj_227_LC_19_15_5.LUT_INIT=16'b1111111111101110;
    LogicCell40 i1_2_lut_3_lut_adj_227_LC_19_15_5 (
            .in0(N__54885),
            .in1(N__54409),
            .in2(_gnd_net_),
            .in3(N__54002),
            .lcout(n10804),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i11_4_lut_LC_20_6_0 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i11_4_lut_LC_20_6_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i11_4_lut_LC_20_6_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i11_4_lut_LC_20_6_0  (
            .in0(N__53760),
            .in1(N__53741),
            .in2(N__53727),
            .in3(N__53712),
            .lcout(),
            .ltout(\ADC_VDC.genclk.n27_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i19142_4_lut_LC_20_6_1 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i19142_4_lut_LC_20_6_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i19142_4_lut_LC_20_6_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i19142_4_lut_LC_20_6_1  (
            .in0(N__56526),
            .in1(N__56238),
            .in2(N__53697),
            .in3(N__56328),
            .lcout(\ADC_VDC.genclk.n21598 ),
            .ltout(\ADC_VDC.genclk.n21598_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i19468_2_lut_4_lut_LC_20_6_2 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i19468_2_lut_4_lut_LC_20_6_2 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i19468_2_lut_4_lut_LC_20_6_2 .LUT_INIT=16'b0001101111111111;
    LogicCell40 \ADC_VDC.genclk.i19468_2_lut_4_lut_LC_20_6_2  (
            .in0(N__56578),
            .in1(N__56319),
            .in2(N__53694),
            .in3(N__56231),
            .lcout(\ADC_VDC.genclk.n6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i19033_4_lut_LC_20_6_3 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i19033_4_lut_LC_20_6_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i19033_4_lut_LC_20_6_3 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \ADC_VDC.genclk.i19033_4_lut_LC_20_6_3  (
            .in0(N__56381),
            .in1(N__56369),
            .in2(N__56357),
            .in3(N__56339),
            .lcout(\ADC_VDC.genclk.n21600 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i11_4_lut_adj_25_LC_20_7_0 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i11_4_lut_adj_25_LC_20_7_0 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i11_4_lut_adj_25_LC_20_7_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i11_4_lut_adj_25_LC_20_7_0  (
            .in0(N__57677),
            .in1(N__57816),
            .in2(N__57567),
            .in3(N__57858),
            .lcout(),
            .ltout(\ADC_VDC.genclk.n27_adj_1449_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i19193_4_lut_LC_20_7_1 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i19193_4_lut_LC_20_7_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i19193_4_lut_LC_20_7_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i19193_4_lut_LC_20_7_1  (
            .in0(N__56205),
            .in1(N__56517),
            .in2(N__56322),
            .in3(N__56304),
            .lcout(\ADC_VDC.genclk.n21597 ),
            .ltout(\ADC_VDC.genclk.n21597_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.div_state_i0_LC_20_7_2 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.div_state_i0_LC_20_7_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.div_state_i0_LC_20_7_2 .LUT_INIT=16'b1101100011111111;
    LogicCell40 \ADC_VDC.genclk.div_state_i0_LC_20_7_2  (
            .in0(N__56572),
            .in1(N__56313),
            .in2(N__56307),
            .in3(N__56232),
            .lcout(\ADC_VDC.genclk.div_state_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVADC_VDC.genclk.div_state_i0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i19022_4_lut_LC_20_7_3 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i19022_4_lut_LC_20_7_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i19022_4_lut_LC_20_7_3 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \ADC_VDC.genclk.i19022_4_lut_LC_20_7_3  (
            .in0(N__57587),
            .in1(N__57714),
            .in2(N__57636),
            .in3(N__57696),
            .lcout(\ADC_VDC.genclk.n21603 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i10_4_lut_LC_20_7_5 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i10_4_lut_LC_20_7_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i10_4_lut_LC_20_7_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i10_4_lut_LC_20_7_5  (
            .in0(N__56297),
            .in1(N__56280),
            .in2(N__56265),
            .in3(N__56249),
            .lcout(\ADC_VDC.genclk.n26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i19414_2_lut_LC_20_7_7 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i19414_2_lut_LC_20_7_7 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i19414_2_lut_LC_20_7_7 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \ADC_VDC.genclk.i19414_2_lut_LC_20_7_7  (
            .in0(_gnd_net_),
            .in1(N__56228),
            .in2(_gnd_net_),
            .in3(N__56571),
            .lcout(\ADC_VDC.genclk.n14894 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i12_4_lut_adj_23_LC_20_8_3 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i12_4_lut_adj_23_LC_20_8_3 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i12_4_lut_adj_23_LC_20_8_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i12_4_lut_adj_23_LC_20_8_3  (
            .in0(N__57774),
            .in1(N__57878),
            .in2(N__57753),
            .in3(N__57836),
            .lcout(\ADC_VDC.genclk.n28_adj_1447 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i12_4_lut_LC_20_8_4 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i12_4_lut_LC_20_8_4 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i12_4_lut_LC_20_8_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i12_4_lut_LC_20_8_4  (
            .in0(N__56198),
            .in1(N__56180),
            .in2(N__56169),
            .in3(N__56537),
            .lcout(\ADC_VDC.genclk.n28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.i10_4_lut_adj_24_LC_20_8_5 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.i10_4_lut_adj_24_LC_20_8_5 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.i10_4_lut_adj_24_LC_20_8_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \ADC_VDC.genclk.i10_4_lut_adj_24_LC_20_8_5  (
            .in0(N__57794),
            .in1(N__57897),
            .in2(N__57612),
            .in3(N__57657),
            .lcout(\ADC_VDC.genclk.n26_adj_1448 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i4_12317_12318_reset_LC_20_9_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i4_12317_12318_reset_LC_20_9_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i4_12317_12318_reset_LC_20_9_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i4_12317_12318_reset_LC_20_9_0  (
            .in0(N__56511),
            .in1(N__56486),
            .in2(_gnd_net_),
            .in3(N__57371),
            .lcout(\comm_spi.n14839 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__58384),
            .ce(),
            .sr(N__56466));
    defparam \comm_spi.data_tx_i2_12309_12310_set_LC_20_10_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i2_12309_12310_set_LC_20_10_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i2_12309_12310_set_LC_20_10_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i2_12309_12310_set_LC_20_10_0  (
            .in0(N__58800),
            .in1(N__58860),
            .in2(_gnd_net_),
            .in3(N__58910),
            .lcout(\comm_spi.n14830 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__58406),
            .ce(),
            .sr(N__56457));
    defparam \comm_spi.RESET_I_0_103_2_lut_LC_20_10_1 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_103_2_lut_LC_20_10_1 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_103_2_lut_LC_20_10_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \comm_spi.RESET_I_0_103_2_lut_LC_20_10_1  (
            .in0(_gnd_net_),
            .in1(N__56446),
            .in2(_gnd_net_),
            .in3(N__58131),
            .lcout(\comm_spi.data_tx_7__N_823 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_97_2_lut_LC_20_10_2 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_97_2_lut_LC_20_10_2 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_97_2_lut_LC_20_10_2 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \comm_spi.RESET_I_0_97_2_lut_LC_20_10_2  (
            .in0(N__56402),
            .in1(_gnd_net_),
            .in2(N__58162),
            .in3(_gnd_net_),
            .lcout(\comm_spi.data_tx_7__N_811 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_105_2_lut_LC_20_10_3 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_105_2_lut_LC_20_10_3 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_105_2_lut_LC_20_10_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \comm_spi.RESET_I_0_105_2_lut_LC_20_10_3  (
            .in0(_gnd_net_),
            .in1(N__56401),
            .in2(_gnd_net_),
            .in3(N__58132),
            .lcout(\comm_spi.data_tx_7__N_829 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_95_2_lut_LC_20_10_4 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_95_2_lut_LC_20_10_4 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_95_2_lut_LC_20_10_4 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \comm_spi.RESET_I_0_95_2_lut_LC_20_10_4  (
            .in0(N__56447),
            .in1(_gnd_net_),
            .in2(N__58161),
            .in3(_gnd_net_),
            .lcout(\comm_spi.data_tx_7__N_809 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i19505_4_lut_3_lut_LC_20_10_5 .C_ON=1'b0;
    defparam \comm_spi.i19505_4_lut_3_lut_LC_20_10_5 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19505_4_lut_3_lut_LC_20_10_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \comm_spi.i19505_4_lut_3_lut_LC_20_10_5  (
            .in0(N__57430),
            .in1(N__56403),
            .in2(_gnd_net_),
            .in3(N__58139),
            .lcout(\comm_spi.n23104 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i2_12309_12310_reset_LC_20_11_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i2_12309_12310_reset_LC_20_11_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i2_12309_12310_reset_LC_20_11_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i2_12309_12310_reset_LC_20_11_0  (
            .in0(N__58796),
            .in1(N__58856),
            .in2(_gnd_net_),
            .in3(N__58914),
            .lcout(\comm_spi.n14831 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__58367),
            .ce(),
            .sr(N__57546));
    defparam \comm_spi.data_tx_i5_12321_12322_reset_LC_20_12_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i5_12321_12322_reset_LC_20_12_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i5_12321_12322_reset_LC_20_12_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i5_12321_12322_reset_LC_20_12_0  (
            .in0(N__57536),
            .in1(N__57519),
            .in2(_gnd_net_),
            .in3(N__57491),
            .lcout(\comm_spi.n14843 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__58407),
            .ce(),
            .sr(N__57450));
    defparam \comm_spi.data_tx_i3_12313_12314_reset_LC_20_13_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i3_12313_12314_reset_LC_20_13_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i3_12313_12314_reset_LC_20_13_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i3_12313_12314_reset_LC_20_13_0  (
            .in0(N__57437),
            .in1(N__57413),
            .in2(_gnd_net_),
            .in3(N__57395),
            .lcout(\comm_spi.n14835 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__58412),
            .ce(),
            .sr(N__57354));
    defparam i19378_2_lut_LC_20_14_2.C_ON=1'b0;
    defparam i19378_2_lut_LC_20_14_2.SEQ_MODE=4'b0000;
    defparam i19378_2_lut_LC_20_14_2.LUT_INIT=16'b0000000011001100;
    LogicCell40 i19378_2_lut_LC_20_14_2 (
            .in0(_gnd_net_),
            .in1(N__57342),
            .in2(_gnd_net_),
            .in3(N__57127),
            .lcout(n21456),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19099_2_lut_LC_20_15_0.C_ON=1'b0;
    defparam i19099_2_lut_LC_20_15_0.SEQ_MODE=4'b0000;
    defparam i19099_2_lut_LC_20_15_0.LUT_INIT=16'b0000000011001100;
    LogicCell40 i19099_2_lut_LC_20_15_0 (
            .in0(_gnd_net_),
            .in1(N__57324),
            .in2(_gnd_net_),
            .in3(N__57264),
            .lcout(n21447),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19145_2_lut_LC_20_16_2.C_ON=1'b0;
    defparam i19145_2_lut_LC_20_16_2.SEQ_MODE=4'b0000;
    defparam i19145_2_lut_LC_20_16_2.LUT_INIT=16'b0000000010101010;
    LogicCell40 i19145_2_lut_LC_20_16_2 (
            .in0(N__57300),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57265),
            .lcout(n21512),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam i19302_2_lut_LC_20_17_4.C_ON=1'b0;
    defparam i19302_2_lut_LC_20_17_4.SEQ_MODE=4'b0000;
    defparam i19302_2_lut_LC_20_17_4.LUT_INIT=16'b0000000011001100;
    LogicCell40 i19302_2_lut_LC_20_17_4 (
            .in0(_gnd_net_),
            .in1(N__57279),
            .in2(_gnd_net_),
            .in3(N__57263),
            .lcout(n21434),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i0_12279_12280_reset_LC_22_5_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i0_12279_12280_reset_LC_22_5_0 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i0_12279_12280_reset_LC_22_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \comm_spi.data_tx_i0_12279_12280_reset_LC_22_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58721),
            .lcout(\comm_spi.n14801 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__58371),
            .ce(),
            .sr(N__58926));
    defparam \ADC_VDC.genclk.div_state_1__I_0_1_lut_LC_22_6_1 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.div_state_1__I_0_1_lut_LC_22_6_1 .SEQ_MODE=4'b0000;
    defparam \ADC_VDC.genclk.div_state_1__I_0_1_lut_LC_22_6_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \ADC_VDC.genclk.div_state_1__I_0_1_lut_LC_22_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56582),
            .lcout(\ADC_VDC.genclk.div_state_1__N_1432 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ADC_VDC.genclk.t0on_i0_LC_22_7_0 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i0_LC_22_7_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i0_LC_22_7_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i0_LC_22_7_0  (
            .in0(_gnd_net_),
            .in1(N__57713),
            .in2(_gnd_net_),
            .in3(N__57699),
            .lcout(\ADC_VDC.genclk.t0on_0 ),
            .ltout(),
            .carryin(bfn_22_7_0_),
            .carryout(\ADC_VDC.genclk.n19903 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__57735),
            .sr(N__58973));
    defparam \ADC_VDC.genclk.t0on_i1_LC_22_7_1 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i1_LC_22_7_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i1_LC_22_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i1_LC_22_7_1  (
            .in0(_gnd_net_),
            .in1(N__57695),
            .in2(N__58751),
            .in3(N__57681),
            .lcout(\ADC_VDC.genclk.t0on_1 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19903 ),
            .carryout(\ADC_VDC.genclk.n19904 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__57735),
            .sr(N__58973));
    defparam \ADC_VDC.genclk.t0on_i2_LC_22_7_2 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i2_LC_22_7_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i2_LC_22_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i2_LC_22_7_2  (
            .in0(_gnd_net_),
            .in1(N__58687),
            .in2(N__57678),
            .in3(N__57660),
            .lcout(\ADC_VDC.genclk.t0on_2 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19904 ),
            .carryout(\ADC_VDC.genclk.n19905 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__57735),
            .sr(N__58973));
    defparam \ADC_VDC.genclk.t0on_i3_LC_22_7_3 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i3_LC_22_7_3 .SEQ_MODE=4'b1001;
    defparam \ADC_VDC.genclk.t0on_i3_LC_22_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i3_LC_22_7_3  (
            .in0(_gnd_net_),
            .in1(N__57653),
            .in2(N__58752),
            .in3(N__57639),
            .lcout(\ADC_VDC.genclk.t0on_3 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19905 ),
            .carryout(\ADC_VDC.genclk.n19906 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__57735),
            .sr(N__58973));
    defparam \ADC_VDC.genclk.t0on_i4_LC_22_7_4 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i4_LC_22_7_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i4_LC_22_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i4_LC_22_7_4  (
            .in0(_gnd_net_),
            .in1(N__58691),
            .in2(N__57635),
            .in3(N__57615),
            .lcout(\ADC_VDC.genclk.t0on_4 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19906 ),
            .carryout(\ADC_VDC.genclk.n19907 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__57735),
            .sr(N__58973));
    defparam \ADC_VDC.genclk.t0on_i5_LC_22_7_5 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i5_LC_22_7_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i5_LC_22_7_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i5_LC_22_7_5  (
            .in0(_gnd_net_),
            .in1(N__57605),
            .in2(N__58753),
            .in3(N__57591),
            .lcout(\ADC_VDC.genclk.t0on_5 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19907 ),
            .carryout(\ADC_VDC.genclk.n19908 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__57735),
            .sr(N__58973));
    defparam \ADC_VDC.genclk.t0on_i6_LC_22_7_6 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i6_LC_22_7_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i6_LC_22_7_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i6_LC_22_7_6  (
            .in0(_gnd_net_),
            .in1(N__58695),
            .in2(N__57588),
            .in3(N__57570),
            .lcout(\ADC_VDC.genclk.t0on_6 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19908 ),
            .carryout(\ADC_VDC.genclk.n19909 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__57735),
            .sr(N__58973));
    defparam \ADC_VDC.genclk.t0on_i7_LC_22_7_7 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i7_LC_22_7_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i7_LC_22_7_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i7_LC_22_7_7  (
            .in0(_gnd_net_),
            .in1(N__57563),
            .in2(N__58754),
            .in3(N__57549),
            .lcout(\ADC_VDC.genclk.t0on_7 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19909 ),
            .carryout(\ADC_VDC.genclk.n19910 ),
            .clk(\INVADC_VDC.genclk.t0on_i0C_net ),
            .ce(N__57735),
            .sr(N__58973));
    defparam \ADC_VDC.genclk.t0on_i8_LC_22_8_0 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i8_LC_22_8_0 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i8_LC_22_8_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i8_LC_22_8_0  (
            .in0(_gnd_net_),
            .in1(N__57896),
            .in2(N__58750),
            .in3(N__57882),
            .lcout(\ADC_VDC.genclk.t0on_8 ),
            .ltout(),
            .carryin(bfn_22_8_0_),
            .carryout(\ADC_VDC.genclk.n19911 ),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__57734),
            .sr(N__58968));
    defparam \ADC_VDC.genclk.t0on_i9_LC_22_8_1 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i9_LC_22_8_1 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i9_LC_22_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i9_LC_22_8_1  (
            .in0(_gnd_net_),
            .in1(N__58683),
            .in2(N__57879),
            .in3(N__57861),
            .lcout(\ADC_VDC.genclk.t0on_9 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19911 ),
            .carryout(\ADC_VDC.genclk.n19912 ),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__57734),
            .sr(N__58968));
    defparam \ADC_VDC.genclk.t0on_i10_LC_22_8_2 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i10_LC_22_8_2 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i10_LC_22_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i10_LC_22_8_2  (
            .in0(_gnd_net_),
            .in1(N__57854),
            .in2(N__58747),
            .in3(N__57840),
            .lcout(\ADC_VDC.genclk.t0on_10 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19912 ),
            .carryout(\ADC_VDC.genclk.n19913 ),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__57734),
            .sr(N__58968));
    defparam \ADC_VDC.genclk.t0on_i11_LC_22_8_3 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i11_LC_22_8_3 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i11_LC_22_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i11_LC_22_8_3  (
            .in0(_gnd_net_),
            .in1(N__58671),
            .in2(N__57837),
            .in3(N__57819),
            .lcout(\ADC_VDC.genclk.t0on_11 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19913 ),
            .carryout(\ADC_VDC.genclk.n19914 ),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__57734),
            .sr(N__58968));
    defparam \ADC_VDC.genclk.t0on_i12_LC_22_8_4 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i12_LC_22_8_4 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i12_LC_22_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i12_LC_22_8_4  (
            .in0(_gnd_net_),
            .in1(N__57812),
            .in2(N__58748),
            .in3(N__57798),
            .lcout(\ADC_VDC.genclk.t0on_12 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19914 ),
            .carryout(\ADC_VDC.genclk.n19915 ),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__57734),
            .sr(N__58968));
    defparam \ADC_VDC.genclk.t0on_i13_LC_22_8_5 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i13_LC_22_8_5 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i13_LC_22_8_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i13_LC_22_8_5  (
            .in0(_gnd_net_),
            .in1(N__58675),
            .in2(N__57795),
            .in3(N__57777),
            .lcout(\ADC_VDC.genclk.t0on_13 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19915 ),
            .carryout(\ADC_VDC.genclk.n19916 ),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__57734),
            .sr(N__58968));
    defparam \ADC_VDC.genclk.t0on_i14_LC_22_8_6 .C_ON=1'b1;
    defparam \ADC_VDC.genclk.t0on_i14_LC_22_8_6 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i14_LC_22_8_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ADC_VDC.genclk.t0on_i14_LC_22_8_6  (
            .in0(_gnd_net_),
            .in1(N__57773),
            .in2(N__58749),
            .in3(N__57759),
            .lcout(\ADC_VDC.genclk.t0on_14 ),
            .ltout(),
            .carryin(\ADC_VDC.genclk.n19916 ),
            .carryout(\ADC_VDC.genclk.n19917 ),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__57734),
            .sr(N__58968));
    defparam \ADC_VDC.genclk.t0on_i15_LC_22_8_7 .C_ON=1'b0;
    defparam \ADC_VDC.genclk.t0on_i15_LC_22_8_7 .SEQ_MODE=4'b1000;
    defparam \ADC_VDC.genclk.t0on_i15_LC_22_8_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \ADC_VDC.genclk.t0on_i15_LC_22_8_7  (
            .in0(N__57749),
            .in1(N__58679),
            .in2(_gnd_net_),
            .in3(N__57756),
            .lcout(\ADC_VDC.genclk.t0on_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVADC_VDC.genclk.t0on_i8C_net ),
            .ce(N__57734),
            .sr(N__58968));
    defparam \comm_spi.RESET_I_0_2_lut_LC_22_9_1 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_2_lut_LC_22_9_1 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_2_lut_LC_22_9_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \comm_spi.RESET_I_0_2_lut_LC_22_9_1  (
            .in0(N__58163),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58193),
            .lcout(\comm_spi.data_tx_7__N_835 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i19530_4_lut_3_lut_LC_22_9_6 .C_ON=1'b0;
    defparam \comm_spi.i19530_4_lut_3_lut_LC_22_9_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19530_4_lut_3_lut_LC_22_9_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \comm_spi.i19530_4_lut_3_lut_LC_22_9_6  (
            .in0(N__58194),
            .in1(N__58891),
            .in2(_gnd_net_),
            .in3(N__58164),
            .lcout(\comm_spi.n23110 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i1_12305_12306_reset_LC_22_10_7 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i1_12305_12306_reset_LC_22_10_7 .SEQ_MODE=4'b1010;
    defparam \comm_spi.data_tx_i1_12305_12306_reset_LC_22_10_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i1_12305_12306_reset_LC_22_10_7  (
            .in0(N__58892),
            .in1(N__58431),
            .in2(_gnd_net_),
            .in3(N__58874),
            .lcout(\comm_spi.n14827 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__58408),
            .ce(),
            .sr(N__58830));
    defparam \comm_spi.data_tx_i1_12305_12306_set_LC_22_11_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i1_12305_12306_set_LC_22_11_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i1_12305_12306_set_LC_22_11_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \comm_spi.data_tx_i1_12305_12306_set_LC_22_11_0  (
            .in0(N__58896),
            .in1(N__58430),
            .in2(_gnd_net_),
            .in3(N__58875),
            .lcout(\comm_spi.n14826 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__58399),
            .ce(),
            .sr(N__58839));
    defparam \comm_spi.RESET_I_0_98_2_lut_LC_22_11_2 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_98_2_lut_LC_22_11_2 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_98_2_lut_LC_22_11_2 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \comm_spi.RESET_I_0_98_2_lut_LC_22_11_2  (
            .in0(N__58817),
            .in1(_gnd_net_),
            .in2(N__58166),
            .in3(_gnd_net_),
            .lcout(\comm_spi.data_tx_7__N_812 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.RESET_I_0_106_2_lut_LC_22_11_3 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_106_2_lut_LC_22_11_3 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_106_2_lut_LC_22_11_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \comm_spi.RESET_I_0_106_2_lut_LC_22_11_3  (
            .in0(_gnd_net_),
            .in1(N__58816),
            .in2(_gnd_net_),
            .in3(N__58149),
            .lcout(\comm_spi.data_tx_7__N_832 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.i19495_4_lut_3_lut_LC_22_11_6 .C_ON=1'b0;
    defparam \comm_spi.i19495_4_lut_3_lut_LC_22_11_6 .SEQ_MODE=4'b0000;
    defparam \comm_spi.i19495_4_lut_3_lut_LC_22_11_6 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \comm_spi.i19495_4_lut_3_lut_LC_22_11_6  (
            .in0(N__58818),
            .in1(_gnd_net_),
            .in2(N__58167),
            .in3(N__58789),
            .lcout(\comm_spi.n23107 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \comm_spi.data_tx_i0_12279_12280_set_LC_22_13_0 .C_ON=1'b0;
    defparam \comm_spi.data_tx_i0_12279_12280_set_LC_22_13_0 .SEQ_MODE=4'b1011;
    defparam \comm_spi.data_tx_i0_12279_12280_set_LC_22_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \comm_spi.data_tx_i0_12279_12280_set_LC_22_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58765),
            .lcout(\comm_spi.n14800 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__58413),
            .ce(),
            .sr(N__57903));
    defparam \comm_spi.RESET_I_0_99_2_lut_LC_22_14_5 .C_ON=1'b0;
    defparam \comm_spi.RESET_I_0_99_2_lut_LC_22_14_5 .SEQ_MODE=4'b0000;
    defparam \comm_spi.RESET_I_0_99_2_lut_LC_22_14_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \comm_spi.RESET_I_0_99_2_lut_LC_22_14_5  (
            .in0(N__58192),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58157),
            .lcout(\comm_spi.data_tx_7__N_813 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // zim
